magic
tech sky130
magscale 1 2
timestamp 1667449939
<< error_p >>
rect -1 2144 0 2158
rect -2 1984 -1 2000
rect -8 1942 0 1984
rect -2 1932 -1 1942
rect -2 1926 0 1932
rect -1 1918 0 1926
rect -1 1874 0 1888
rect -2 1714 -1 1730
rect -8 1672 0 1714
rect -2 1662 -1 1672
rect -2 1656 0 1662
rect -1 1648 0 1656
rect -1 1604 0 1618
rect -2 1444 -1 1460
rect -8 1402 0 1444
rect -2 1392 -1 1402
rect -2 1386 0 1392
rect -1 1378 0 1386
rect -1 1334 0 1348
rect -2 -1256 -1 -1250
rect -8 -1298 0 -1256
rect -2 -1308 -1 -1298
rect -2 -1314 0 -1308
rect -1 -1322 0 -1314
rect -1 -1366 0 -1352
rect -2 -1526 -1 -1510
rect -8 -1568 0 -1526
rect -2 -1578 -1 -1568
rect -2 -1584 0 -1578
rect -1 -1592 0 -1584
rect -1 -1636 0 -1622
rect -2 -1796 -1 -1780
rect -8 -1838 0 -1796
rect -2 -1848 -1 -1838
rect -2 -1854 0 -1848
rect -1 -1862 0 -1854
rect -1 -1906 0 -1892
rect -2 -2066 -1 -2050
rect -8 -2108 0 -2066
rect -2 -2118 -1 -2108
rect -2 -2124 0 -2118
rect -1 -2132 0 -2124
<< error_s >>
rect 14 2158 27 2174
rect 116 2172 129 2174
rect 82 2158 97 2172
rect 106 2158 136 2172
rect 197 2170 350 2216
rect 179 2158 371 2170
rect 414 2158 444 2172
rect 450 2158 463 2174
rect 551 2158 564 2174
rect 594 2158 607 2174
rect 696 2172 709 2174
rect 662 2158 677 2172
rect 686 2158 716 2172
rect 777 2170 930 2216
rect 759 2158 951 2170
rect 994 2158 1024 2172
rect 1030 2158 1043 2174
rect 1131 2158 1144 2174
rect 1174 2158 1187 2174
rect 1276 2172 1289 2174
rect 1242 2158 1257 2172
rect 1266 2158 1296 2172
rect 1357 2170 1510 2216
rect 1339 2158 1531 2170
rect 1574 2158 1604 2172
rect 1610 2158 1623 2174
rect 1711 2158 1724 2174
rect 1754 2158 1767 2174
rect 1856 2172 1869 2174
rect 1822 2158 1837 2172
rect 1846 2158 1876 2172
rect 1937 2170 2090 2216
rect 1919 2158 2111 2170
rect 2154 2158 2184 2172
rect 2190 2158 2203 2174
rect 2291 2158 2304 2174
rect 2334 2158 2347 2174
rect 2436 2172 2449 2174
rect 2402 2158 2417 2172
rect 2426 2158 2456 2172
rect 2517 2170 2670 2216
rect 2499 2158 2691 2170
rect 2734 2158 2764 2172
rect 2770 2158 2783 2174
rect 2871 2158 2884 2174
rect 2914 2158 2927 2174
rect 3016 2172 3029 2174
rect 2982 2158 2997 2172
rect 3006 2158 3036 2172
rect 3097 2170 3250 2216
rect 3079 2158 3271 2170
rect 3314 2158 3344 2172
rect 3350 2158 3363 2174
rect 3451 2158 3464 2174
rect 3494 2158 3507 2174
rect 3596 2172 3609 2174
rect 3562 2158 3577 2172
rect 3586 2158 3616 2172
rect 3677 2170 3830 2216
rect 3659 2158 3851 2170
rect 3894 2158 3924 2172
rect 3930 2158 3943 2174
rect 4031 2158 4044 2174
rect 4074 2158 4087 2174
rect 4176 2172 4189 2174
rect 4142 2158 4157 2172
rect 4166 2158 4196 2172
rect 4257 2170 4410 2216
rect 4239 2158 4431 2170
rect 4474 2158 4504 2172
rect 4510 2158 4523 2174
rect 4611 2158 4624 2174
rect 4654 2158 4667 2174
rect 4756 2172 4769 2222
rect 4722 2158 4737 2172
rect 4746 2158 4776 2172
rect 4837 2170 4990 2216
rect 4819 2158 5011 2170
rect 5054 2158 5084 2172
rect 5090 2158 5103 2222
rect 5191 2158 5204 2174
rect 5234 2158 5247 2174
rect 5336 2172 5349 2222
rect 5302 2158 5317 2172
rect 5326 2158 5356 2172
rect 5417 2170 5570 2216
rect 5399 2158 5591 2170
rect 5634 2158 5664 2172
rect 5670 2158 5683 2222
rect 5771 2158 5784 2174
rect 5814 2158 5827 2174
rect 5916 2172 5929 2222
rect 5882 2158 5897 2172
rect 5906 2158 5936 2172
rect 5997 2170 6150 2216
rect 5979 2158 6171 2170
rect 6214 2158 6244 2172
rect 6250 2158 6263 2222
rect 6351 2158 6364 2174
rect 6394 2158 6407 2174
rect 6496 2172 6509 2222
rect 6462 2158 6477 2172
rect 6486 2158 6516 2172
rect 6577 2170 6730 2216
rect 6559 2158 6751 2170
rect 6794 2158 6824 2172
rect 6830 2158 6843 2222
rect 6931 2158 6944 2174
rect 0 2144 6944 2158
rect 14 2040 27 2144
rect 72 2122 73 2132
rect 88 2122 101 2132
rect 72 2118 101 2122
rect 106 2118 136 2144
rect 154 2130 170 2132
rect 242 2130 295 2144
rect 243 2128 307 2130
rect 350 2128 365 2144
rect 414 2141 444 2144
rect 414 2138 450 2141
rect 380 2130 396 2132
rect 154 2118 169 2122
rect 72 2116 169 2118
rect 197 2116 365 2128
rect 381 2118 396 2122
rect 414 2119 453 2138
rect 472 2132 479 2133
rect 478 2125 479 2132
rect 462 2122 463 2125
rect 478 2122 491 2125
rect 414 2118 444 2119
rect 453 2118 459 2119
rect 462 2118 491 2122
rect 381 2117 491 2118
rect 381 2116 497 2117
rect 56 2108 107 2116
rect 56 2096 81 2108
rect 88 2096 107 2108
rect 138 2108 188 2116
rect 138 2100 154 2108
rect 161 2106 188 2108
rect 197 2106 418 2116
rect 161 2096 418 2106
rect 447 2108 497 2116
rect 447 2099 463 2108
rect 56 2088 107 2096
rect 154 2088 418 2096
rect 444 2096 463 2099
rect 470 2096 497 2108
rect 444 2088 497 2096
rect 72 2080 73 2088
rect 88 2080 101 2088
rect 72 2072 88 2080
rect 69 2065 88 2068
rect 69 2056 91 2065
rect 42 2046 91 2056
rect 42 2040 72 2046
rect 91 2041 96 2046
rect 14 2024 88 2040
rect 106 2032 136 2088
rect 171 2078 379 2088
rect 414 2084 459 2088
rect 462 2087 463 2088
rect 478 2087 491 2088
rect 197 2048 386 2078
rect 212 2045 386 2048
rect 205 2042 386 2045
rect 14 2022 27 2024
rect 42 2022 76 2024
rect 14 2006 88 2022
rect 115 2018 128 2032
rect 143 2018 159 2034
rect 205 2029 216 2042
rect 14 1984 27 2006
rect 42 1984 72 2006
rect 115 2002 177 2018
rect 205 2011 216 2027
rect 221 2022 231 2042
rect 241 2022 255 2042
rect 258 2029 267 2042
rect 283 2029 292 2042
rect 221 2011 255 2022
rect 258 2011 267 2027
rect 283 2011 292 2027
rect 299 2022 309 2042
rect 319 2022 333 2042
rect 334 2029 345 2042
rect 299 2011 333 2022
rect 334 2011 345 2027
rect 391 2018 407 2034
rect 414 2032 444 2084
rect 478 2080 479 2087
rect 463 2072 479 2080
rect 450 2040 463 2059
rect 478 2040 508 2056
rect 450 2024 524 2040
rect 450 2022 463 2024
rect 478 2022 512 2024
rect 115 2000 128 2002
rect 143 2000 177 2002
rect 115 1984 177 2000
rect 221 1995 237 1998
rect 299 1995 329 2006
rect 377 2002 423 2018
rect 450 2006 524 2022
rect 377 2000 411 2002
rect 376 1984 423 2000
rect 450 1984 463 2006
rect 478 1984 508 2006
rect 535 1984 536 2000
rect 551 1984 564 2144
rect 594 2040 607 2144
rect 652 2122 653 2132
rect 668 2122 681 2132
rect 652 2118 681 2122
rect 686 2118 716 2144
rect 734 2130 750 2132
rect 822 2130 875 2144
rect 823 2128 887 2130
rect 930 2128 945 2144
rect 994 2141 1024 2144
rect 994 2138 1030 2141
rect 960 2130 976 2132
rect 734 2118 749 2122
rect 652 2116 749 2118
rect 777 2116 945 2128
rect 961 2118 976 2122
rect 994 2119 1033 2138
rect 1052 2132 1059 2133
rect 1058 2125 1059 2132
rect 1042 2122 1043 2125
rect 1058 2122 1071 2125
rect 994 2118 1024 2119
rect 1033 2118 1039 2119
rect 1042 2118 1071 2122
rect 961 2117 1071 2118
rect 961 2116 1077 2117
rect 636 2108 687 2116
rect 636 2096 661 2108
rect 668 2096 687 2108
rect 718 2108 768 2116
rect 718 2100 734 2108
rect 741 2106 768 2108
rect 777 2106 998 2116
rect 741 2096 998 2106
rect 1027 2108 1077 2116
rect 1027 2099 1043 2108
rect 636 2088 687 2096
rect 734 2088 998 2096
rect 1024 2096 1043 2099
rect 1050 2096 1077 2108
rect 1024 2088 1077 2096
rect 652 2080 653 2088
rect 668 2080 681 2088
rect 652 2072 668 2080
rect 649 2065 668 2068
rect 649 2056 671 2065
rect 622 2046 671 2056
rect 622 2040 652 2046
rect 671 2041 676 2046
rect 594 2024 668 2040
rect 686 2032 716 2088
rect 751 2078 959 2088
rect 994 2084 1039 2088
rect 1042 2087 1043 2088
rect 1058 2087 1071 2088
rect 777 2048 966 2078
rect 792 2045 966 2048
rect 785 2042 966 2045
rect 594 2022 607 2024
rect 622 2022 656 2024
rect 594 2006 668 2022
rect 695 2018 708 2032
rect 723 2018 739 2034
rect 785 2029 796 2042
rect 578 1984 579 2000
rect 594 1984 607 2006
rect 622 1984 652 2006
rect 695 2002 757 2018
rect 785 2011 796 2027
rect 801 2022 811 2042
rect 821 2022 835 2042
rect 838 2029 847 2042
rect 863 2029 872 2042
rect 801 2011 835 2022
rect 838 2011 847 2027
rect 863 2011 872 2027
rect 879 2022 889 2042
rect 899 2022 913 2042
rect 914 2029 925 2042
rect 879 2011 913 2022
rect 914 2011 925 2027
rect 971 2018 987 2034
rect 994 2032 1024 2084
rect 1058 2080 1059 2087
rect 1043 2072 1059 2080
rect 1030 2040 1043 2059
rect 1058 2040 1088 2056
rect 1030 2024 1104 2040
rect 1030 2022 1043 2024
rect 1058 2022 1092 2024
rect 695 2000 708 2002
rect 723 2000 757 2002
rect 695 1984 757 2000
rect 801 1995 817 1998
rect 879 1995 909 2006
rect 957 2002 1003 2018
rect 1030 2006 1104 2022
rect 957 2000 991 2002
rect 956 1984 1003 2000
rect 1030 1984 1043 2006
rect 1058 1984 1088 2006
rect 1115 1984 1116 2000
rect 1131 1984 1144 2144
rect 1174 2040 1187 2144
rect 1232 2122 1233 2132
rect 1248 2122 1261 2132
rect 1232 2118 1261 2122
rect 1266 2118 1296 2144
rect 1314 2130 1330 2132
rect 1402 2130 1455 2144
rect 1403 2128 1467 2130
rect 1510 2128 1525 2144
rect 1574 2141 1604 2144
rect 1574 2138 1610 2141
rect 1540 2130 1556 2132
rect 1314 2118 1329 2122
rect 1232 2116 1329 2118
rect 1357 2116 1525 2128
rect 1541 2118 1556 2122
rect 1574 2119 1613 2138
rect 1632 2132 1639 2133
rect 1638 2125 1639 2132
rect 1622 2122 1623 2125
rect 1638 2122 1651 2125
rect 1574 2118 1604 2119
rect 1613 2118 1619 2119
rect 1622 2118 1651 2122
rect 1541 2117 1651 2118
rect 1541 2116 1657 2117
rect 1216 2108 1267 2116
rect 1216 2096 1241 2108
rect 1248 2096 1267 2108
rect 1298 2108 1348 2116
rect 1298 2100 1314 2108
rect 1321 2106 1348 2108
rect 1357 2106 1578 2116
rect 1321 2096 1578 2106
rect 1607 2108 1657 2116
rect 1607 2099 1623 2108
rect 1216 2088 1267 2096
rect 1314 2088 1578 2096
rect 1604 2096 1623 2099
rect 1630 2096 1657 2108
rect 1604 2088 1657 2096
rect 1232 2080 1233 2088
rect 1248 2080 1261 2088
rect 1232 2072 1248 2080
rect 1229 2065 1248 2068
rect 1229 2056 1251 2065
rect 1202 2046 1251 2056
rect 1202 2040 1232 2046
rect 1251 2041 1256 2046
rect 1174 2024 1248 2040
rect 1266 2032 1296 2088
rect 1331 2078 1539 2088
rect 1574 2084 1619 2088
rect 1622 2087 1623 2088
rect 1638 2087 1651 2088
rect 1357 2048 1546 2078
rect 1372 2045 1546 2048
rect 1365 2042 1546 2045
rect 1174 2022 1187 2024
rect 1202 2022 1236 2024
rect 1174 2006 1248 2022
rect 1275 2018 1288 2032
rect 1303 2018 1319 2034
rect 1365 2029 1376 2042
rect 1158 1984 1159 2000
rect 1174 1984 1187 2006
rect 1202 1984 1232 2006
rect 1275 2002 1337 2018
rect 1365 2011 1376 2027
rect 1381 2022 1391 2042
rect 1401 2022 1415 2042
rect 1418 2029 1427 2042
rect 1443 2029 1452 2042
rect 1381 2011 1415 2022
rect 1418 2011 1427 2027
rect 1443 2011 1452 2027
rect 1459 2022 1469 2042
rect 1479 2022 1493 2042
rect 1494 2029 1505 2042
rect 1459 2011 1493 2022
rect 1494 2011 1505 2027
rect 1551 2018 1567 2034
rect 1574 2032 1604 2084
rect 1638 2080 1639 2087
rect 1623 2072 1639 2080
rect 1610 2040 1623 2059
rect 1638 2040 1668 2056
rect 1610 2024 1684 2040
rect 1610 2022 1623 2024
rect 1638 2022 1672 2024
rect 1275 2000 1288 2002
rect 1303 2000 1337 2002
rect 1275 1984 1337 2000
rect 1381 1995 1397 1998
rect 1459 1995 1489 2006
rect 1537 2002 1583 2018
rect 1610 2006 1684 2022
rect 1537 2000 1571 2002
rect 1536 1984 1583 2000
rect 1610 1984 1623 2006
rect 1638 1984 1668 2006
rect 1695 1984 1696 2000
rect 1711 1984 1724 2144
rect 1754 2040 1767 2144
rect 1812 2122 1813 2132
rect 1828 2122 1841 2132
rect 1812 2118 1841 2122
rect 1846 2118 1876 2144
rect 1894 2130 1910 2132
rect 1982 2130 2035 2144
rect 1983 2128 2047 2130
rect 2090 2128 2105 2144
rect 2154 2141 2184 2144
rect 2154 2138 2190 2141
rect 2120 2130 2136 2132
rect 1894 2118 1909 2122
rect 1812 2116 1909 2118
rect 1937 2116 2105 2128
rect 2121 2118 2136 2122
rect 2154 2119 2193 2138
rect 2212 2132 2219 2133
rect 2218 2125 2219 2132
rect 2202 2122 2203 2125
rect 2218 2122 2231 2125
rect 2154 2118 2184 2119
rect 2193 2118 2199 2119
rect 2202 2118 2231 2122
rect 2121 2117 2231 2118
rect 2121 2116 2237 2117
rect 1796 2108 1847 2116
rect 1796 2096 1821 2108
rect 1828 2096 1847 2108
rect 1878 2108 1928 2116
rect 1878 2100 1894 2108
rect 1901 2106 1928 2108
rect 1937 2106 2158 2116
rect 1901 2096 2158 2106
rect 2187 2108 2237 2116
rect 2187 2099 2203 2108
rect 1796 2088 1847 2096
rect 1894 2088 2158 2096
rect 2184 2096 2203 2099
rect 2210 2096 2237 2108
rect 2184 2088 2237 2096
rect 1812 2080 1813 2088
rect 1828 2080 1841 2088
rect 1812 2072 1828 2080
rect 1809 2065 1828 2068
rect 1809 2056 1831 2065
rect 1782 2046 1831 2056
rect 1782 2040 1812 2046
rect 1831 2041 1836 2046
rect 1754 2024 1828 2040
rect 1846 2032 1876 2088
rect 1911 2078 2119 2088
rect 2154 2084 2199 2088
rect 2202 2087 2203 2088
rect 2218 2087 2231 2088
rect 1937 2048 2126 2078
rect 1952 2045 2126 2048
rect 1945 2043 2126 2045
rect 1945 2042 2116 2043
rect 1754 2022 1767 2024
rect 1782 2022 1816 2024
rect 1754 2006 1828 2022
rect 1855 2018 1868 2032
rect 1883 2018 1899 2034
rect 1945 2029 1956 2042
rect 1738 1984 1739 2000
rect 1754 1984 1767 2006
rect 1782 1984 1812 2006
rect 1855 2002 1917 2018
rect 1945 2011 1956 2027
rect 1961 2022 1971 2042
rect 1981 2022 1995 2042
rect 1998 2029 2007 2042
rect 2023 2029 2032 2042
rect 1961 2011 1995 2022
rect 1998 2011 2007 2027
rect 2023 2011 2032 2027
rect 2039 2022 2049 2042
rect 2059 2022 2073 2042
rect 2074 2029 2085 2042
rect 2039 2011 2073 2022
rect 2074 2011 2085 2027
rect 2131 2018 2147 2034
rect 2154 2032 2184 2084
rect 2218 2080 2219 2087
rect 2203 2072 2219 2080
rect 2190 2040 2203 2059
rect 2218 2040 2248 2056
rect 2190 2024 2264 2040
rect 2190 2022 2203 2024
rect 2218 2022 2252 2024
rect 1855 2000 1868 2002
rect 1883 2000 1917 2002
rect 1855 1984 1917 2000
rect 1961 1995 1977 1998
rect 2039 1995 2069 2006
rect 2117 2002 2163 2018
rect 2190 2006 2264 2022
rect 2117 2000 2151 2002
rect 2116 1984 2163 2000
rect 2190 1984 2203 2006
rect 2218 1984 2248 2006
rect 2275 1984 2276 2000
rect 2291 1984 2304 2144
rect 2334 2040 2347 2144
rect 2392 2122 2393 2132
rect 2408 2122 2421 2132
rect 2392 2118 2421 2122
rect 2426 2118 2456 2144
rect 2474 2130 2490 2132
rect 2562 2130 2615 2144
rect 2563 2128 2627 2130
rect 2670 2128 2685 2144
rect 2734 2141 2764 2144
rect 2734 2138 2770 2141
rect 2700 2130 2716 2132
rect 2474 2118 2489 2122
rect 2392 2116 2489 2118
rect 2517 2116 2685 2128
rect 2701 2118 2716 2122
rect 2734 2119 2773 2138
rect 2792 2132 2799 2133
rect 2798 2125 2799 2132
rect 2782 2122 2783 2125
rect 2798 2122 2811 2125
rect 2734 2118 2764 2119
rect 2773 2118 2779 2119
rect 2782 2118 2811 2122
rect 2701 2117 2811 2118
rect 2701 2116 2817 2117
rect 2376 2108 2427 2116
rect 2376 2096 2401 2108
rect 2408 2096 2427 2108
rect 2458 2108 2508 2116
rect 2458 2100 2474 2108
rect 2481 2106 2508 2108
rect 2517 2106 2738 2116
rect 2481 2096 2738 2106
rect 2767 2108 2817 2116
rect 2767 2099 2783 2108
rect 2376 2088 2427 2096
rect 2474 2088 2738 2096
rect 2764 2096 2783 2099
rect 2790 2096 2817 2108
rect 2764 2088 2817 2096
rect 2392 2080 2393 2088
rect 2408 2080 2421 2088
rect 2392 2072 2408 2080
rect 2389 2065 2408 2068
rect 2389 2056 2411 2065
rect 2362 2046 2411 2056
rect 2362 2040 2392 2046
rect 2411 2041 2416 2046
rect 2334 2024 2408 2040
rect 2426 2032 2456 2088
rect 2491 2078 2699 2088
rect 2734 2084 2779 2088
rect 2782 2087 2783 2088
rect 2798 2087 2811 2088
rect 2517 2048 2706 2078
rect 2532 2045 2706 2048
rect 2525 2042 2706 2045
rect 2334 2022 2347 2024
rect 2362 2022 2396 2024
rect 2334 2006 2408 2022
rect 2435 2018 2448 2032
rect 2463 2018 2479 2034
rect 2525 2029 2536 2042
rect 2318 1984 2319 2000
rect 2334 1984 2347 2006
rect 2362 1984 2392 2006
rect 2435 2002 2497 2018
rect 2525 2011 2536 2027
rect 2541 2022 2551 2042
rect 2561 2022 2575 2042
rect 2578 2029 2587 2042
rect 2603 2029 2612 2042
rect 2541 2011 2575 2022
rect 2578 2011 2587 2027
rect 2603 2011 2612 2027
rect 2619 2022 2629 2042
rect 2639 2022 2653 2042
rect 2654 2029 2665 2042
rect 2619 2011 2653 2022
rect 2654 2011 2665 2027
rect 2711 2018 2727 2034
rect 2734 2032 2764 2084
rect 2798 2080 2799 2087
rect 2783 2072 2799 2080
rect 2770 2040 2783 2059
rect 2798 2040 2828 2056
rect 2770 2024 2844 2040
rect 2770 2022 2783 2024
rect 2798 2022 2832 2024
rect 2435 2000 2448 2002
rect 2463 2000 2497 2002
rect 2435 1984 2497 2000
rect 2541 1995 2557 1998
rect 2619 1995 2649 2006
rect 2697 2002 2743 2018
rect 2770 2006 2844 2022
rect 2697 2000 2731 2002
rect 2696 1984 2743 2000
rect 2770 1984 2783 2006
rect 2798 1984 2828 2006
rect 2855 1984 2856 2000
rect 2871 1984 2884 2144
rect 2914 2040 2927 2144
rect 2972 2122 2973 2132
rect 2988 2122 3001 2132
rect 2972 2118 3001 2122
rect 3006 2118 3036 2144
rect 3054 2130 3070 2132
rect 3142 2130 3195 2144
rect 3143 2128 3205 2130
rect 3250 2128 3265 2144
rect 3314 2141 3344 2144
rect 3314 2138 3350 2141
rect 3280 2130 3296 2132
rect 3054 2118 3069 2122
rect 2972 2116 3069 2118
rect 3097 2116 3265 2128
rect 3281 2118 3296 2122
rect 3314 2119 3353 2138
rect 3372 2132 3379 2133
rect 3378 2125 3379 2132
rect 3362 2122 3363 2125
rect 3378 2122 3391 2125
rect 3314 2118 3344 2119
rect 3353 2118 3359 2119
rect 3362 2118 3391 2122
rect 3281 2117 3391 2118
rect 3281 2116 3397 2117
rect 2956 2108 3007 2116
rect 2956 2096 2981 2108
rect 2988 2096 3007 2108
rect 3038 2108 3088 2116
rect 3038 2100 3054 2108
rect 3061 2106 3088 2108
rect 3097 2106 3318 2116
rect 3061 2096 3318 2106
rect 3347 2108 3397 2116
rect 3347 2099 3363 2108
rect 2956 2088 3007 2096
rect 3054 2088 3318 2096
rect 3344 2096 3363 2099
rect 3370 2096 3397 2108
rect 3344 2088 3397 2096
rect 2972 2080 2973 2088
rect 2988 2080 3001 2088
rect 2972 2072 2988 2080
rect 2969 2065 2988 2068
rect 2969 2056 2991 2065
rect 2942 2046 2991 2056
rect 2942 2040 2972 2046
rect 2991 2041 2996 2046
rect 2914 2024 2988 2040
rect 3006 2032 3036 2088
rect 3071 2078 3279 2088
rect 3314 2084 3359 2088
rect 3362 2087 3363 2088
rect 3378 2087 3391 2088
rect 3097 2048 3286 2078
rect 3112 2045 3286 2048
rect 3105 2042 3286 2045
rect 2914 2022 2927 2024
rect 2942 2022 2976 2024
rect 2914 2006 2988 2022
rect 3015 2018 3028 2032
rect 3043 2018 3059 2034
rect 3105 2029 3116 2042
rect 2898 1984 2899 2000
rect 2914 1984 2927 2006
rect 2942 1984 2972 2006
rect 3015 2002 3077 2018
rect 3105 2011 3116 2027
rect 3121 2022 3131 2042
rect 3141 2022 3155 2042
rect 3158 2029 3167 2042
rect 3183 2029 3192 2042
rect 3121 2011 3155 2022
rect 3158 2011 3167 2027
rect 3183 2011 3192 2027
rect 3199 2022 3209 2042
rect 3219 2022 3233 2042
rect 3234 2029 3245 2042
rect 3199 2011 3233 2022
rect 3234 2011 3245 2027
rect 3291 2018 3307 2034
rect 3314 2032 3344 2084
rect 3378 2080 3379 2087
rect 3363 2072 3379 2080
rect 3350 2040 3363 2059
rect 3378 2040 3408 2056
rect 3350 2024 3424 2040
rect 3350 2022 3363 2024
rect 3378 2022 3412 2024
rect 3015 2000 3028 2002
rect 3043 2000 3077 2002
rect 3015 1984 3077 2000
rect 3121 1995 3137 1998
rect 3199 1995 3229 2006
rect 3277 2002 3323 2018
rect 3350 2006 3424 2022
rect 3277 2000 3311 2002
rect 3276 1984 3323 2000
rect 3350 1984 3363 2006
rect 3378 1984 3408 2006
rect 3435 1984 3436 2000
rect 3451 1984 3464 2144
rect 3494 2040 3507 2144
rect 3552 2122 3553 2132
rect 3568 2122 3581 2132
rect 3552 2118 3581 2122
rect 3586 2118 3616 2144
rect 3634 2130 3650 2132
rect 3722 2130 3775 2144
rect 3723 2128 3787 2130
rect 3830 2128 3845 2144
rect 3894 2141 3924 2144
rect 3894 2138 3930 2141
rect 3860 2130 3876 2132
rect 3634 2118 3649 2122
rect 3552 2116 3649 2118
rect 3677 2116 3845 2128
rect 3861 2118 3876 2122
rect 3894 2119 3933 2138
rect 3952 2132 3959 2133
rect 3958 2125 3959 2132
rect 3942 2122 3943 2125
rect 3958 2122 3971 2125
rect 3894 2118 3924 2119
rect 3933 2118 3939 2119
rect 3942 2118 3971 2122
rect 3861 2117 3971 2118
rect 3861 2116 3977 2117
rect 3536 2108 3587 2116
rect 3536 2096 3561 2108
rect 3568 2096 3587 2108
rect 3618 2108 3668 2116
rect 3618 2100 3634 2108
rect 3641 2106 3668 2108
rect 3677 2106 3898 2116
rect 3641 2096 3898 2106
rect 3927 2108 3977 2116
rect 3927 2099 3943 2108
rect 3536 2088 3587 2096
rect 3634 2088 3898 2096
rect 3924 2096 3943 2099
rect 3950 2096 3977 2108
rect 3924 2088 3977 2096
rect 3552 2080 3553 2088
rect 3568 2080 3581 2088
rect 3552 2072 3568 2080
rect 3549 2065 3568 2068
rect 3549 2056 3571 2065
rect 3522 2046 3571 2056
rect 3522 2040 3552 2046
rect 3571 2041 3576 2046
rect 3494 2024 3568 2040
rect 3586 2032 3616 2088
rect 3651 2078 3859 2088
rect 3894 2084 3939 2088
rect 3942 2087 3943 2088
rect 3958 2087 3971 2088
rect 3677 2048 3866 2078
rect 3692 2045 3866 2048
rect 3685 2042 3866 2045
rect 3494 2022 3507 2024
rect 3522 2022 3556 2024
rect 3494 2006 3568 2022
rect 3595 2018 3608 2032
rect 3623 2018 3639 2034
rect 3685 2029 3696 2042
rect 3478 1984 3479 2000
rect 3494 1984 3507 2006
rect 3522 1984 3552 2006
rect 3595 2002 3657 2018
rect 3685 2011 3696 2027
rect 3701 2022 3711 2042
rect 3721 2022 3735 2042
rect 3738 2029 3747 2042
rect 3763 2029 3772 2042
rect 3701 2011 3735 2022
rect 3738 2011 3747 2027
rect 3763 2011 3772 2027
rect 3779 2022 3789 2042
rect 3799 2022 3813 2042
rect 3814 2029 3825 2042
rect 3779 2011 3813 2022
rect 3814 2011 3825 2027
rect 3871 2018 3887 2034
rect 3894 2032 3924 2084
rect 3958 2080 3959 2087
rect 3943 2072 3959 2080
rect 3930 2040 3943 2059
rect 3958 2040 3988 2056
rect 3930 2024 4004 2040
rect 3930 2022 3943 2024
rect 3958 2022 3992 2024
rect 3595 2000 3608 2002
rect 3623 2000 3657 2002
rect 3595 1984 3657 2000
rect 3701 1995 3717 1998
rect 3779 1995 3809 2006
rect 3857 2002 3903 2018
rect 3930 2006 4004 2022
rect 3857 2000 3891 2002
rect 3856 1984 3903 2000
rect 3930 1984 3943 2006
rect 3958 1984 3988 2006
rect 4015 1984 4016 2000
rect 4031 1984 4044 2144
rect 4074 2040 4087 2144
rect 4132 2122 4133 2132
rect 4148 2122 4161 2132
rect 4132 2118 4161 2122
rect 4166 2118 4196 2144
rect 4214 2130 4230 2132
rect 4302 2130 4355 2144
rect 4303 2128 4367 2130
rect 4410 2128 4425 2144
rect 4474 2141 4504 2144
rect 4474 2138 4510 2141
rect 4440 2130 4456 2132
rect 4214 2118 4229 2122
rect 4132 2116 4229 2118
rect 4257 2116 4425 2128
rect 4441 2118 4456 2122
rect 4474 2119 4513 2138
rect 4532 2132 4539 2133
rect 4538 2125 4539 2132
rect 4522 2122 4523 2125
rect 4538 2122 4551 2125
rect 4474 2118 4504 2119
rect 4513 2118 4519 2119
rect 4522 2118 4551 2122
rect 4441 2117 4551 2118
rect 4441 2116 4557 2117
rect 4116 2108 4167 2116
rect 4116 2096 4141 2108
rect 4148 2096 4167 2108
rect 4198 2108 4248 2116
rect 4198 2100 4214 2108
rect 4221 2106 4248 2108
rect 4257 2106 4478 2116
rect 4221 2096 4478 2106
rect 4507 2108 4557 2116
rect 4507 2099 4523 2108
rect 4116 2088 4167 2096
rect 4214 2088 4478 2096
rect 4504 2096 4523 2099
rect 4530 2096 4557 2108
rect 4504 2088 4557 2096
rect 4132 2080 4133 2088
rect 4148 2080 4161 2088
rect 4132 2072 4148 2080
rect 4129 2065 4148 2068
rect 4129 2056 4151 2065
rect 4102 2046 4151 2056
rect 4102 2040 4132 2046
rect 4151 2041 4156 2046
rect 4074 2024 4148 2040
rect 4166 2032 4196 2088
rect 4231 2078 4439 2088
rect 4474 2084 4519 2088
rect 4522 2087 4523 2088
rect 4538 2087 4551 2088
rect 4257 2048 4446 2078
rect 4272 2045 4446 2048
rect 4265 2042 4446 2045
rect 4074 2022 4087 2024
rect 4102 2022 4136 2024
rect 4074 2006 4148 2022
rect 4175 2018 4188 2032
rect 4203 2018 4219 2034
rect 4265 2029 4276 2042
rect 4058 1984 4059 2000
rect 4074 1984 4087 2006
rect 4102 1984 4132 2006
rect 4175 2002 4237 2018
rect 4265 2011 4276 2027
rect 4281 2022 4291 2042
rect 4301 2022 4315 2042
rect 4318 2029 4327 2042
rect 4343 2029 4352 2042
rect 4281 2011 4315 2022
rect 4318 2011 4327 2027
rect 4343 2011 4352 2027
rect 4359 2022 4369 2042
rect 4379 2022 4393 2042
rect 4394 2029 4405 2042
rect 4359 2011 4393 2022
rect 4394 2011 4405 2027
rect 4451 2018 4467 2034
rect 4474 2032 4504 2084
rect 4538 2080 4539 2087
rect 4523 2072 4539 2080
rect 4510 2040 4523 2059
rect 4538 2040 4568 2056
rect 4510 2024 4584 2040
rect 4510 2022 4523 2024
rect 4538 2022 4572 2024
rect 4175 2000 4188 2002
rect 4203 2000 4237 2002
rect 4175 1984 4237 2000
rect 4281 1995 4297 1998
rect 4359 1995 4389 2006
rect 4437 2002 4483 2018
rect 4510 2006 4584 2022
rect 4437 2000 4471 2002
rect 4436 1984 4483 2000
rect 4510 1984 4523 2006
rect 4538 1984 4568 2006
rect 4595 1984 4596 2000
rect 4611 1984 4624 2144
rect 4654 2040 4667 2144
rect 4712 2122 4713 2132
rect 4733 2130 4741 2132
rect 4731 2128 4741 2130
rect 4728 2122 4741 2128
rect 4712 2118 4741 2122
rect 4746 2118 4776 2144
rect 4794 2130 4810 2132
rect 4882 2130 4933 2144
rect 4883 2128 4947 2130
rect 4990 2128 5005 2144
rect 5054 2141 5084 2144
rect 5054 2138 5090 2141
rect 5020 2130 5036 2132
rect 4794 2118 4809 2122
rect 4712 2116 4809 2118
rect 4837 2116 5005 2128
rect 5021 2118 5036 2122
rect 5054 2119 5093 2138
rect 5112 2132 5119 2133
rect 5118 2125 5119 2132
rect 5102 2122 5103 2125
rect 5118 2122 5131 2125
rect 5054 2118 5084 2119
rect 5093 2118 5099 2119
rect 5102 2118 5131 2122
rect 5021 2117 5131 2118
rect 5021 2116 5137 2117
rect 4696 2108 4747 2116
rect 4696 2096 4721 2108
rect 4728 2096 4747 2108
rect 4778 2108 4828 2116
rect 4778 2100 4794 2108
rect 4801 2106 4828 2108
rect 4837 2106 5058 2116
rect 4801 2096 5058 2106
rect 5087 2108 5137 2116
rect 5087 2099 5103 2108
rect 4696 2088 4747 2096
rect 4794 2088 5058 2096
rect 5084 2096 5103 2099
rect 5110 2096 5137 2108
rect 5084 2088 5137 2096
rect 4712 2080 4713 2088
rect 4728 2080 4741 2088
rect 4712 2072 4728 2080
rect 4709 2065 4728 2068
rect 4709 2056 4731 2065
rect 4682 2046 4731 2056
rect 4682 2040 4712 2046
rect 4731 2041 4736 2046
rect 4654 2024 4728 2040
rect 4746 2032 4776 2088
rect 4811 2078 5019 2088
rect 5054 2084 5099 2088
rect 5102 2087 5103 2088
rect 5118 2087 5131 2088
rect 4837 2048 5026 2078
rect 4852 2045 5026 2048
rect 4845 2042 5026 2045
rect 4654 2022 4667 2024
rect 4682 2022 4716 2024
rect 4654 2006 4728 2022
rect 4755 2018 4768 2032
rect 4783 2018 4799 2034
rect 4845 2029 4856 2042
rect 4638 1984 4639 2000
rect 4654 1984 4667 2006
rect 4682 1984 4712 2006
rect 4755 2002 4817 2018
rect 4845 2011 4856 2027
rect 4861 2022 4871 2042
rect 4881 2022 4895 2042
rect 4898 2029 4907 2042
rect 4923 2029 4932 2042
rect 4861 2011 4895 2022
rect 4898 2011 4907 2027
rect 4923 2011 4932 2027
rect 4939 2022 4949 2042
rect 4959 2022 4973 2042
rect 4974 2029 4985 2042
rect 4939 2011 4973 2022
rect 4974 2011 4985 2027
rect 5031 2018 5047 2034
rect 5054 2032 5084 2084
rect 5118 2080 5119 2087
rect 5103 2072 5119 2080
rect 5090 2040 5103 2059
rect 5118 2040 5148 2056
rect 5090 2024 5164 2040
rect 5090 2022 5103 2024
rect 5118 2022 5152 2024
rect 4755 2000 4768 2002
rect 4783 2000 4817 2002
rect 4755 1984 4817 2000
rect 4861 1995 4877 1998
rect 4939 1995 4969 2006
rect 5017 2002 5063 2018
rect 5090 2006 5164 2022
rect 5017 2000 5051 2002
rect 5016 1984 5063 2000
rect 5090 1984 5103 2006
rect 5118 1984 5148 2006
rect 5175 1984 5176 2000
rect 5191 1984 5204 2144
rect 5234 2040 5247 2144
rect 5292 2122 5293 2132
rect 5313 2130 5321 2132
rect 5311 2128 5321 2130
rect 5308 2122 5321 2128
rect 5292 2118 5321 2122
rect 5326 2118 5356 2144
rect 5374 2130 5390 2132
rect 5462 2130 5513 2144
rect 5463 2128 5527 2130
rect 5570 2128 5585 2144
rect 5634 2141 5664 2144
rect 5634 2138 5670 2141
rect 5600 2130 5616 2132
rect 5374 2118 5389 2122
rect 5292 2116 5389 2118
rect 5417 2116 5585 2128
rect 5601 2118 5616 2122
rect 5634 2119 5673 2138
rect 5692 2132 5699 2133
rect 5698 2125 5699 2132
rect 5682 2122 5683 2125
rect 5698 2122 5711 2125
rect 5634 2118 5664 2119
rect 5673 2118 5679 2119
rect 5682 2118 5711 2122
rect 5601 2117 5711 2118
rect 5601 2116 5717 2117
rect 5276 2108 5327 2116
rect 5276 2096 5301 2108
rect 5308 2096 5327 2108
rect 5358 2108 5408 2116
rect 5358 2100 5374 2108
rect 5381 2106 5408 2108
rect 5417 2106 5638 2116
rect 5381 2096 5638 2106
rect 5667 2108 5717 2116
rect 5667 2099 5683 2108
rect 5276 2088 5327 2096
rect 5374 2088 5638 2096
rect 5664 2096 5683 2099
rect 5690 2096 5717 2108
rect 5664 2088 5717 2096
rect 5292 2080 5293 2088
rect 5308 2080 5321 2088
rect 5292 2072 5308 2080
rect 5289 2065 5308 2068
rect 5289 2056 5311 2065
rect 5262 2046 5311 2056
rect 5262 2040 5292 2046
rect 5311 2041 5316 2046
rect 5234 2024 5308 2040
rect 5326 2032 5356 2088
rect 5391 2078 5599 2088
rect 5634 2084 5679 2088
rect 5682 2087 5683 2088
rect 5698 2087 5711 2088
rect 5417 2048 5606 2078
rect 5432 2045 5606 2048
rect 5425 2042 5606 2045
rect 5234 2022 5247 2024
rect 5262 2022 5296 2024
rect 5234 2006 5308 2022
rect 5335 2018 5348 2032
rect 5363 2018 5379 2034
rect 5425 2029 5436 2042
rect 5218 1984 5219 2000
rect 5234 1984 5247 2006
rect 5262 1984 5292 2006
rect 5335 2002 5397 2018
rect 5425 2011 5436 2027
rect 5441 2022 5451 2042
rect 5461 2022 5475 2042
rect 5478 2029 5487 2042
rect 5503 2029 5512 2042
rect 5441 2011 5475 2022
rect 5478 2011 5487 2027
rect 5503 2011 5512 2027
rect 5519 2022 5529 2042
rect 5539 2022 5553 2042
rect 5554 2029 5565 2042
rect 5519 2011 5553 2022
rect 5554 2011 5565 2027
rect 5611 2018 5627 2034
rect 5634 2032 5664 2084
rect 5698 2080 5699 2087
rect 5683 2072 5699 2080
rect 5670 2040 5683 2059
rect 5698 2040 5728 2056
rect 5670 2024 5744 2040
rect 5670 2022 5683 2024
rect 5698 2022 5732 2024
rect 5335 2000 5348 2002
rect 5363 2000 5397 2002
rect 5335 1984 5397 2000
rect 5441 1995 5457 1998
rect 5519 1995 5549 2006
rect 5597 2002 5643 2018
rect 5670 2006 5744 2022
rect 5597 2000 5631 2002
rect 5596 1984 5643 2000
rect 5670 1984 5683 2006
rect 5698 1984 5728 2006
rect 5755 1984 5756 2000
rect 5771 1984 5784 2144
rect 5814 2040 5827 2144
rect 5872 2122 5873 2132
rect 5893 2130 5901 2132
rect 5891 2128 5901 2130
rect 5888 2122 5901 2128
rect 5872 2118 5901 2122
rect 5906 2118 5936 2144
rect 5954 2130 5970 2132
rect 6042 2130 6093 2144
rect 6043 2128 6107 2130
rect 6150 2128 6165 2144
rect 6214 2141 6244 2144
rect 6214 2138 6250 2141
rect 6180 2130 6196 2132
rect 5954 2118 5969 2122
rect 5872 2116 5969 2118
rect 5997 2116 6165 2128
rect 6181 2118 6196 2122
rect 6214 2119 6253 2138
rect 6272 2132 6279 2133
rect 6278 2125 6279 2132
rect 6262 2122 6263 2125
rect 6278 2122 6291 2125
rect 6214 2118 6244 2119
rect 6253 2118 6259 2119
rect 6262 2118 6291 2122
rect 6181 2117 6291 2118
rect 6181 2116 6297 2117
rect 5856 2108 5907 2116
rect 5856 2096 5881 2108
rect 5888 2096 5907 2108
rect 5938 2108 5988 2116
rect 5938 2100 5954 2108
rect 5961 2106 5988 2108
rect 5997 2106 6218 2116
rect 5961 2096 6218 2106
rect 6247 2108 6297 2116
rect 6247 2099 6263 2108
rect 5856 2088 5907 2096
rect 5954 2088 6218 2096
rect 6244 2096 6263 2099
rect 6270 2096 6297 2108
rect 6244 2088 6297 2096
rect 5872 2080 5873 2088
rect 5888 2080 5901 2088
rect 5872 2072 5888 2080
rect 5869 2065 5888 2068
rect 5869 2056 5891 2065
rect 5842 2046 5891 2056
rect 5842 2040 5872 2046
rect 5891 2041 5896 2046
rect 5814 2024 5888 2040
rect 5906 2032 5936 2088
rect 5971 2078 6179 2088
rect 6214 2084 6259 2088
rect 6262 2087 6263 2088
rect 6278 2087 6291 2088
rect 5997 2048 6186 2078
rect 6012 2045 6186 2048
rect 6005 2042 6186 2045
rect 5814 2022 5827 2024
rect 5842 2022 5876 2024
rect 5814 2006 5888 2022
rect 5915 2018 5928 2032
rect 5943 2018 5959 2034
rect 6005 2029 6016 2042
rect 5798 1984 5799 2000
rect 5814 1984 5827 2006
rect 5842 1984 5872 2006
rect 5915 2002 5977 2018
rect 6005 2011 6016 2027
rect 6021 2022 6031 2042
rect 6041 2022 6055 2042
rect 6058 2029 6067 2042
rect 6083 2029 6092 2042
rect 6021 2011 6055 2022
rect 6058 2011 6067 2027
rect 6083 2011 6092 2027
rect 6099 2022 6109 2042
rect 6119 2022 6133 2042
rect 6134 2029 6145 2042
rect 6099 2011 6133 2022
rect 6134 2011 6145 2027
rect 6191 2018 6207 2034
rect 6214 2032 6244 2084
rect 6278 2080 6279 2087
rect 6263 2072 6279 2080
rect 6250 2040 6263 2059
rect 6278 2040 6308 2056
rect 6250 2024 6324 2040
rect 6250 2022 6263 2024
rect 6278 2022 6312 2024
rect 5915 2000 5928 2002
rect 5943 2000 5977 2002
rect 5915 1984 5977 2000
rect 6021 1995 6037 1998
rect 6099 1995 6129 2006
rect 6177 2002 6223 2018
rect 6250 2006 6324 2022
rect 6177 2000 6211 2002
rect 6176 1984 6223 2000
rect 6250 1984 6263 2006
rect 6278 1984 6308 2006
rect 6335 1984 6336 2000
rect 6351 1984 6364 2144
rect 6394 2040 6407 2144
rect 6452 2122 6453 2132
rect 6473 2130 6481 2132
rect 6471 2128 6481 2130
rect 6468 2122 6481 2128
rect 6452 2118 6481 2122
rect 6486 2118 6516 2144
rect 6534 2130 6550 2132
rect 6622 2130 6673 2144
rect 6623 2128 6687 2130
rect 6730 2128 6745 2144
rect 6794 2141 6824 2144
rect 6794 2138 6830 2141
rect 6760 2130 6776 2132
rect 6534 2118 6549 2122
rect 6452 2116 6549 2118
rect 6577 2116 6745 2128
rect 6761 2118 6776 2122
rect 6794 2119 6833 2138
rect 6852 2132 6859 2133
rect 6858 2125 6859 2132
rect 6842 2122 6843 2125
rect 6858 2122 6871 2125
rect 6794 2118 6824 2119
rect 6833 2118 6839 2119
rect 6842 2118 6871 2122
rect 6761 2117 6871 2118
rect 6761 2116 6877 2117
rect 6436 2108 6487 2116
rect 6436 2096 6461 2108
rect 6468 2096 6487 2108
rect 6518 2108 6568 2116
rect 6518 2100 6534 2108
rect 6541 2106 6568 2108
rect 6577 2106 6798 2116
rect 6541 2096 6798 2106
rect 6827 2108 6877 2116
rect 6827 2099 6843 2108
rect 6436 2088 6487 2096
rect 6534 2088 6798 2096
rect 6824 2096 6843 2099
rect 6850 2096 6877 2108
rect 6824 2088 6877 2096
rect 6452 2080 6453 2088
rect 6468 2080 6481 2088
rect 6452 2072 6468 2080
rect 6449 2065 6468 2068
rect 6449 2056 6471 2065
rect 6422 2046 6471 2056
rect 6422 2040 6452 2046
rect 6471 2041 6476 2046
rect 6394 2024 6468 2040
rect 6486 2032 6516 2088
rect 6551 2078 6759 2088
rect 6794 2084 6839 2088
rect 6842 2087 6843 2088
rect 6858 2087 6871 2088
rect 6577 2048 6766 2078
rect 6592 2045 6766 2048
rect 6585 2042 6766 2045
rect 6394 2022 6407 2024
rect 6422 2022 6456 2024
rect 6394 2006 6468 2022
rect 6495 2018 6508 2032
rect 6523 2018 6539 2034
rect 6585 2029 6596 2042
rect 6378 1984 6379 2000
rect 6394 1984 6407 2006
rect 6422 1984 6452 2006
rect 6495 2002 6557 2018
rect 6585 2011 6596 2027
rect 6601 2022 6611 2042
rect 6621 2022 6635 2042
rect 6638 2029 6647 2042
rect 6663 2029 6672 2042
rect 6601 2011 6635 2022
rect 6638 2011 6647 2027
rect 6663 2011 6672 2027
rect 6679 2022 6689 2042
rect 6699 2022 6713 2042
rect 6714 2029 6725 2042
rect 6679 2011 6713 2022
rect 6714 2011 6725 2027
rect 6771 2018 6787 2034
rect 6794 2032 6824 2084
rect 6858 2080 6859 2087
rect 6843 2072 6859 2080
rect 6830 2040 6843 2059
rect 6858 2040 6888 2056
rect 6830 2024 6904 2040
rect 6830 2022 6843 2024
rect 6858 2022 6892 2024
rect 6495 2000 6508 2002
rect 6523 2000 6557 2002
rect 6495 1984 6557 2000
rect 6601 1995 6617 1998
rect 6679 1995 6709 2006
rect 6757 2002 6803 2018
rect 6830 2006 6904 2022
rect 6757 2000 6791 2002
rect 6756 1984 6803 2000
rect 6830 1984 6843 2006
rect 6858 1984 6888 2006
rect 6915 1984 6916 2000
rect 6931 1984 6944 2144
rect 0 1976 33 1984
rect 0 1950 7 1976
rect 14 1950 33 1976
rect 97 1972 159 1984
rect 171 1972 246 1984
rect 304 1972 379 1984
rect 391 1972 422 1984
rect 428 1972 463 1984
rect 97 1970 259 1972
rect 0 1942 33 1950
rect 115 1946 128 1970
rect 143 1968 158 1970
rect 14 1932 27 1942
rect 42 1932 72 1946
rect 115 1932 158 1946
rect 182 1943 189 1950
rect 192 1946 259 1970
rect 291 1970 463 1972
rect 261 1948 289 1952
rect 291 1948 371 1970
rect 392 1968 407 1970
rect 261 1946 371 1948
rect 192 1942 371 1946
rect 165 1932 195 1942
rect 197 1932 350 1942
rect 358 1932 388 1942
rect 392 1932 422 1946
rect 450 1932 463 1970
rect 535 1976 570 1984
rect 535 1950 536 1976
rect 543 1950 570 1976
rect 478 1932 508 1946
rect 535 1942 570 1950
rect 572 1976 613 1984
rect 572 1950 587 1976
rect 594 1950 613 1976
rect 677 1972 739 1984
rect 751 1972 826 1984
rect 884 1972 959 1984
rect 971 1972 1002 1984
rect 1008 1972 1043 1984
rect 677 1970 839 1972
rect 572 1942 613 1950
rect 695 1946 708 1970
rect 723 1968 738 1970
rect 535 1932 536 1942
rect 551 1932 564 1942
rect 578 1932 579 1942
rect 594 1932 607 1942
rect 622 1932 652 1946
rect 695 1932 738 1946
rect 762 1943 769 1950
rect 772 1946 839 1970
rect 871 1970 1043 1972
rect 841 1948 869 1952
rect 871 1948 951 1970
rect 972 1968 987 1970
rect 841 1946 951 1948
rect 772 1942 951 1946
rect 745 1932 775 1942
rect 777 1932 930 1942
rect 938 1932 968 1942
rect 972 1932 1002 1946
rect 1030 1932 1043 1970
rect 1115 1976 1150 1984
rect 1115 1950 1116 1976
rect 1123 1950 1150 1976
rect 1058 1932 1088 1946
rect 1115 1942 1150 1950
rect 1152 1976 1193 1984
rect 1152 1950 1167 1976
rect 1174 1950 1193 1976
rect 1257 1972 1319 1984
rect 1331 1972 1406 1984
rect 1464 1972 1539 1984
rect 1551 1972 1582 1984
rect 1588 1972 1623 1984
rect 1257 1970 1419 1972
rect 1152 1942 1193 1950
rect 1275 1946 1288 1970
rect 1303 1968 1318 1970
rect 1115 1932 1116 1942
rect 1131 1932 1144 1942
rect 1158 1932 1159 1942
rect 1174 1932 1187 1942
rect 1202 1932 1232 1946
rect 1275 1932 1318 1946
rect 1342 1943 1349 1950
rect 1352 1946 1419 1970
rect 1451 1970 1623 1972
rect 1421 1948 1449 1952
rect 1451 1948 1531 1970
rect 1552 1968 1567 1970
rect 1421 1946 1531 1948
rect 1352 1942 1531 1946
rect 1325 1932 1355 1942
rect 1357 1932 1510 1942
rect 1518 1932 1548 1942
rect 1552 1932 1582 1946
rect 1610 1932 1623 1970
rect 1695 1976 1730 1984
rect 1695 1950 1696 1976
rect 1703 1950 1730 1976
rect 1638 1932 1668 1946
rect 1695 1942 1730 1950
rect 1732 1976 1773 1984
rect 1732 1950 1747 1976
rect 1754 1950 1773 1976
rect 1837 1972 1899 1984
rect 1911 1972 1986 1984
rect 2044 1972 2119 1984
rect 2131 1972 2162 1984
rect 2168 1972 2203 1984
rect 1837 1970 1999 1972
rect 1732 1942 1773 1950
rect 1855 1946 1868 1970
rect 1883 1968 1898 1970
rect 1695 1932 1696 1942
rect 1711 1932 1724 1942
rect 1738 1932 1739 1942
rect 1754 1932 1767 1942
rect 1782 1932 1812 1946
rect 1855 1932 1898 1946
rect 1922 1943 1929 1950
rect 1932 1946 1999 1970
rect 2031 1970 2203 1972
rect 2001 1948 2029 1952
rect 2031 1948 2111 1970
rect 2132 1968 2147 1970
rect 2001 1946 2111 1948
rect 1932 1942 2111 1946
rect 1905 1932 1935 1942
rect 1937 1932 2090 1942
rect 2098 1932 2128 1942
rect 2132 1932 2162 1946
rect 2190 1932 2203 1970
rect 2275 1976 2310 1984
rect 2275 1950 2276 1976
rect 2283 1950 2310 1976
rect 2218 1932 2248 1946
rect 2275 1942 2310 1950
rect 2312 1976 2353 1984
rect 2312 1950 2327 1976
rect 2334 1950 2353 1976
rect 2417 1972 2479 1984
rect 2491 1972 2566 1984
rect 2624 1972 2699 1984
rect 2711 1972 2742 1984
rect 2748 1972 2783 1984
rect 2417 1970 2579 1972
rect 2312 1942 2353 1950
rect 2435 1946 2448 1970
rect 2463 1968 2478 1970
rect 2275 1932 2276 1942
rect 2291 1932 2304 1942
rect 2318 1932 2319 1942
rect 2334 1932 2347 1942
rect 2362 1932 2392 1946
rect 2435 1932 2478 1946
rect 2502 1943 2509 1950
rect 2512 1946 2579 1970
rect 2611 1970 2783 1972
rect 2581 1948 2609 1952
rect 2611 1948 2691 1970
rect 2712 1968 2727 1970
rect 2581 1946 2691 1948
rect 2512 1942 2691 1946
rect 2485 1932 2515 1942
rect 2517 1932 2670 1942
rect 2678 1932 2708 1942
rect 2712 1932 2742 1946
rect 2770 1932 2783 1970
rect 2855 1976 2890 1984
rect 2855 1950 2856 1976
rect 2863 1950 2890 1976
rect 2798 1932 2828 1946
rect 2855 1942 2890 1950
rect 2892 1976 2933 1984
rect 2892 1950 2907 1976
rect 2914 1950 2933 1976
rect 2997 1972 3059 1984
rect 3071 1972 3146 1984
rect 3204 1972 3279 1984
rect 3291 1972 3322 1984
rect 3328 1972 3363 1984
rect 2997 1970 3159 1972
rect 2892 1942 2933 1950
rect 3015 1946 3028 1970
rect 3043 1968 3058 1970
rect 2855 1932 2856 1942
rect 2871 1932 2884 1942
rect 2898 1932 2899 1942
rect 2914 1932 2927 1942
rect 2942 1932 2972 1946
rect 3015 1932 3058 1946
rect 3082 1943 3089 1950
rect 3092 1946 3159 1970
rect 3191 1970 3363 1972
rect 3161 1948 3189 1952
rect 3191 1948 3271 1970
rect 3292 1968 3307 1970
rect 3161 1946 3271 1948
rect 3092 1942 3271 1946
rect 3065 1932 3095 1942
rect 3097 1932 3250 1942
rect 3258 1932 3288 1942
rect 3292 1932 3322 1946
rect 3350 1932 3363 1970
rect 3435 1976 3470 1984
rect 3435 1950 3436 1976
rect 3443 1950 3470 1976
rect 3378 1932 3408 1946
rect 3435 1942 3470 1950
rect 3472 1976 3513 1984
rect 3472 1950 3487 1976
rect 3494 1950 3513 1976
rect 3577 1972 3639 1984
rect 3651 1972 3726 1984
rect 3784 1972 3859 1984
rect 3871 1972 3902 1984
rect 3908 1972 3943 1984
rect 3577 1970 3739 1972
rect 3472 1942 3513 1950
rect 3595 1946 3608 1970
rect 3623 1968 3638 1970
rect 3435 1932 3436 1942
rect 3451 1932 3464 1942
rect 3478 1932 3479 1942
rect 3494 1932 3507 1942
rect 3522 1932 3552 1946
rect 3595 1932 3638 1946
rect 3662 1943 3669 1950
rect 3672 1946 3739 1970
rect 3771 1970 3943 1972
rect 3741 1948 3769 1952
rect 3771 1948 3851 1970
rect 3872 1968 3887 1970
rect 3741 1946 3851 1948
rect 3672 1942 3851 1946
rect 3645 1932 3675 1942
rect 3677 1932 3830 1942
rect 3838 1932 3868 1942
rect 3872 1932 3902 1946
rect 3930 1932 3943 1970
rect 4015 1976 4050 1984
rect 4015 1950 4016 1976
rect 4023 1950 4050 1976
rect 3958 1932 3988 1946
rect 4015 1942 4050 1950
rect 4052 1976 4093 1984
rect 4052 1950 4067 1976
rect 4074 1950 4093 1976
rect 4157 1972 4219 1984
rect 4231 1972 4306 1984
rect 4364 1972 4439 1984
rect 4451 1972 4482 1984
rect 4488 1972 4523 1984
rect 4157 1970 4319 1972
rect 4052 1942 4093 1950
rect 4175 1946 4188 1970
rect 4203 1968 4218 1970
rect 4015 1932 4016 1942
rect 4031 1932 4044 1942
rect 4058 1932 4059 1942
rect 4074 1932 4087 1942
rect 4102 1932 4132 1946
rect 4175 1932 4218 1946
rect 4242 1943 4249 1950
rect 4252 1946 4319 1970
rect 4351 1970 4523 1972
rect 4321 1948 4349 1952
rect 4351 1948 4431 1970
rect 4452 1968 4467 1970
rect 4321 1946 4431 1948
rect 4252 1942 4431 1946
rect 4225 1932 4255 1942
rect 4257 1932 4410 1942
rect 4418 1932 4448 1942
rect 4452 1932 4482 1946
rect 4510 1932 4523 1970
rect 4595 1976 4630 1984
rect 4595 1950 4596 1976
rect 4603 1950 4630 1976
rect 4538 1932 4568 1946
rect 4595 1942 4630 1950
rect 4632 1976 4673 1984
rect 4632 1950 4647 1976
rect 4654 1950 4673 1976
rect 4737 1972 4799 1984
rect 4811 1972 4886 1984
rect 4944 1972 5019 1984
rect 5031 1972 5062 1984
rect 5068 1972 5103 1984
rect 4737 1970 4899 1972
rect 4632 1942 4673 1950
rect 4755 1946 4768 1970
rect 4783 1968 4798 1970
rect 4832 1952 4899 1970
rect 4931 1970 5103 1972
rect 4931 1952 5011 1970
rect 5032 1968 5047 1970
rect 4595 1932 4596 1942
rect 4611 1932 4624 1942
rect 4638 1932 4639 1942
rect 4654 1932 4667 1942
rect 4682 1932 4712 1946
rect 4755 1932 4798 1946
rect 4822 1943 4829 1950
rect 4832 1942 5011 1952
rect 4805 1932 4835 1942
rect 4837 1932 4990 1942
rect 4998 1932 5028 1942
rect 5032 1932 5062 1946
rect 5090 1932 5103 1970
rect 5175 1976 5210 1984
rect 5175 1950 5176 1976
rect 5183 1950 5210 1976
rect 5118 1932 5148 1946
rect 5175 1942 5210 1950
rect 5212 1976 5253 1984
rect 5212 1950 5227 1976
rect 5234 1950 5253 1976
rect 5317 1972 5379 1984
rect 5391 1972 5466 1984
rect 5524 1972 5599 1984
rect 5611 1972 5642 1984
rect 5648 1972 5683 1984
rect 5317 1970 5479 1972
rect 5212 1942 5253 1950
rect 5335 1946 5348 1970
rect 5363 1968 5378 1970
rect 5412 1952 5479 1970
rect 5511 1970 5683 1972
rect 5511 1952 5591 1970
rect 5612 1968 5627 1970
rect 5175 1932 5176 1942
rect 5191 1932 5204 1942
rect 5218 1932 5219 1942
rect 5234 1932 5247 1942
rect 5262 1932 5292 1946
rect 5335 1932 5378 1946
rect 5402 1943 5409 1950
rect 5412 1942 5591 1952
rect 5385 1932 5415 1942
rect 5417 1932 5570 1942
rect 5578 1932 5608 1942
rect 5612 1932 5642 1946
rect 5670 1932 5683 1970
rect 5755 1976 5790 1984
rect 5755 1950 5756 1976
rect 5763 1950 5790 1976
rect 5698 1932 5728 1946
rect 5755 1942 5790 1950
rect 5792 1976 5833 1984
rect 5792 1950 5807 1976
rect 5814 1950 5833 1976
rect 5897 1972 5959 1984
rect 5971 1972 6046 1984
rect 6104 1972 6179 1984
rect 6191 1972 6222 1984
rect 6228 1972 6263 1984
rect 5897 1970 6059 1972
rect 5792 1942 5833 1950
rect 5915 1946 5928 1970
rect 5943 1968 5958 1970
rect 5992 1952 6059 1970
rect 6091 1970 6263 1972
rect 6091 1952 6171 1970
rect 6192 1968 6207 1970
rect 5755 1932 5756 1942
rect 5771 1932 5784 1942
rect 5798 1932 5799 1942
rect 5814 1932 5827 1942
rect 5842 1932 5872 1946
rect 5915 1932 5958 1946
rect 5982 1943 5989 1950
rect 5992 1942 6171 1952
rect 5965 1932 5995 1942
rect 5997 1932 6150 1942
rect 6158 1932 6188 1942
rect 6192 1932 6222 1946
rect 6250 1932 6263 1970
rect 6335 1976 6370 1984
rect 6335 1950 6336 1976
rect 6343 1950 6370 1976
rect 6278 1932 6308 1946
rect 6335 1942 6370 1950
rect 6372 1976 6413 1984
rect 6372 1950 6387 1976
rect 6394 1950 6413 1976
rect 6477 1972 6539 1984
rect 6551 1972 6626 1984
rect 6684 1972 6759 1984
rect 6771 1972 6802 1984
rect 6808 1972 6843 1984
rect 6477 1970 6639 1972
rect 6372 1942 6413 1950
rect 6495 1946 6508 1970
rect 6523 1968 6538 1970
rect 6572 1952 6639 1970
rect 6671 1970 6843 1972
rect 6671 1952 6751 1970
rect 6772 1968 6787 1970
rect 6335 1932 6336 1942
rect 6351 1932 6364 1942
rect 6378 1932 6379 1942
rect 6394 1932 6407 1942
rect 6422 1932 6452 1946
rect 6495 1932 6538 1946
rect 6562 1943 6569 1950
rect 6572 1942 6751 1952
rect 6545 1932 6575 1942
rect 6577 1932 6730 1942
rect 6738 1932 6768 1942
rect 6772 1932 6802 1946
rect 6830 1932 6843 1970
rect 6915 1976 6950 1984
rect 6915 1950 6916 1976
rect 6923 1950 6950 1976
rect 6858 1932 6888 1946
rect 6915 1942 6950 1950
rect 6915 1932 6916 1942
rect 6931 1932 6944 1942
rect 0 1918 6944 1932
rect 14 1888 27 1918
rect 42 1900 72 1918
rect 115 1904 129 1918
rect 165 1904 385 1918
rect 116 1902 129 1904
rect 82 1890 97 1902
rect 79 1888 101 1890
rect 106 1888 136 1902
rect 197 1900 350 1904
rect 179 1888 371 1900
rect 414 1888 444 1902
rect 450 1888 463 1918
rect 478 1900 508 1918
rect 551 1888 564 1918
rect 594 1888 607 1918
rect 622 1900 652 1918
rect 695 1904 709 1918
rect 745 1904 965 1918
rect 696 1902 709 1904
rect 662 1890 677 1902
rect 659 1888 681 1890
rect 686 1888 716 1902
rect 777 1900 930 1904
rect 759 1888 951 1900
rect 994 1888 1024 1902
rect 1030 1888 1043 1918
rect 1058 1900 1088 1918
rect 1131 1888 1144 1918
rect 1174 1888 1187 1918
rect 1202 1900 1232 1918
rect 1275 1904 1289 1918
rect 1325 1904 1545 1918
rect 1276 1902 1289 1904
rect 1242 1890 1257 1902
rect 1239 1888 1261 1890
rect 1266 1888 1296 1902
rect 1357 1900 1510 1904
rect 1339 1888 1531 1900
rect 1574 1888 1604 1902
rect 1610 1888 1623 1918
rect 1638 1900 1668 1918
rect 1711 1888 1724 1918
rect 1754 1888 1767 1918
rect 1782 1900 1812 1918
rect 1855 1904 1869 1918
rect 1905 1904 2125 1918
rect 1856 1902 1869 1904
rect 1822 1890 1837 1902
rect 1819 1888 1841 1890
rect 1846 1888 1876 1902
rect 1937 1900 2090 1904
rect 1919 1888 2111 1900
rect 2154 1888 2184 1902
rect 2190 1888 2203 1918
rect 2218 1900 2248 1918
rect 2291 1888 2304 1918
rect 2334 1888 2347 1918
rect 2362 1900 2392 1918
rect 2435 1904 2449 1918
rect 2485 1904 2705 1918
rect 2436 1902 2449 1904
rect 2402 1890 2417 1902
rect 2399 1888 2421 1890
rect 2426 1888 2456 1902
rect 2517 1900 2670 1904
rect 2499 1888 2691 1900
rect 2734 1888 2764 1902
rect 2770 1888 2783 1918
rect 2798 1900 2828 1918
rect 2871 1888 2884 1918
rect 2914 1888 2927 1918
rect 2942 1900 2972 1918
rect 3015 1904 3029 1918
rect 3065 1904 3285 1918
rect 3016 1902 3029 1904
rect 2982 1890 2997 1902
rect 2979 1888 3001 1890
rect 3006 1888 3036 1902
rect 3097 1900 3250 1904
rect 3079 1888 3271 1900
rect 3314 1888 3344 1902
rect 3350 1888 3363 1918
rect 3378 1900 3408 1918
rect 3451 1888 3464 1918
rect 3494 1888 3507 1918
rect 3522 1900 3552 1918
rect 3595 1904 3609 1918
rect 3645 1904 3865 1918
rect 3596 1902 3609 1904
rect 3562 1890 3577 1902
rect 3559 1888 3581 1890
rect 3586 1888 3616 1902
rect 3677 1900 3830 1904
rect 3659 1888 3851 1900
rect 3894 1888 3924 1902
rect 3930 1888 3943 1918
rect 3958 1900 3988 1918
rect 4031 1888 4044 1918
rect 4074 1888 4087 1918
rect 4102 1900 4132 1918
rect 4175 1904 4189 1918
rect 4225 1904 4445 1918
rect 4176 1902 4189 1904
rect 4142 1890 4157 1902
rect 4139 1888 4161 1890
rect 4166 1888 4196 1902
rect 4257 1900 4410 1904
rect 4239 1888 4431 1900
rect 4474 1888 4504 1902
rect 4510 1888 4523 1918
rect 4538 1900 4568 1918
rect 4611 1888 4624 1918
rect 4654 1888 4667 1918
rect 4682 1900 4712 1918
rect 4755 1904 4769 1918
rect 4805 1904 5025 1918
rect 4756 1902 4769 1904
rect 4722 1890 4737 1902
rect 4719 1888 4741 1890
rect 4746 1888 4776 1902
rect 4837 1900 4990 1904
rect 4819 1888 5011 1900
rect 5054 1888 5084 1902
rect 5090 1888 5103 1918
rect 5118 1900 5148 1918
rect 5191 1888 5204 1918
rect 5234 1888 5247 1918
rect 5262 1900 5292 1918
rect 5335 1904 5349 1918
rect 5385 1904 5605 1918
rect 5336 1902 5349 1904
rect 5302 1890 5317 1902
rect 5299 1888 5321 1890
rect 5326 1888 5356 1902
rect 5417 1900 5570 1904
rect 5399 1888 5591 1900
rect 5634 1888 5664 1902
rect 5670 1888 5683 1918
rect 5698 1900 5728 1918
rect 5771 1888 5784 1918
rect 5814 1888 5827 1918
rect 5842 1900 5872 1918
rect 5915 1904 5929 1918
rect 5965 1904 6185 1918
rect 5916 1902 5929 1904
rect 5882 1890 5897 1902
rect 5879 1888 5901 1890
rect 5906 1888 5936 1902
rect 5997 1900 6150 1904
rect 5979 1888 6171 1900
rect 6214 1888 6244 1902
rect 6250 1888 6263 1918
rect 6278 1900 6308 1918
rect 6351 1888 6364 1918
rect 6394 1888 6407 1918
rect 6422 1900 6452 1918
rect 6495 1904 6509 1918
rect 6545 1904 6765 1918
rect 6496 1902 6509 1904
rect 6462 1890 6477 1902
rect 6459 1888 6481 1890
rect 6486 1888 6516 1902
rect 6577 1900 6730 1904
rect 6559 1888 6751 1900
rect 6794 1888 6824 1902
rect 6830 1888 6843 1918
rect 6858 1900 6888 1918
rect 6931 1888 6944 1918
rect 0 1874 6944 1888
rect 14 1770 27 1874
rect 72 1852 73 1862
rect 88 1852 101 1862
rect 72 1848 101 1852
rect 106 1848 136 1874
rect 154 1860 170 1862
rect 242 1860 295 1874
rect 243 1858 307 1860
rect 350 1858 365 1874
rect 414 1871 444 1874
rect 414 1868 450 1871
rect 380 1860 396 1862
rect 154 1848 169 1852
rect 72 1846 169 1848
rect 197 1846 365 1858
rect 381 1848 396 1852
rect 414 1849 453 1868
rect 472 1862 479 1863
rect 478 1855 479 1862
rect 462 1852 463 1855
rect 478 1852 491 1855
rect 414 1848 444 1849
rect 453 1848 459 1849
rect 462 1848 491 1852
rect 381 1847 491 1848
rect 381 1846 497 1847
rect 56 1838 107 1846
rect 56 1826 81 1838
rect 88 1826 107 1838
rect 138 1838 188 1846
rect 138 1830 154 1838
rect 161 1836 188 1838
rect 197 1836 418 1846
rect 161 1826 418 1836
rect 447 1838 497 1846
rect 447 1829 463 1838
rect 56 1818 107 1826
rect 154 1818 418 1826
rect 444 1826 463 1829
rect 470 1826 497 1838
rect 444 1818 497 1826
rect 72 1810 73 1818
rect 88 1810 101 1818
rect 72 1802 88 1810
rect 69 1795 88 1798
rect 69 1786 91 1795
rect 42 1776 91 1786
rect 42 1770 72 1776
rect 91 1771 96 1776
rect 14 1754 88 1770
rect 106 1762 136 1818
rect 171 1808 379 1818
rect 414 1814 459 1818
rect 462 1817 463 1818
rect 478 1817 491 1818
rect 197 1778 386 1808
rect 212 1775 386 1778
rect 205 1772 386 1775
rect 14 1752 27 1754
rect 42 1752 76 1754
rect 14 1736 88 1752
rect 115 1748 128 1762
rect 143 1748 159 1764
rect 205 1759 216 1772
rect 14 1714 27 1736
rect 42 1714 72 1736
rect 115 1732 177 1748
rect 205 1741 216 1757
rect 221 1752 231 1772
rect 241 1752 255 1772
rect 258 1759 267 1772
rect 283 1759 292 1772
rect 221 1741 255 1752
rect 258 1741 267 1757
rect 283 1741 292 1757
rect 299 1752 309 1772
rect 319 1752 333 1772
rect 334 1759 345 1772
rect 299 1741 333 1752
rect 334 1741 345 1757
rect 391 1748 407 1764
rect 414 1762 444 1814
rect 478 1810 479 1817
rect 463 1802 479 1810
rect 450 1770 463 1789
rect 478 1770 508 1786
rect 450 1754 524 1770
rect 450 1752 463 1754
rect 478 1752 512 1754
rect 115 1730 128 1732
rect 143 1730 177 1732
rect 115 1714 177 1730
rect 221 1725 237 1728
rect 299 1725 329 1736
rect 377 1732 423 1748
rect 450 1736 524 1752
rect 377 1730 411 1732
rect 376 1714 423 1730
rect 450 1714 463 1736
rect 478 1714 508 1736
rect 535 1714 536 1730
rect 551 1714 564 1874
rect 594 1770 607 1874
rect 652 1852 653 1862
rect 668 1852 681 1862
rect 652 1848 681 1852
rect 686 1848 716 1874
rect 734 1860 750 1862
rect 822 1860 875 1874
rect 823 1858 887 1860
rect 930 1858 945 1874
rect 994 1871 1024 1874
rect 994 1868 1030 1871
rect 960 1860 976 1862
rect 734 1848 749 1852
rect 652 1846 749 1848
rect 777 1846 945 1858
rect 961 1848 976 1852
rect 994 1849 1033 1868
rect 1052 1862 1059 1863
rect 1058 1855 1059 1862
rect 1042 1852 1043 1855
rect 1058 1852 1071 1855
rect 994 1848 1024 1849
rect 1033 1848 1039 1849
rect 1042 1848 1071 1852
rect 961 1847 1071 1848
rect 961 1846 1077 1847
rect 636 1838 687 1846
rect 636 1826 661 1838
rect 668 1826 687 1838
rect 718 1838 768 1846
rect 718 1830 734 1838
rect 741 1836 768 1838
rect 777 1836 998 1846
rect 741 1826 998 1836
rect 1027 1838 1077 1846
rect 1027 1829 1043 1838
rect 636 1818 687 1826
rect 734 1818 998 1826
rect 1024 1826 1043 1829
rect 1050 1826 1077 1838
rect 1024 1818 1077 1826
rect 652 1810 653 1818
rect 668 1810 681 1818
rect 652 1802 668 1810
rect 649 1795 668 1798
rect 649 1786 671 1795
rect 622 1776 671 1786
rect 622 1770 652 1776
rect 671 1771 676 1776
rect 594 1754 668 1770
rect 686 1762 716 1818
rect 751 1808 959 1818
rect 994 1814 1039 1818
rect 1042 1817 1043 1818
rect 1058 1817 1071 1818
rect 777 1778 966 1808
rect 792 1775 966 1778
rect 785 1772 966 1775
rect 594 1752 607 1754
rect 622 1752 656 1754
rect 594 1736 668 1752
rect 695 1748 708 1762
rect 723 1748 739 1764
rect 785 1759 796 1772
rect 578 1714 579 1730
rect 594 1714 607 1736
rect 622 1714 652 1736
rect 695 1732 757 1748
rect 785 1741 796 1757
rect 801 1752 811 1772
rect 821 1752 835 1772
rect 838 1759 847 1772
rect 863 1759 872 1772
rect 801 1741 835 1752
rect 838 1741 847 1757
rect 863 1741 872 1757
rect 879 1752 889 1772
rect 899 1752 913 1772
rect 914 1759 925 1772
rect 879 1741 913 1752
rect 914 1741 925 1757
rect 971 1748 987 1764
rect 994 1762 1024 1814
rect 1058 1810 1059 1817
rect 1043 1802 1059 1810
rect 1030 1770 1043 1789
rect 1058 1770 1088 1786
rect 1030 1754 1104 1770
rect 1030 1752 1043 1754
rect 1058 1752 1092 1754
rect 695 1730 708 1732
rect 723 1730 757 1732
rect 695 1714 757 1730
rect 801 1725 817 1728
rect 879 1725 909 1736
rect 957 1732 1003 1748
rect 1030 1736 1104 1752
rect 957 1730 991 1732
rect 956 1714 1003 1730
rect 1030 1714 1043 1736
rect 1058 1714 1088 1736
rect 1115 1714 1116 1730
rect 1131 1714 1144 1874
rect 1174 1770 1187 1874
rect 1232 1852 1233 1862
rect 1248 1852 1261 1862
rect 1232 1848 1261 1852
rect 1266 1848 1296 1874
rect 1314 1860 1330 1862
rect 1402 1860 1455 1874
rect 1403 1858 1467 1860
rect 1510 1858 1525 1874
rect 1574 1871 1604 1874
rect 1574 1868 1610 1871
rect 1540 1860 1556 1862
rect 1314 1848 1329 1852
rect 1232 1846 1329 1848
rect 1357 1846 1525 1858
rect 1541 1848 1556 1852
rect 1574 1849 1613 1868
rect 1632 1862 1639 1863
rect 1638 1855 1639 1862
rect 1622 1852 1623 1855
rect 1638 1852 1651 1855
rect 1574 1848 1604 1849
rect 1613 1848 1619 1849
rect 1622 1848 1651 1852
rect 1541 1847 1651 1848
rect 1541 1846 1657 1847
rect 1216 1838 1267 1846
rect 1216 1826 1241 1838
rect 1248 1826 1267 1838
rect 1298 1838 1348 1846
rect 1298 1830 1314 1838
rect 1321 1836 1348 1838
rect 1357 1836 1578 1846
rect 1321 1826 1578 1836
rect 1607 1838 1657 1846
rect 1607 1829 1623 1838
rect 1216 1818 1267 1826
rect 1314 1818 1578 1826
rect 1604 1826 1623 1829
rect 1630 1826 1657 1838
rect 1604 1818 1657 1826
rect 1232 1810 1233 1818
rect 1248 1810 1261 1818
rect 1232 1802 1248 1810
rect 1229 1795 1248 1798
rect 1229 1786 1251 1795
rect 1202 1776 1251 1786
rect 1202 1770 1232 1776
rect 1251 1771 1256 1776
rect 1174 1754 1248 1770
rect 1266 1762 1296 1818
rect 1331 1808 1539 1818
rect 1574 1814 1619 1818
rect 1622 1817 1623 1818
rect 1638 1817 1651 1818
rect 1357 1778 1546 1808
rect 1372 1775 1546 1778
rect 1365 1772 1546 1775
rect 1174 1752 1187 1754
rect 1202 1752 1236 1754
rect 1174 1736 1248 1752
rect 1275 1748 1288 1762
rect 1303 1748 1319 1764
rect 1365 1759 1376 1772
rect 1158 1714 1159 1730
rect 1174 1714 1187 1736
rect 1202 1714 1232 1736
rect 1275 1732 1337 1748
rect 1365 1741 1376 1757
rect 1381 1752 1391 1772
rect 1401 1752 1415 1772
rect 1418 1759 1427 1772
rect 1443 1759 1452 1772
rect 1381 1741 1415 1752
rect 1418 1741 1427 1757
rect 1443 1741 1452 1757
rect 1459 1752 1469 1772
rect 1479 1752 1493 1772
rect 1494 1759 1505 1772
rect 1459 1741 1493 1752
rect 1494 1741 1505 1757
rect 1551 1748 1567 1764
rect 1574 1762 1604 1814
rect 1638 1810 1639 1817
rect 1623 1802 1639 1810
rect 1610 1770 1623 1789
rect 1638 1770 1668 1786
rect 1610 1754 1684 1770
rect 1610 1752 1623 1754
rect 1638 1752 1672 1754
rect 1275 1730 1288 1732
rect 1303 1730 1337 1732
rect 1275 1714 1337 1730
rect 1381 1725 1397 1728
rect 1459 1725 1489 1736
rect 1537 1732 1583 1748
rect 1610 1736 1684 1752
rect 1537 1730 1571 1732
rect 1536 1714 1583 1730
rect 1610 1714 1623 1736
rect 1638 1714 1668 1736
rect 1695 1714 1696 1730
rect 1711 1714 1724 1874
rect 1754 1770 1767 1874
rect 1812 1852 1813 1862
rect 1828 1852 1841 1862
rect 1812 1848 1841 1852
rect 1846 1848 1876 1874
rect 1894 1860 1910 1862
rect 1982 1860 2035 1874
rect 1983 1858 2047 1860
rect 2090 1858 2105 1874
rect 2154 1871 2184 1874
rect 2154 1868 2190 1871
rect 2120 1860 2136 1862
rect 1894 1848 1909 1852
rect 1812 1846 1909 1848
rect 1937 1846 2105 1858
rect 2121 1848 2136 1852
rect 2154 1849 2193 1868
rect 2212 1862 2219 1863
rect 2218 1855 2219 1862
rect 2202 1852 2203 1855
rect 2218 1852 2231 1855
rect 2154 1848 2184 1849
rect 2193 1848 2199 1849
rect 2202 1848 2231 1852
rect 2121 1847 2231 1848
rect 2121 1846 2237 1847
rect 1796 1838 1847 1846
rect 1796 1826 1821 1838
rect 1828 1826 1847 1838
rect 1878 1838 1928 1846
rect 1878 1830 1894 1838
rect 1901 1836 1928 1838
rect 1937 1836 2158 1846
rect 1901 1826 2158 1836
rect 2187 1838 2237 1846
rect 2187 1829 2203 1838
rect 1796 1818 1847 1826
rect 1894 1818 2158 1826
rect 2184 1826 2203 1829
rect 2210 1826 2237 1838
rect 2184 1818 2237 1826
rect 1812 1810 1813 1818
rect 1828 1810 1841 1818
rect 1812 1802 1828 1810
rect 1809 1795 1828 1798
rect 1809 1786 1831 1795
rect 1782 1776 1831 1786
rect 1782 1770 1812 1776
rect 1831 1771 1836 1776
rect 1754 1754 1828 1770
rect 1846 1762 1876 1818
rect 1911 1808 2119 1818
rect 2154 1814 2199 1818
rect 2202 1817 2203 1818
rect 2218 1817 2231 1818
rect 1937 1778 2126 1808
rect 1952 1775 2126 1778
rect 1945 1772 2126 1775
rect 1754 1752 1767 1754
rect 1782 1752 1816 1754
rect 1754 1736 1828 1752
rect 1855 1748 1868 1762
rect 1883 1748 1899 1764
rect 1945 1759 1956 1772
rect 1738 1714 1739 1730
rect 1754 1714 1767 1736
rect 1782 1714 1812 1736
rect 1855 1732 1917 1748
rect 1945 1741 1956 1757
rect 1961 1752 1971 1772
rect 1981 1752 1995 1772
rect 1998 1759 2007 1772
rect 2023 1759 2032 1772
rect 1961 1741 1995 1752
rect 1998 1741 2007 1757
rect 2023 1741 2032 1757
rect 2039 1752 2049 1772
rect 2059 1752 2073 1772
rect 2074 1759 2085 1772
rect 2039 1741 2073 1752
rect 2074 1741 2085 1757
rect 2131 1748 2147 1764
rect 2154 1762 2184 1814
rect 2218 1810 2219 1817
rect 2203 1802 2219 1810
rect 2190 1770 2203 1789
rect 2218 1770 2248 1786
rect 2190 1754 2264 1770
rect 2190 1752 2203 1754
rect 2218 1752 2252 1754
rect 1855 1730 1868 1732
rect 1883 1730 1917 1732
rect 1855 1714 1917 1730
rect 1961 1725 1977 1728
rect 2039 1725 2069 1736
rect 2117 1732 2163 1748
rect 2190 1736 2264 1752
rect 2117 1730 2151 1732
rect 2116 1714 2163 1730
rect 2190 1714 2203 1736
rect 2218 1714 2248 1736
rect 2275 1714 2276 1730
rect 2291 1714 2304 1874
rect 2334 1770 2347 1874
rect 2392 1852 2393 1862
rect 2408 1852 2421 1862
rect 2392 1848 2421 1852
rect 2426 1848 2456 1874
rect 2474 1860 2490 1862
rect 2562 1860 2615 1874
rect 2563 1858 2627 1860
rect 2670 1858 2685 1874
rect 2734 1871 2764 1874
rect 2734 1868 2770 1871
rect 2700 1860 2716 1862
rect 2474 1848 2489 1852
rect 2392 1846 2489 1848
rect 2517 1846 2685 1858
rect 2701 1848 2716 1852
rect 2734 1849 2773 1868
rect 2792 1862 2799 1863
rect 2798 1855 2799 1862
rect 2782 1852 2783 1855
rect 2798 1852 2811 1855
rect 2734 1848 2764 1849
rect 2773 1848 2779 1849
rect 2782 1848 2811 1852
rect 2701 1847 2811 1848
rect 2701 1846 2817 1847
rect 2376 1838 2427 1846
rect 2376 1826 2401 1838
rect 2408 1826 2427 1838
rect 2458 1838 2508 1846
rect 2458 1830 2474 1838
rect 2481 1836 2508 1838
rect 2517 1836 2738 1846
rect 2481 1826 2738 1836
rect 2767 1838 2817 1846
rect 2767 1829 2783 1838
rect 2376 1818 2427 1826
rect 2474 1818 2738 1826
rect 2764 1826 2783 1829
rect 2790 1826 2817 1838
rect 2764 1818 2817 1826
rect 2392 1810 2393 1818
rect 2408 1810 2421 1818
rect 2392 1802 2408 1810
rect 2389 1795 2408 1798
rect 2389 1786 2411 1795
rect 2362 1776 2411 1786
rect 2362 1770 2392 1776
rect 2411 1771 2416 1776
rect 2334 1754 2408 1770
rect 2426 1762 2456 1818
rect 2491 1808 2699 1818
rect 2734 1814 2779 1818
rect 2782 1817 2783 1818
rect 2798 1817 2811 1818
rect 2517 1778 2706 1808
rect 2532 1775 2706 1778
rect 2525 1772 2706 1775
rect 2334 1752 2347 1754
rect 2362 1752 2396 1754
rect 2334 1736 2408 1752
rect 2435 1748 2448 1762
rect 2463 1748 2479 1764
rect 2525 1759 2536 1772
rect 2318 1714 2319 1730
rect 2334 1714 2347 1736
rect 2362 1714 2392 1736
rect 2435 1732 2497 1748
rect 2525 1741 2536 1757
rect 2541 1752 2551 1772
rect 2561 1752 2575 1772
rect 2578 1759 2587 1772
rect 2603 1759 2612 1772
rect 2541 1741 2575 1752
rect 2578 1741 2587 1757
rect 2603 1741 2612 1757
rect 2619 1752 2629 1772
rect 2639 1752 2653 1772
rect 2654 1759 2665 1772
rect 2619 1741 2653 1752
rect 2654 1741 2665 1757
rect 2711 1748 2727 1764
rect 2734 1762 2764 1814
rect 2798 1810 2799 1817
rect 2783 1802 2799 1810
rect 2770 1770 2783 1789
rect 2798 1770 2828 1786
rect 2770 1754 2844 1770
rect 2770 1752 2783 1754
rect 2798 1752 2832 1754
rect 2435 1730 2448 1732
rect 2463 1730 2497 1732
rect 2435 1714 2497 1730
rect 2541 1725 2557 1728
rect 2619 1725 2649 1736
rect 2697 1732 2743 1748
rect 2770 1736 2844 1752
rect 2697 1730 2731 1732
rect 2696 1714 2743 1730
rect 2770 1714 2783 1736
rect 2798 1714 2828 1736
rect 2855 1714 2856 1730
rect 2871 1714 2884 1874
rect 2914 1770 2927 1874
rect 2972 1852 2973 1862
rect 2988 1852 3001 1862
rect 2972 1848 3001 1852
rect 3006 1848 3036 1874
rect 3054 1860 3070 1862
rect 3142 1860 3195 1874
rect 3143 1858 3205 1860
rect 3250 1858 3265 1874
rect 3314 1871 3344 1874
rect 3314 1868 3350 1871
rect 3280 1860 3296 1862
rect 3054 1848 3069 1852
rect 2972 1846 3069 1848
rect 3097 1846 3265 1858
rect 3281 1848 3296 1852
rect 3314 1849 3353 1868
rect 3372 1862 3379 1863
rect 3378 1855 3379 1862
rect 3362 1852 3363 1855
rect 3378 1852 3391 1855
rect 3314 1848 3344 1849
rect 3353 1848 3359 1849
rect 3362 1848 3391 1852
rect 3281 1847 3391 1848
rect 3281 1846 3397 1847
rect 2956 1838 3007 1846
rect 2956 1826 2981 1838
rect 2988 1826 3007 1838
rect 3038 1838 3088 1846
rect 3038 1830 3054 1838
rect 3061 1836 3088 1838
rect 3097 1836 3318 1846
rect 3061 1826 3318 1836
rect 3347 1838 3397 1846
rect 3347 1829 3363 1838
rect 2956 1818 3007 1826
rect 3054 1818 3318 1826
rect 3344 1826 3363 1829
rect 3370 1826 3397 1838
rect 3344 1818 3397 1826
rect 2972 1810 2973 1818
rect 2988 1810 3001 1818
rect 2972 1802 2988 1810
rect 2969 1795 2988 1798
rect 2969 1786 2991 1795
rect 2942 1776 2991 1786
rect 2942 1770 2972 1776
rect 2991 1771 2996 1776
rect 2914 1754 2988 1770
rect 3006 1762 3036 1818
rect 3071 1808 3279 1818
rect 3314 1814 3359 1818
rect 3362 1817 3363 1818
rect 3378 1817 3391 1818
rect 3097 1778 3286 1808
rect 3112 1775 3286 1778
rect 3105 1772 3286 1775
rect 2914 1752 2927 1754
rect 2942 1752 2976 1754
rect 2914 1736 2988 1752
rect 3015 1748 3028 1762
rect 3043 1748 3059 1764
rect 3105 1759 3116 1772
rect 2898 1714 2899 1730
rect 2914 1714 2927 1736
rect 2942 1714 2972 1736
rect 3015 1732 3077 1748
rect 3105 1741 3116 1757
rect 3121 1752 3131 1772
rect 3141 1752 3155 1772
rect 3158 1759 3167 1772
rect 3183 1759 3192 1772
rect 3121 1741 3155 1752
rect 3158 1741 3167 1757
rect 3183 1741 3192 1757
rect 3199 1752 3209 1772
rect 3219 1752 3233 1772
rect 3234 1759 3245 1772
rect 3199 1741 3233 1752
rect 3234 1741 3245 1757
rect 3291 1748 3307 1764
rect 3314 1762 3344 1814
rect 3378 1810 3379 1817
rect 3363 1802 3379 1810
rect 3350 1770 3363 1789
rect 3378 1770 3408 1786
rect 3350 1754 3424 1770
rect 3350 1752 3363 1754
rect 3378 1752 3412 1754
rect 3015 1730 3028 1732
rect 3043 1730 3077 1732
rect 3015 1714 3077 1730
rect 3121 1725 3137 1728
rect 3199 1725 3229 1736
rect 3277 1732 3323 1748
rect 3350 1736 3424 1752
rect 3277 1730 3311 1732
rect 3276 1714 3323 1730
rect 3350 1714 3363 1736
rect 3378 1714 3408 1736
rect 3435 1714 3436 1730
rect 3451 1714 3464 1874
rect 3494 1770 3507 1874
rect 3552 1852 3553 1862
rect 3568 1852 3581 1862
rect 3552 1848 3581 1852
rect 3586 1848 3616 1874
rect 3634 1860 3650 1862
rect 3722 1860 3775 1874
rect 3723 1858 3787 1860
rect 3830 1858 3845 1874
rect 3894 1871 3924 1874
rect 3894 1868 3930 1871
rect 3860 1860 3876 1862
rect 3634 1848 3649 1852
rect 3552 1846 3649 1848
rect 3677 1846 3845 1858
rect 3861 1848 3876 1852
rect 3894 1849 3933 1868
rect 3952 1862 3959 1863
rect 3958 1855 3959 1862
rect 3942 1852 3943 1855
rect 3958 1852 3971 1855
rect 3894 1848 3924 1849
rect 3933 1848 3939 1849
rect 3942 1848 3971 1852
rect 3861 1847 3971 1848
rect 3861 1846 3977 1847
rect 3536 1838 3587 1846
rect 3536 1826 3561 1838
rect 3568 1826 3587 1838
rect 3618 1838 3668 1846
rect 3618 1830 3634 1838
rect 3641 1836 3668 1838
rect 3677 1836 3898 1846
rect 3641 1826 3898 1836
rect 3927 1838 3977 1846
rect 3927 1829 3943 1838
rect 3536 1818 3587 1826
rect 3634 1818 3898 1826
rect 3924 1826 3943 1829
rect 3950 1826 3977 1838
rect 3924 1818 3977 1826
rect 3552 1810 3553 1818
rect 3568 1810 3581 1818
rect 3552 1802 3568 1810
rect 3549 1795 3568 1798
rect 3549 1786 3571 1795
rect 3522 1776 3571 1786
rect 3522 1770 3552 1776
rect 3571 1771 3576 1776
rect 3494 1754 3568 1770
rect 3586 1762 3616 1818
rect 3651 1808 3859 1818
rect 3894 1814 3939 1818
rect 3942 1817 3943 1818
rect 3958 1817 3971 1818
rect 3677 1778 3866 1808
rect 3692 1775 3866 1778
rect 3685 1772 3866 1775
rect 3494 1752 3507 1754
rect 3522 1752 3556 1754
rect 3494 1736 3568 1752
rect 3595 1748 3608 1762
rect 3623 1748 3639 1764
rect 3685 1759 3696 1772
rect 3478 1714 3479 1730
rect 3494 1714 3507 1736
rect 3522 1714 3552 1736
rect 3595 1732 3657 1748
rect 3685 1741 3696 1757
rect 3701 1752 3711 1772
rect 3721 1752 3735 1772
rect 3738 1759 3747 1772
rect 3763 1759 3772 1772
rect 3701 1741 3735 1752
rect 3738 1741 3747 1757
rect 3763 1741 3772 1757
rect 3779 1752 3789 1772
rect 3799 1752 3813 1772
rect 3814 1759 3825 1772
rect 3779 1741 3813 1752
rect 3814 1741 3825 1757
rect 3871 1748 3887 1764
rect 3894 1762 3924 1814
rect 3958 1810 3959 1817
rect 3943 1802 3959 1810
rect 3930 1770 3943 1789
rect 3958 1770 3988 1786
rect 3930 1754 4004 1770
rect 3930 1752 3943 1754
rect 3958 1752 3992 1754
rect 3595 1730 3608 1732
rect 3623 1730 3657 1732
rect 3595 1714 3657 1730
rect 3701 1725 3717 1728
rect 3779 1725 3809 1736
rect 3857 1732 3903 1748
rect 3930 1736 4004 1752
rect 3857 1730 3891 1732
rect 3856 1714 3903 1730
rect 3930 1714 3943 1736
rect 3958 1714 3988 1736
rect 4015 1714 4016 1730
rect 4031 1714 4044 1874
rect 4074 1770 4087 1874
rect 4132 1852 4133 1862
rect 4148 1852 4161 1862
rect 4132 1848 4161 1852
rect 4166 1848 4196 1874
rect 4214 1860 4230 1862
rect 4302 1860 4355 1874
rect 4303 1858 4367 1860
rect 4410 1858 4425 1874
rect 4474 1871 4504 1874
rect 4474 1868 4510 1871
rect 4440 1860 4456 1862
rect 4214 1848 4229 1852
rect 4132 1846 4229 1848
rect 4257 1846 4425 1858
rect 4441 1848 4456 1852
rect 4474 1849 4513 1868
rect 4532 1862 4539 1863
rect 4538 1855 4539 1862
rect 4522 1852 4523 1855
rect 4538 1852 4551 1855
rect 4474 1848 4504 1849
rect 4513 1848 4519 1849
rect 4522 1848 4551 1852
rect 4441 1847 4551 1848
rect 4441 1846 4557 1847
rect 4116 1838 4167 1846
rect 4116 1826 4141 1838
rect 4148 1826 4167 1838
rect 4198 1838 4248 1846
rect 4198 1830 4214 1838
rect 4221 1836 4248 1838
rect 4257 1836 4478 1846
rect 4221 1826 4478 1836
rect 4507 1838 4557 1846
rect 4507 1829 4523 1838
rect 4116 1818 4167 1826
rect 4214 1818 4478 1826
rect 4504 1826 4523 1829
rect 4530 1826 4557 1838
rect 4504 1818 4557 1826
rect 4132 1810 4133 1818
rect 4148 1810 4161 1818
rect 4132 1802 4148 1810
rect 4129 1795 4148 1798
rect 4129 1786 4151 1795
rect 4102 1776 4151 1786
rect 4102 1770 4132 1776
rect 4151 1771 4156 1776
rect 4074 1754 4148 1770
rect 4166 1762 4196 1818
rect 4231 1808 4439 1818
rect 4474 1814 4519 1818
rect 4522 1817 4523 1818
rect 4538 1817 4551 1818
rect 4257 1778 4446 1808
rect 4272 1775 4446 1778
rect 4265 1772 4446 1775
rect 4074 1752 4087 1754
rect 4102 1752 4136 1754
rect 4074 1736 4148 1752
rect 4175 1748 4188 1762
rect 4203 1748 4219 1764
rect 4265 1759 4276 1772
rect 4058 1714 4059 1730
rect 4074 1714 4087 1736
rect 4102 1714 4132 1736
rect 4175 1732 4237 1748
rect 4265 1741 4276 1757
rect 4281 1752 4291 1772
rect 4301 1752 4315 1772
rect 4318 1759 4327 1772
rect 4343 1759 4352 1772
rect 4281 1741 4315 1752
rect 4318 1741 4327 1757
rect 4343 1741 4352 1757
rect 4359 1752 4369 1772
rect 4379 1752 4393 1772
rect 4394 1759 4405 1772
rect 4359 1741 4393 1752
rect 4394 1741 4405 1757
rect 4451 1748 4467 1764
rect 4474 1762 4504 1814
rect 4538 1810 4539 1817
rect 4523 1802 4539 1810
rect 4510 1770 4523 1789
rect 4538 1770 4568 1786
rect 4510 1754 4584 1770
rect 4510 1752 4523 1754
rect 4538 1752 4572 1754
rect 4175 1730 4188 1732
rect 4203 1730 4237 1732
rect 4175 1714 4237 1730
rect 4281 1725 4297 1728
rect 4359 1725 4389 1736
rect 4437 1732 4483 1748
rect 4510 1736 4584 1752
rect 4437 1730 4471 1732
rect 4436 1714 4483 1730
rect 4510 1714 4523 1736
rect 4538 1714 4568 1736
rect 4595 1714 4596 1730
rect 4611 1714 4624 1874
rect 4654 1770 4667 1874
rect 4712 1852 4713 1862
rect 4733 1860 4741 1862
rect 4731 1858 4741 1860
rect 4728 1852 4741 1858
rect 4712 1848 4741 1852
rect 4746 1848 4776 1874
rect 4794 1860 4810 1862
rect 4882 1860 4933 1874
rect 4883 1858 4947 1860
rect 4990 1858 5005 1874
rect 5054 1871 5084 1874
rect 5054 1868 5090 1871
rect 5020 1860 5036 1862
rect 4794 1848 4809 1852
rect 4712 1846 4809 1848
rect 4837 1846 5005 1858
rect 5021 1848 5036 1852
rect 5054 1849 5093 1868
rect 5112 1862 5119 1863
rect 5118 1855 5119 1862
rect 5102 1852 5103 1855
rect 5118 1852 5131 1855
rect 5054 1848 5084 1849
rect 5093 1848 5099 1849
rect 5102 1848 5131 1852
rect 5021 1847 5131 1848
rect 5021 1846 5137 1847
rect 4696 1838 4747 1846
rect 4696 1826 4721 1838
rect 4728 1826 4747 1838
rect 4778 1838 4828 1846
rect 4778 1830 4794 1838
rect 4801 1836 4828 1838
rect 4837 1836 5058 1846
rect 4801 1826 5058 1836
rect 5087 1838 5137 1846
rect 5087 1829 5103 1838
rect 4696 1818 4747 1826
rect 4794 1818 5058 1826
rect 5084 1826 5103 1829
rect 5110 1826 5137 1838
rect 5084 1818 5137 1826
rect 4712 1810 4713 1818
rect 4728 1810 4741 1818
rect 4712 1802 4728 1810
rect 4709 1795 4728 1798
rect 4709 1786 4731 1795
rect 4682 1776 4731 1786
rect 4682 1770 4712 1776
rect 4731 1771 4736 1776
rect 4654 1754 4728 1770
rect 4746 1762 4776 1818
rect 4811 1808 5019 1818
rect 5054 1814 5099 1818
rect 5102 1817 5103 1818
rect 5118 1817 5131 1818
rect 4837 1778 5026 1808
rect 4852 1775 5026 1778
rect 4845 1772 5026 1775
rect 4654 1752 4667 1754
rect 4682 1752 4716 1754
rect 4654 1736 4728 1752
rect 4755 1748 4768 1762
rect 4783 1748 4799 1764
rect 4845 1759 4856 1772
rect 4638 1714 4639 1730
rect 4654 1714 4667 1736
rect 4682 1714 4712 1736
rect 4755 1732 4817 1748
rect 4845 1741 4856 1757
rect 4861 1752 4871 1772
rect 4881 1752 4895 1772
rect 4898 1759 4907 1772
rect 4923 1759 4932 1772
rect 4861 1741 4895 1752
rect 4898 1741 4907 1757
rect 4923 1741 4932 1757
rect 4939 1752 4949 1772
rect 4959 1752 4973 1772
rect 4974 1759 4985 1772
rect 4939 1741 4973 1752
rect 4974 1741 4985 1757
rect 5031 1748 5047 1764
rect 5054 1762 5084 1814
rect 5118 1810 5119 1817
rect 5103 1802 5119 1810
rect 5090 1770 5103 1789
rect 5118 1770 5148 1786
rect 5090 1754 5164 1770
rect 5090 1752 5103 1754
rect 5118 1752 5152 1754
rect 4755 1730 4768 1732
rect 4783 1730 4817 1732
rect 4755 1714 4817 1730
rect 4861 1725 4877 1728
rect 4939 1725 4969 1736
rect 5017 1732 5063 1748
rect 5090 1736 5164 1752
rect 5017 1730 5051 1732
rect 5016 1714 5063 1730
rect 5090 1714 5103 1736
rect 5118 1714 5148 1736
rect 5175 1714 5176 1730
rect 5191 1714 5204 1874
rect 5234 1770 5247 1874
rect 5292 1852 5293 1862
rect 5313 1860 5321 1862
rect 5311 1858 5321 1860
rect 5308 1852 5321 1858
rect 5292 1848 5321 1852
rect 5326 1848 5356 1874
rect 5374 1860 5390 1862
rect 5462 1860 5513 1874
rect 5463 1858 5527 1860
rect 5570 1858 5585 1874
rect 5634 1871 5664 1874
rect 5634 1868 5670 1871
rect 5600 1860 5616 1862
rect 5374 1848 5389 1852
rect 5292 1846 5389 1848
rect 5417 1846 5585 1858
rect 5601 1848 5616 1852
rect 5634 1849 5673 1868
rect 5692 1862 5699 1863
rect 5698 1855 5699 1862
rect 5682 1852 5683 1855
rect 5698 1852 5711 1855
rect 5634 1848 5664 1849
rect 5673 1848 5679 1849
rect 5682 1848 5711 1852
rect 5601 1847 5711 1848
rect 5601 1846 5717 1847
rect 5276 1838 5327 1846
rect 5276 1826 5301 1838
rect 5308 1826 5327 1838
rect 5358 1838 5408 1846
rect 5358 1830 5374 1838
rect 5381 1836 5408 1838
rect 5417 1836 5638 1846
rect 5381 1826 5638 1836
rect 5667 1838 5717 1846
rect 5667 1829 5683 1838
rect 5276 1818 5327 1826
rect 5374 1818 5638 1826
rect 5664 1826 5683 1829
rect 5690 1826 5717 1838
rect 5664 1818 5717 1826
rect 5292 1810 5293 1818
rect 5308 1810 5321 1818
rect 5292 1802 5308 1810
rect 5289 1795 5308 1798
rect 5289 1786 5311 1795
rect 5262 1776 5311 1786
rect 5262 1770 5292 1776
rect 5311 1771 5316 1776
rect 5234 1754 5308 1770
rect 5326 1762 5356 1818
rect 5391 1808 5599 1818
rect 5634 1814 5679 1818
rect 5682 1817 5683 1818
rect 5698 1817 5711 1818
rect 5417 1778 5606 1808
rect 5432 1775 5606 1778
rect 5425 1772 5606 1775
rect 5234 1752 5247 1754
rect 5262 1752 5296 1754
rect 5234 1736 5308 1752
rect 5335 1748 5348 1762
rect 5363 1748 5379 1764
rect 5425 1759 5436 1772
rect 5218 1714 5219 1730
rect 5234 1714 5247 1736
rect 5262 1714 5292 1736
rect 5335 1732 5397 1748
rect 5425 1741 5436 1757
rect 5441 1752 5451 1772
rect 5461 1752 5475 1772
rect 5478 1759 5487 1772
rect 5503 1759 5512 1772
rect 5441 1741 5475 1752
rect 5478 1741 5487 1757
rect 5503 1741 5512 1757
rect 5519 1752 5529 1772
rect 5539 1752 5553 1772
rect 5554 1759 5565 1772
rect 5519 1741 5553 1752
rect 5554 1741 5565 1757
rect 5611 1748 5627 1764
rect 5634 1762 5664 1814
rect 5698 1810 5699 1817
rect 5683 1802 5699 1810
rect 5670 1770 5683 1789
rect 5698 1770 5728 1786
rect 5670 1754 5744 1770
rect 5670 1752 5683 1754
rect 5698 1752 5732 1754
rect 5335 1730 5348 1732
rect 5363 1730 5397 1732
rect 5335 1714 5397 1730
rect 5441 1725 5457 1728
rect 5519 1725 5549 1736
rect 5597 1732 5643 1748
rect 5670 1736 5744 1752
rect 5597 1730 5631 1732
rect 5596 1714 5643 1730
rect 5670 1714 5683 1736
rect 5698 1714 5728 1736
rect 5755 1714 5756 1730
rect 5771 1714 5784 1874
rect 5814 1770 5827 1874
rect 5872 1852 5873 1862
rect 5893 1860 5901 1862
rect 5891 1858 5901 1860
rect 5888 1852 5901 1858
rect 5872 1848 5901 1852
rect 5906 1848 5936 1874
rect 5954 1860 5970 1862
rect 6042 1860 6093 1874
rect 6043 1858 6107 1860
rect 6150 1858 6165 1874
rect 6214 1871 6244 1874
rect 6214 1868 6250 1871
rect 6180 1860 6196 1862
rect 5954 1848 5969 1852
rect 5872 1846 5969 1848
rect 5997 1846 6165 1858
rect 6181 1848 6196 1852
rect 6214 1849 6253 1868
rect 6272 1862 6279 1863
rect 6278 1855 6279 1862
rect 6262 1852 6263 1855
rect 6278 1852 6291 1855
rect 6214 1848 6244 1849
rect 6253 1848 6259 1849
rect 6262 1848 6291 1852
rect 6181 1847 6291 1848
rect 6181 1846 6297 1847
rect 5856 1838 5907 1846
rect 5856 1826 5881 1838
rect 5888 1826 5907 1838
rect 5938 1838 5988 1846
rect 5938 1830 5954 1838
rect 5961 1836 5988 1838
rect 5997 1836 6218 1846
rect 5961 1826 6218 1836
rect 6247 1838 6297 1846
rect 6247 1829 6263 1838
rect 5856 1818 5907 1826
rect 5954 1818 6218 1826
rect 6244 1826 6263 1829
rect 6270 1826 6297 1838
rect 6244 1818 6297 1826
rect 5872 1810 5873 1818
rect 5888 1810 5901 1818
rect 5872 1802 5888 1810
rect 5869 1795 5888 1798
rect 5869 1786 5891 1795
rect 5842 1776 5891 1786
rect 5842 1770 5872 1776
rect 5891 1771 5896 1776
rect 5814 1754 5888 1770
rect 5906 1762 5936 1818
rect 5971 1808 6179 1818
rect 6214 1814 6259 1818
rect 6262 1817 6263 1818
rect 6278 1817 6291 1818
rect 5997 1778 6186 1808
rect 6012 1775 6186 1778
rect 6005 1772 6186 1775
rect 5814 1752 5827 1754
rect 5842 1752 5876 1754
rect 5814 1736 5888 1752
rect 5915 1748 5928 1762
rect 5943 1748 5959 1764
rect 6005 1759 6016 1772
rect 5798 1714 5799 1730
rect 5814 1714 5827 1736
rect 5842 1714 5872 1736
rect 5915 1732 5977 1748
rect 6005 1741 6016 1757
rect 6021 1752 6031 1772
rect 6041 1752 6055 1772
rect 6058 1759 6067 1772
rect 6083 1759 6092 1772
rect 6021 1741 6055 1752
rect 6058 1741 6067 1757
rect 6083 1741 6092 1757
rect 6099 1752 6109 1772
rect 6119 1752 6133 1772
rect 6134 1759 6145 1772
rect 6099 1741 6133 1752
rect 6134 1741 6145 1757
rect 6191 1748 6207 1764
rect 6214 1762 6244 1814
rect 6278 1810 6279 1817
rect 6263 1802 6279 1810
rect 6250 1770 6263 1789
rect 6278 1770 6308 1786
rect 6250 1754 6324 1770
rect 6250 1752 6263 1754
rect 6278 1752 6312 1754
rect 5915 1730 5928 1732
rect 5943 1730 5977 1732
rect 5915 1714 5977 1730
rect 6021 1725 6037 1728
rect 6099 1725 6129 1736
rect 6177 1732 6223 1748
rect 6250 1736 6324 1752
rect 6177 1730 6211 1732
rect 6176 1714 6223 1730
rect 6250 1714 6263 1736
rect 6278 1714 6308 1736
rect 6335 1714 6336 1730
rect 6351 1714 6364 1874
rect 6394 1770 6407 1874
rect 6452 1852 6453 1862
rect 6473 1860 6481 1862
rect 6471 1858 6481 1860
rect 6468 1852 6481 1858
rect 6452 1848 6481 1852
rect 6486 1848 6516 1874
rect 6534 1860 6550 1862
rect 6622 1860 6673 1874
rect 6623 1858 6687 1860
rect 6730 1858 6745 1874
rect 6794 1871 6824 1874
rect 6794 1868 6830 1871
rect 6760 1860 6776 1862
rect 6534 1848 6549 1852
rect 6452 1846 6549 1848
rect 6577 1846 6745 1858
rect 6761 1848 6776 1852
rect 6794 1849 6833 1868
rect 6852 1862 6859 1863
rect 6858 1855 6859 1862
rect 6842 1852 6843 1855
rect 6858 1852 6871 1855
rect 6794 1848 6824 1849
rect 6833 1848 6839 1849
rect 6842 1848 6871 1852
rect 6761 1847 6871 1848
rect 6761 1846 6877 1847
rect 6436 1838 6487 1846
rect 6436 1826 6461 1838
rect 6468 1826 6487 1838
rect 6518 1838 6568 1846
rect 6518 1830 6534 1838
rect 6541 1836 6568 1838
rect 6577 1836 6798 1846
rect 6541 1826 6798 1836
rect 6827 1838 6877 1846
rect 6827 1829 6843 1838
rect 6436 1818 6487 1826
rect 6534 1818 6798 1826
rect 6824 1826 6843 1829
rect 6850 1826 6877 1838
rect 6824 1818 6877 1826
rect 6452 1810 6453 1818
rect 6468 1810 6481 1818
rect 6452 1802 6468 1810
rect 6449 1795 6468 1798
rect 6449 1786 6471 1795
rect 6422 1776 6471 1786
rect 6422 1770 6452 1776
rect 6471 1771 6476 1776
rect 6394 1754 6468 1770
rect 6486 1762 6516 1818
rect 6551 1808 6759 1818
rect 6794 1814 6839 1818
rect 6842 1817 6843 1818
rect 6858 1817 6871 1818
rect 6577 1778 6766 1808
rect 6592 1775 6766 1778
rect 6585 1772 6766 1775
rect 6394 1752 6407 1754
rect 6422 1752 6456 1754
rect 6394 1736 6468 1752
rect 6495 1748 6508 1762
rect 6523 1748 6539 1764
rect 6585 1759 6596 1772
rect 6378 1714 6379 1730
rect 6394 1714 6407 1736
rect 6422 1714 6452 1736
rect 6495 1732 6557 1748
rect 6585 1741 6596 1757
rect 6601 1752 6611 1772
rect 6621 1752 6635 1772
rect 6638 1759 6647 1772
rect 6663 1759 6672 1772
rect 6601 1741 6635 1752
rect 6638 1741 6647 1757
rect 6663 1741 6672 1757
rect 6679 1752 6689 1772
rect 6699 1752 6713 1772
rect 6714 1759 6725 1772
rect 6679 1741 6713 1752
rect 6714 1741 6725 1757
rect 6771 1748 6787 1764
rect 6794 1762 6824 1814
rect 6858 1810 6859 1817
rect 6843 1802 6859 1810
rect 6830 1770 6843 1789
rect 6858 1770 6888 1786
rect 6830 1754 6904 1770
rect 6830 1752 6843 1754
rect 6858 1752 6892 1754
rect 6495 1730 6508 1732
rect 6523 1730 6557 1732
rect 6495 1714 6557 1730
rect 6601 1725 6617 1728
rect 6679 1725 6709 1736
rect 6757 1732 6803 1748
rect 6830 1736 6904 1752
rect 6757 1730 6791 1732
rect 6756 1714 6803 1730
rect 6830 1714 6843 1736
rect 6858 1714 6888 1736
rect 6915 1714 6916 1730
rect 6931 1714 6944 1874
rect 0 1706 33 1714
rect 0 1680 7 1706
rect 14 1680 33 1706
rect 97 1702 159 1714
rect 171 1702 246 1714
rect 304 1702 379 1714
rect 391 1702 422 1714
rect 428 1702 463 1714
rect 97 1700 259 1702
rect 0 1672 33 1680
rect 115 1676 128 1700
rect 143 1698 158 1700
rect 14 1662 27 1672
rect 42 1662 72 1676
rect 115 1662 158 1676
rect 182 1673 189 1680
rect 192 1676 259 1700
rect 291 1700 463 1702
rect 261 1678 289 1682
rect 291 1678 371 1700
rect 392 1698 407 1700
rect 261 1676 371 1678
rect 192 1672 371 1676
rect 165 1662 195 1672
rect 197 1662 350 1672
rect 358 1662 388 1672
rect 392 1662 422 1676
rect 450 1662 463 1700
rect 535 1706 570 1714
rect 535 1680 536 1706
rect 543 1680 570 1706
rect 478 1662 508 1676
rect 535 1672 570 1680
rect 572 1706 613 1714
rect 572 1680 587 1706
rect 594 1680 613 1706
rect 677 1702 739 1714
rect 751 1702 826 1714
rect 884 1702 959 1714
rect 971 1702 1002 1714
rect 1008 1702 1043 1714
rect 677 1700 839 1702
rect 572 1672 613 1680
rect 695 1676 708 1700
rect 723 1698 738 1700
rect 535 1662 536 1672
rect 551 1662 564 1672
rect 578 1662 579 1672
rect 594 1662 607 1672
rect 622 1662 652 1676
rect 695 1662 738 1676
rect 762 1673 769 1680
rect 772 1676 839 1700
rect 871 1700 1043 1702
rect 841 1678 869 1682
rect 871 1678 951 1700
rect 972 1698 987 1700
rect 841 1676 951 1678
rect 772 1672 951 1676
rect 745 1662 775 1672
rect 777 1662 930 1672
rect 938 1662 968 1672
rect 972 1662 1002 1676
rect 1030 1662 1043 1700
rect 1115 1706 1150 1714
rect 1115 1680 1116 1706
rect 1123 1680 1150 1706
rect 1058 1662 1088 1676
rect 1115 1672 1150 1680
rect 1152 1706 1193 1714
rect 1152 1680 1167 1706
rect 1174 1680 1193 1706
rect 1257 1702 1319 1714
rect 1331 1702 1406 1714
rect 1464 1702 1539 1714
rect 1551 1702 1582 1714
rect 1588 1702 1623 1714
rect 1257 1700 1419 1702
rect 1152 1672 1193 1680
rect 1275 1676 1288 1700
rect 1303 1698 1318 1700
rect 1115 1662 1116 1672
rect 1131 1662 1144 1672
rect 1158 1662 1159 1672
rect 1174 1662 1187 1672
rect 1202 1662 1232 1676
rect 1275 1662 1318 1676
rect 1342 1673 1349 1680
rect 1352 1676 1419 1700
rect 1451 1700 1623 1702
rect 1421 1678 1449 1682
rect 1451 1678 1531 1700
rect 1552 1698 1567 1700
rect 1421 1676 1531 1678
rect 1352 1672 1531 1676
rect 1325 1662 1355 1672
rect 1357 1662 1510 1672
rect 1518 1662 1548 1672
rect 1552 1662 1582 1676
rect 1610 1662 1623 1700
rect 1695 1706 1730 1714
rect 1695 1680 1696 1706
rect 1703 1680 1730 1706
rect 1638 1662 1668 1676
rect 1695 1672 1730 1680
rect 1732 1706 1773 1714
rect 1732 1680 1747 1706
rect 1754 1680 1773 1706
rect 1837 1702 1899 1714
rect 1911 1702 1986 1714
rect 2044 1702 2119 1714
rect 2131 1702 2162 1714
rect 2168 1702 2203 1714
rect 1837 1700 1999 1702
rect 1732 1672 1773 1680
rect 1855 1676 1868 1700
rect 1883 1698 1898 1700
rect 1695 1662 1696 1672
rect 1711 1662 1724 1672
rect 1738 1662 1739 1672
rect 1754 1662 1767 1672
rect 1782 1662 1812 1676
rect 1855 1662 1898 1676
rect 1922 1673 1929 1680
rect 1932 1676 1999 1700
rect 2031 1700 2203 1702
rect 2001 1678 2029 1682
rect 2031 1678 2111 1700
rect 2132 1698 2147 1700
rect 2001 1676 2111 1678
rect 1932 1672 2111 1676
rect 1905 1662 1935 1672
rect 1937 1662 2090 1672
rect 2098 1662 2128 1672
rect 2132 1662 2162 1676
rect 2190 1662 2203 1700
rect 2275 1706 2310 1714
rect 2275 1680 2276 1706
rect 2283 1680 2310 1706
rect 2218 1662 2248 1676
rect 2275 1672 2310 1680
rect 2312 1706 2353 1714
rect 2312 1680 2327 1706
rect 2334 1680 2353 1706
rect 2417 1702 2479 1714
rect 2491 1702 2566 1714
rect 2624 1702 2699 1714
rect 2711 1702 2742 1714
rect 2748 1702 2783 1714
rect 2417 1700 2579 1702
rect 2312 1672 2353 1680
rect 2435 1676 2448 1700
rect 2463 1698 2478 1700
rect 2275 1662 2276 1672
rect 2291 1662 2304 1672
rect 2318 1662 2319 1672
rect 2334 1662 2347 1672
rect 2362 1662 2392 1676
rect 2435 1662 2478 1676
rect 2502 1673 2509 1680
rect 2512 1676 2579 1700
rect 2611 1700 2783 1702
rect 2581 1678 2609 1682
rect 2611 1678 2691 1700
rect 2712 1698 2727 1700
rect 2581 1676 2691 1678
rect 2512 1672 2691 1676
rect 2485 1662 2515 1672
rect 2517 1662 2670 1672
rect 2678 1662 2708 1672
rect 2712 1662 2742 1676
rect 2770 1662 2783 1700
rect 2855 1706 2890 1714
rect 2855 1680 2856 1706
rect 2863 1680 2890 1706
rect 2798 1662 2828 1676
rect 2855 1672 2890 1680
rect 2892 1706 2933 1714
rect 2892 1680 2907 1706
rect 2914 1680 2933 1706
rect 2997 1702 3059 1714
rect 3071 1702 3146 1714
rect 3204 1702 3279 1714
rect 3291 1702 3322 1714
rect 3328 1702 3363 1714
rect 2997 1700 3159 1702
rect 2892 1672 2933 1680
rect 3015 1676 3028 1700
rect 3043 1698 3058 1700
rect 2855 1662 2856 1672
rect 2871 1662 2884 1672
rect 2898 1662 2899 1672
rect 2914 1662 2927 1672
rect 2942 1662 2972 1676
rect 3015 1662 3058 1676
rect 3082 1673 3089 1680
rect 3092 1676 3159 1700
rect 3191 1700 3363 1702
rect 3161 1678 3189 1682
rect 3191 1678 3271 1700
rect 3292 1698 3307 1700
rect 3161 1676 3271 1678
rect 3092 1672 3271 1676
rect 3065 1662 3095 1672
rect 3097 1662 3250 1672
rect 3258 1662 3288 1672
rect 3292 1662 3322 1676
rect 3350 1662 3363 1700
rect 3435 1706 3470 1714
rect 3435 1680 3436 1706
rect 3443 1680 3470 1706
rect 3378 1662 3408 1676
rect 3435 1672 3470 1680
rect 3472 1706 3513 1714
rect 3472 1680 3487 1706
rect 3494 1680 3513 1706
rect 3577 1702 3639 1714
rect 3651 1702 3726 1714
rect 3784 1702 3859 1714
rect 3871 1702 3902 1714
rect 3908 1702 3943 1714
rect 3577 1700 3739 1702
rect 3472 1672 3513 1680
rect 3595 1676 3608 1700
rect 3623 1698 3638 1700
rect 3435 1662 3436 1672
rect 3451 1662 3464 1672
rect 3478 1662 3479 1672
rect 3494 1662 3507 1672
rect 3522 1662 3552 1676
rect 3595 1662 3638 1676
rect 3662 1673 3669 1680
rect 3672 1676 3739 1700
rect 3771 1700 3943 1702
rect 3741 1678 3769 1682
rect 3771 1678 3851 1700
rect 3872 1698 3887 1700
rect 3741 1676 3851 1678
rect 3672 1672 3851 1676
rect 3645 1662 3675 1672
rect 3677 1662 3830 1672
rect 3838 1662 3868 1672
rect 3872 1662 3902 1676
rect 3930 1662 3943 1700
rect 4015 1706 4050 1714
rect 4015 1680 4016 1706
rect 4023 1680 4050 1706
rect 3958 1662 3988 1676
rect 4015 1672 4050 1680
rect 4052 1706 4093 1714
rect 4052 1680 4067 1706
rect 4074 1680 4093 1706
rect 4157 1702 4219 1714
rect 4231 1702 4306 1714
rect 4364 1702 4439 1714
rect 4451 1702 4482 1714
rect 4488 1702 4523 1714
rect 4157 1700 4319 1702
rect 4052 1672 4093 1680
rect 4175 1676 4188 1700
rect 4203 1698 4218 1700
rect 4015 1662 4016 1672
rect 4031 1662 4044 1672
rect 4058 1662 4059 1672
rect 4074 1662 4087 1672
rect 4102 1662 4132 1676
rect 4175 1662 4218 1676
rect 4242 1673 4249 1680
rect 4252 1676 4319 1700
rect 4351 1700 4523 1702
rect 4321 1678 4349 1682
rect 4351 1678 4431 1700
rect 4452 1698 4467 1700
rect 4321 1676 4431 1678
rect 4252 1672 4431 1676
rect 4225 1662 4255 1672
rect 4257 1662 4410 1672
rect 4418 1662 4448 1672
rect 4452 1662 4482 1676
rect 4510 1662 4523 1700
rect 4595 1706 4630 1714
rect 4595 1680 4596 1706
rect 4603 1680 4630 1706
rect 4538 1662 4568 1676
rect 4595 1672 4630 1680
rect 4632 1706 4673 1714
rect 4632 1680 4647 1706
rect 4654 1680 4673 1706
rect 4737 1702 4799 1714
rect 4811 1702 4886 1714
rect 4944 1702 5019 1714
rect 5031 1702 5062 1714
rect 5068 1702 5103 1714
rect 4737 1700 4899 1702
rect 4755 1682 4768 1700
rect 4783 1698 4798 1700
rect 4632 1672 4673 1680
rect 4756 1676 4768 1682
rect 4832 1682 4899 1700
rect 4931 1700 5103 1702
rect 4931 1682 5011 1700
rect 5032 1698 5047 1700
rect 4595 1662 4596 1672
rect 4611 1662 4624 1672
rect 4638 1662 4639 1672
rect 4654 1662 4667 1672
rect 4682 1662 4712 1676
rect 4756 1662 4798 1676
rect 4822 1673 4829 1680
rect 4832 1672 5011 1682
rect 4805 1662 4835 1672
rect 4837 1662 4990 1672
rect 4998 1662 5028 1672
rect 5032 1662 5062 1676
rect 5090 1662 5103 1700
rect 5175 1706 5210 1714
rect 5175 1680 5176 1706
rect 5183 1680 5210 1706
rect 5118 1662 5148 1676
rect 5175 1672 5210 1680
rect 5212 1706 5253 1714
rect 5212 1680 5227 1706
rect 5234 1680 5253 1706
rect 5317 1702 5379 1714
rect 5391 1702 5466 1714
rect 5524 1702 5599 1714
rect 5611 1702 5642 1714
rect 5648 1702 5683 1714
rect 5317 1700 5479 1702
rect 5335 1682 5348 1700
rect 5363 1698 5378 1700
rect 5212 1672 5253 1680
rect 5336 1676 5348 1682
rect 5412 1682 5479 1700
rect 5511 1700 5683 1702
rect 5511 1682 5591 1700
rect 5612 1698 5627 1700
rect 5175 1662 5176 1672
rect 5191 1662 5204 1672
rect 5218 1662 5219 1672
rect 5234 1662 5247 1672
rect 5262 1662 5292 1676
rect 5336 1662 5378 1676
rect 5402 1673 5409 1680
rect 5412 1672 5591 1682
rect 5385 1662 5415 1672
rect 5417 1662 5570 1672
rect 5578 1662 5608 1672
rect 5612 1662 5642 1676
rect 5670 1662 5683 1700
rect 5755 1706 5790 1714
rect 5755 1680 5756 1706
rect 5763 1680 5790 1706
rect 5698 1662 5728 1676
rect 5755 1672 5790 1680
rect 5792 1706 5833 1714
rect 5792 1680 5807 1706
rect 5814 1680 5833 1706
rect 5897 1702 5959 1714
rect 5971 1702 6046 1714
rect 6104 1702 6179 1714
rect 6191 1702 6222 1714
rect 6228 1702 6263 1714
rect 5897 1700 6059 1702
rect 5915 1682 5928 1700
rect 5943 1698 5958 1700
rect 5792 1672 5833 1680
rect 5916 1676 5928 1682
rect 5992 1682 6059 1700
rect 6091 1700 6263 1702
rect 6091 1682 6171 1700
rect 6192 1698 6207 1700
rect 5755 1662 5756 1672
rect 5771 1662 5784 1672
rect 5798 1662 5799 1672
rect 5814 1662 5827 1672
rect 5842 1662 5872 1676
rect 5916 1662 5958 1676
rect 5982 1673 5989 1680
rect 5992 1672 6171 1682
rect 5965 1662 5995 1672
rect 5997 1662 6150 1672
rect 6158 1662 6188 1672
rect 6192 1662 6222 1676
rect 6250 1662 6263 1700
rect 6335 1706 6370 1714
rect 6335 1680 6336 1706
rect 6343 1680 6370 1706
rect 6278 1662 6308 1676
rect 6335 1672 6370 1680
rect 6372 1706 6413 1714
rect 6372 1680 6387 1706
rect 6394 1680 6413 1706
rect 6477 1702 6539 1714
rect 6551 1702 6626 1714
rect 6684 1702 6759 1714
rect 6771 1702 6802 1714
rect 6808 1702 6843 1714
rect 6477 1700 6639 1702
rect 6495 1682 6508 1700
rect 6523 1698 6538 1700
rect 6372 1672 6413 1680
rect 6496 1676 6508 1682
rect 6572 1682 6639 1700
rect 6671 1700 6843 1702
rect 6671 1682 6751 1700
rect 6772 1698 6787 1700
rect 6335 1662 6336 1672
rect 6351 1662 6364 1672
rect 6378 1662 6379 1672
rect 6394 1662 6407 1672
rect 6422 1662 6452 1676
rect 6496 1662 6538 1676
rect 6562 1673 6569 1680
rect 6572 1672 6751 1682
rect 6545 1662 6575 1672
rect 6577 1662 6730 1672
rect 6738 1662 6768 1672
rect 6772 1662 6802 1676
rect 6830 1662 6843 1700
rect 6915 1706 6950 1714
rect 6915 1680 6916 1706
rect 6923 1680 6950 1706
rect 6858 1662 6888 1676
rect 6915 1672 6950 1680
rect 6915 1662 6916 1672
rect 6931 1662 6944 1672
rect 0 1648 6944 1662
rect 14 1618 27 1648
rect 42 1630 72 1648
rect 115 1634 129 1648
rect 165 1634 385 1648
rect 116 1632 129 1634
rect 82 1620 97 1632
rect 79 1618 101 1620
rect 106 1618 136 1632
rect 197 1630 350 1634
rect 179 1618 371 1630
rect 414 1618 444 1632
rect 450 1618 463 1648
rect 478 1630 508 1648
rect 551 1618 564 1648
rect 594 1618 607 1648
rect 622 1630 652 1648
rect 695 1634 709 1648
rect 745 1634 965 1648
rect 696 1632 709 1634
rect 662 1620 677 1632
rect 659 1618 681 1620
rect 686 1618 716 1632
rect 777 1630 930 1634
rect 759 1618 951 1630
rect 994 1618 1024 1632
rect 1030 1618 1043 1648
rect 1058 1630 1088 1648
rect 1131 1618 1144 1648
rect 1174 1618 1187 1648
rect 1202 1630 1232 1648
rect 1275 1634 1289 1648
rect 1325 1634 1545 1648
rect 1276 1632 1289 1634
rect 1242 1620 1257 1632
rect 1239 1618 1261 1620
rect 1266 1618 1296 1632
rect 1357 1630 1510 1634
rect 1339 1618 1531 1630
rect 1574 1618 1604 1632
rect 1610 1618 1623 1648
rect 1638 1630 1668 1648
rect 1711 1618 1724 1648
rect 1754 1618 1767 1648
rect 1782 1630 1812 1648
rect 1855 1634 1869 1648
rect 1905 1634 2125 1648
rect 1856 1632 1869 1634
rect 1822 1620 1837 1632
rect 1819 1618 1841 1620
rect 1846 1618 1876 1632
rect 1937 1630 2090 1634
rect 1919 1618 2111 1630
rect 2154 1618 2184 1632
rect 2190 1618 2203 1648
rect 2218 1630 2248 1648
rect 2291 1618 2304 1648
rect 2334 1618 2347 1648
rect 2362 1630 2392 1648
rect 2435 1634 2449 1648
rect 2485 1634 2705 1648
rect 2436 1632 2449 1634
rect 2402 1620 2417 1632
rect 2399 1618 2421 1620
rect 2426 1618 2456 1632
rect 2517 1630 2670 1634
rect 2499 1618 2691 1630
rect 2734 1618 2764 1632
rect 2770 1618 2783 1648
rect 2798 1630 2828 1648
rect 2871 1618 2884 1648
rect 2914 1618 2927 1648
rect 2942 1630 2972 1648
rect 3015 1634 3029 1648
rect 3065 1634 3285 1648
rect 3016 1632 3029 1634
rect 2982 1620 2997 1632
rect 2979 1618 3001 1620
rect 3006 1618 3036 1632
rect 3097 1630 3250 1634
rect 3079 1618 3271 1630
rect 3314 1618 3344 1632
rect 3350 1618 3363 1648
rect 3378 1630 3408 1648
rect 3451 1618 3464 1648
rect 3494 1618 3507 1648
rect 3522 1630 3552 1648
rect 3595 1634 3609 1648
rect 3645 1634 3865 1648
rect 3596 1632 3609 1634
rect 3562 1620 3577 1632
rect 3559 1618 3581 1620
rect 3586 1618 3616 1632
rect 3677 1630 3830 1634
rect 3659 1618 3851 1630
rect 3894 1618 3924 1632
rect 3930 1618 3943 1648
rect 3958 1630 3988 1648
rect 4031 1618 4044 1648
rect 4074 1618 4087 1648
rect 4102 1630 4132 1648
rect 4175 1634 4189 1648
rect 4225 1634 4445 1648
rect 4176 1632 4189 1634
rect 4142 1620 4157 1632
rect 4139 1618 4161 1620
rect 4166 1618 4196 1632
rect 4257 1630 4410 1634
rect 4239 1618 4431 1630
rect 4474 1618 4504 1632
rect 4510 1618 4523 1648
rect 4538 1630 4568 1648
rect 4611 1618 4624 1648
rect 4654 1618 4667 1648
rect 4682 1630 4712 1648
rect 4756 1632 4769 1648
rect 4805 1634 5025 1648
rect 4722 1620 4737 1632
rect 4719 1618 4741 1620
rect 4746 1618 4776 1632
rect 4837 1630 4990 1634
rect 4819 1618 5011 1630
rect 5054 1618 5084 1632
rect 5090 1618 5103 1648
rect 5118 1630 5148 1648
rect 5191 1618 5204 1648
rect 5234 1618 5247 1648
rect 5262 1630 5292 1648
rect 5336 1632 5349 1648
rect 5385 1634 5605 1648
rect 5302 1620 5317 1632
rect 5299 1618 5321 1620
rect 5326 1618 5356 1632
rect 5417 1630 5570 1634
rect 5399 1618 5591 1630
rect 5634 1618 5664 1632
rect 5670 1618 5683 1648
rect 5698 1630 5728 1648
rect 5771 1618 5784 1648
rect 5814 1618 5827 1648
rect 5842 1630 5872 1648
rect 5916 1632 5929 1648
rect 5965 1634 6185 1648
rect 5882 1620 5897 1632
rect 5879 1618 5901 1620
rect 5906 1618 5936 1632
rect 5997 1630 6150 1634
rect 5979 1618 6171 1630
rect 6214 1618 6244 1632
rect 6250 1618 6263 1648
rect 6278 1630 6308 1648
rect 6351 1618 6364 1648
rect 6394 1618 6407 1648
rect 6422 1630 6452 1648
rect 6496 1632 6509 1648
rect 6545 1634 6765 1648
rect 6462 1620 6477 1632
rect 6459 1618 6481 1620
rect 6486 1618 6516 1632
rect 6577 1630 6730 1634
rect 6559 1618 6751 1630
rect 6794 1618 6824 1632
rect 6830 1618 6843 1648
rect 6858 1630 6888 1648
rect 6931 1618 6944 1648
rect 0 1604 6944 1618
rect 14 1500 27 1604
rect 72 1582 73 1592
rect 88 1582 101 1592
rect 72 1578 101 1582
rect 106 1578 136 1604
rect 154 1590 170 1592
rect 242 1590 295 1604
rect 243 1588 307 1590
rect 350 1588 365 1604
rect 414 1601 444 1604
rect 414 1598 450 1601
rect 380 1590 396 1592
rect 154 1578 169 1582
rect 72 1576 169 1578
rect 197 1576 365 1588
rect 381 1578 396 1582
rect 414 1579 453 1598
rect 472 1592 479 1593
rect 478 1585 479 1592
rect 462 1582 463 1585
rect 478 1582 491 1585
rect 414 1578 444 1579
rect 453 1578 459 1579
rect 462 1578 491 1582
rect 381 1577 491 1578
rect 381 1576 497 1577
rect 56 1568 107 1576
rect 56 1556 81 1568
rect 88 1556 107 1568
rect 138 1568 188 1576
rect 138 1560 154 1568
rect 161 1566 188 1568
rect 197 1566 418 1576
rect 161 1556 418 1566
rect 447 1568 497 1576
rect 447 1559 463 1568
rect 56 1548 107 1556
rect 154 1548 418 1556
rect 444 1556 463 1559
rect 470 1556 497 1568
rect 444 1548 497 1556
rect 72 1540 73 1548
rect 88 1540 101 1548
rect 72 1532 88 1540
rect 69 1525 88 1528
rect 69 1516 91 1525
rect 42 1506 91 1516
rect 42 1500 72 1506
rect 91 1501 96 1506
rect 14 1484 88 1500
rect 106 1492 136 1548
rect 171 1538 379 1548
rect 414 1544 459 1548
rect 462 1547 463 1548
rect 478 1547 491 1548
rect 197 1508 386 1538
rect 212 1505 386 1508
rect 205 1502 386 1505
rect 14 1482 27 1484
rect 42 1482 76 1484
rect 14 1466 88 1482
rect 115 1478 128 1492
rect 143 1478 159 1494
rect 205 1489 216 1502
rect 14 1444 27 1466
rect 42 1444 72 1466
rect 115 1462 177 1478
rect 205 1471 216 1487
rect 221 1482 231 1502
rect 241 1482 255 1502
rect 258 1489 267 1502
rect 283 1489 292 1502
rect 221 1471 255 1482
rect 258 1471 267 1487
rect 283 1471 292 1487
rect 299 1482 309 1502
rect 319 1482 333 1502
rect 334 1489 345 1502
rect 299 1471 333 1482
rect 334 1471 345 1487
rect 391 1478 407 1494
rect 414 1492 444 1544
rect 478 1540 479 1547
rect 463 1532 479 1540
rect 450 1500 463 1519
rect 478 1500 508 1516
rect 450 1484 524 1500
rect 450 1482 463 1484
rect 478 1482 512 1484
rect 115 1460 128 1462
rect 143 1460 177 1462
rect 115 1444 177 1460
rect 221 1455 237 1458
rect 299 1455 329 1466
rect 377 1462 423 1478
rect 450 1466 524 1482
rect 377 1460 411 1462
rect 376 1444 423 1460
rect 450 1444 463 1466
rect 478 1444 508 1466
rect 535 1444 536 1460
rect 551 1444 564 1604
rect 594 1500 607 1604
rect 652 1582 653 1592
rect 668 1582 681 1592
rect 652 1578 681 1582
rect 686 1578 716 1604
rect 734 1590 750 1592
rect 822 1590 875 1604
rect 823 1588 887 1590
rect 930 1588 945 1604
rect 994 1601 1024 1604
rect 994 1598 1030 1601
rect 960 1590 976 1592
rect 734 1578 749 1582
rect 652 1576 749 1578
rect 777 1576 945 1588
rect 961 1578 976 1582
rect 994 1579 1033 1598
rect 1052 1592 1059 1593
rect 1058 1585 1059 1592
rect 1042 1582 1043 1585
rect 1058 1582 1071 1585
rect 994 1578 1024 1579
rect 1033 1578 1039 1579
rect 1042 1578 1071 1582
rect 961 1577 1071 1578
rect 961 1576 1077 1577
rect 636 1568 687 1576
rect 636 1556 661 1568
rect 668 1556 687 1568
rect 718 1568 768 1576
rect 718 1560 734 1568
rect 741 1566 768 1568
rect 777 1566 998 1576
rect 741 1556 998 1566
rect 1027 1568 1077 1576
rect 1027 1559 1043 1568
rect 636 1548 687 1556
rect 734 1548 998 1556
rect 1024 1556 1043 1559
rect 1050 1556 1077 1568
rect 1024 1548 1077 1556
rect 652 1540 653 1548
rect 668 1540 681 1548
rect 652 1532 668 1540
rect 649 1525 668 1528
rect 649 1516 671 1525
rect 622 1506 671 1516
rect 622 1500 652 1506
rect 671 1501 676 1506
rect 594 1484 668 1500
rect 686 1492 716 1548
rect 751 1538 959 1548
rect 994 1544 1039 1548
rect 1042 1547 1043 1548
rect 1058 1547 1071 1548
rect 777 1508 966 1538
rect 792 1505 966 1508
rect 785 1502 966 1505
rect 594 1482 607 1484
rect 622 1482 656 1484
rect 594 1466 668 1482
rect 695 1478 708 1492
rect 723 1478 739 1494
rect 785 1489 796 1502
rect 578 1444 579 1460
rect 594 1444 607 1466
rect 622 1444 652 1466
rect 695 1462 757 1478
rect 785 1471 796 1487
rect 801 1482 811 1502
rect 821 1482 835 1502
rect 838 1489 847 1502
rect 863 1489 872 1502
rect 801 1471 835 1482
rect 838 1471 847 1487
rect 863 1471 872 1487
rect 879 1482 889 1502
rect 899 1482 913 1502
rect 914 1489 925 1502
rect 879 1471 913 1482
rect 914 1471 925 1487
rect 971 1478 987 1494
rect 994 1492 1024 1544
rect 1058 1540 1059 1547
rect 1043 1532 1059 1540
rect 1030 1500 1043 1519
rect 1058 1500 1088 1516
rect 1030 1484 1104 1500
rect 1030 1482 1043 1484
rect 1058 1482 1092 1484
rect 695 1460 708 1462
rect 723 1460 757 1462
rect 695 1444 757 1460
rect 801 1455 817 1458
rect 879 1455 909 1466
rect 957 1462 1003 1478
rect 1030 1466 1104 1482
rect 957 1460 991 1462
rect 956 1444 1003 1460
rect 1030 1444 1043 1466
rect 1058 1444 1088 1466
rect 1115 1444 1116 1460
rect 1131 1444 1144 1604
rect 1174 1500 1187 1604
rect 1232 1582 1233 1592
rect 1248 1582 1261 1592
rect 1232 1578 1261 1582
rect 1266 1578 1296 1604
rect 1314 1590 1330 1592
rect 1402 1590 1455 1604
rect 1403 1588 1467 1590
rect 1510 1588 1525 1604
rect 1574 1601 1604 1604
rect 1574 1598 1610 1601
rect 1540 1590 1556 1592
rect 1314 1578 1329 1582
rect 1232 1576 1329 1578
rect 1357 1576 1525 1588
rect 1541 1578 1556 1582
rect 1574 1579 1613 1598
rect 1632 1592 1639 1593
rect 1638 1585 1639 1592
rect 1622 1582 1623 1585
rect 1638 1582 1651 1585
rect 1574 1578 1604 1579
rect 1613 1578 1619 1579
rect 1622 1578 1651 1582
rect 1541 1577 1651 1578
rect 1541 1576 1657 1577
rect 1216 1568 1267 1576
rect 1216 1556 1241 1568
rect 1248 1556 1267 1568
rect 1298 1568 1348 1576
rect 1298 1560 1314 1568
rect 1321 1566 1348 1568
rect 1357 1566 1578 1576
rect 1321 1556 1578 1566
rect 1607 1568 1657 1576
rect 1607 1559 1623 1568
rect 1216 1548 1267 1556
rect 1314 1548 1578 1556
rect 1604 1556 1623 1559
rect 1630 1556 1657 1568
rect 1604 1548 1657 1556
rect 1232 1540 1233 1548
rect 1248 1540 1261 1548
rect 1232 1532 1248 1540
rect 1229 1525 1248 1528
rect 1229 1516 1251 1525
rect 1202 1506 1251 1516
rect 1202 1500 1232 1506
rect 1251 1501 1256 1506
rect 1174 1484 1248 1500
rect 1266 1492 1296 1548
rect 1331 1538 1539 1548
rect 1574 1544 1619 1548
rect 1622 1547 1623 1548
rect 1638 1547 1651 1548
rect 1357 1508 1546 1538
rect 1372 1505 1546 1508
rect 1365 1502 1546 1505
rect 1174 1482 1187 1484
rect 1202 1482 1236 1484
rect 1174 1466 1248 1482
rect 1275 1478 1288 1492
rect 1303 1478 1319 1494
rect 1365 1489 1376 1502
rect 1158 1444 1159 1460
rect 1174 1444 1187 1466
rect 1202 1444 1232 1466
rect 1275 1462 1337 1478
rect 1365 1471 1376 1487
rect 1381 1482 1391 1502
rect 1401 1482 1415 1502
rect 1418 1489 1427 1502
rect 1443 1489 1452 1502
rect 1381 1471 1415 1482
rect 1418 1471 1427 1487
rect 1443 1471 1452 1487
rect 1459 1482 1469 1502
rect 1479 1482 1493 1502
rect 1494 1489 1505 1502
rect 1459 1471 1493 1482
rect 1494 1471 1505 1487
rect 1551 1478 1567 1494
rect 1574 1492 1604 1544
rect 1638 1540 1639 1547
rect 1623 1532 1639 1540
rect 1610 1500 1623 1519
rect 1638 1500 1668 1516
rect 1610 1484 1684 1500
rect 1610 1482 1623 1484
rect 1638 1482 1672 1484
rect 1275 1460 1288 1462
rect 1303 1460 1337 1462
rect 1275 1444 1337 1460
rect 1381 1455 1397 1458
rect 1459 1455 1489 1466
rect 1537 1462 1583 1478
rect 1610 1466 1684 1482
rect 1537 1460 1571 1462
rect 1536 1444 1583 1460
rect 1610 1444 1623 1466
rect 1638 1444 1668 1466
rect 1695 1444 1696 1460
rect 1711 1444 1724 1604
rect 1754 1500 1767 1604
rect 1812 1582 1813 1592
rect 1828 1582 1841 1592
rect 1812 1578 1841 1582
rect 1846 1578 1876 1604
rect 1894 1590 1910 1592
rect 1982 1590 2035 1604
rect 1983 1588 2047 1590
rect 2090 1588 2105 1604
rect 2154 1601 2184 1604
rect 2154 1598 2190 1601
rect 2120 1590 2136 1592
rect 1894 1578 1909 1582
rect 1812 1576 1909 1578
rect 1937 1576 2105 1588
rect 2121 1578 2136 1582
rect 2154 1579 2193 1598
rect 2212 1592 2219 1593
rect 2218 1585 2219 1592
rect 2202 1582 2203 1585
rect 2218 1582 2231 1585
rect 2154 1578 2184 1579
rect 2193 1578 2199 1579
rect 2202 1578 2231 1582
rect 2121 1577 2231 1578
rect 2121 1576 2237 1577
rect 1796 1568 1847 1576
rect 1796 1556 1821 1568
rect 1828 1556 1847 1568
rect 1878 1568 1928 1576
rect 1878 1560 1894 1568
rect 1901 1566 1928 1568
rect 1937 1566 2158 1576
rect 1901 1556 2158 1566
rect 2187 1568 2237 1576
rect 2187 1559 2203 1568
rect 1796 1548 1847 1556
rect 1894 1548 2158 1556
rect 2184 1556 2203 1559
rect 2210 1556 2237 1568
rect 2184 1548 2237 1556
rect 1812 1540 1813 1548
rect 1828 1540 1841 1548
rect 1812 1532 1828 1540
rect 1809 1525 1828 1528
rect 1809 1516 1831 1525
rect 1782 1506 1831 1516
rect 1782 1500 1812 1506
rect 1831 1501 1836 1506
rect 1754 1484 1828 1500
rect 1846 1492 1876 1548
rect 1911 1538 2119 1548
rect 2154 1544 2199 1548
rect 2202 1547 2203 1548
rect 2218 1547 2231 1548
rect 1937 1519 2126 1538
rect 1937 1508 2121 1519
rect 1952 1505 2121 1508
rect 1945 1502 2121 1505
rect 1754 1482 1767 1484
rect 1782 1482 1816 1484
rect 1754 1466 1828 1482
rect 1855 1478 1868 1492
rect 1883 1478 1899 1494
rect 1945 1489 1956 1502
rect 1738 1444 1739 1460
rect 1754 1444 1767 1466
rect 1782 1444 1812 1466
rect 1855 1462 1917 1478
rect 1945 1471 1956 1487
rect 1961 1482 1971 1502
rect 1981 1482 1995 1502
rect 1998 1489 2007 1502
rect 2023 1489 2032 1502
rect 1961 1471 1995 1482
rect 1998 1471 2007 1487
rect 2023 1471 2032 1487
rect 2039 1482 2049 1502
rect 2059 1482 2073 1502
rect 2074 1489 2085 1502
rect 2039 1471 2073 1482
rect 2074 1471 2085 1487
rect 2131 1478 2147 1494
rect 2154 1492 2184 1544
rect 2218 1540 2219 1547
rect 2203 1534 2219 1540
rect 2203 1532 2218 1534
rect 2190 1500 2203 1519
rect 2218 1500 2248 1516
rect 2190 1484 2264 1500
rect 2190 1482 2203 1484
rect 2218 1482 2252 1484
rect 1855 1460 1868 1462
rect 1883 1460 1917 1462
rect 1855 1444 1917 1460
rect 1961 1455 1977 1458
rect 2039 1455 2069 1466
rect 2117 1462 2163 1478
rect 2190 1466 2264 1482
rect 2117 1460 2151 1462
rect 2116 1444 2163 1460
rect 2190 1444 2203 1466
rect 2218 1444 2248 1466
rect 2275 1444 2276 1460
rect 2291 1444 2304 1604
rect 2334 1500 2347 1604
rect 2392 1582 2393 1592
rect 2408 1582 2421 1592
rect 2392 1578 2421 1582
rect 2426 1578 2456 1604
rect 2474 1590 2490 1592
rect 2562 1590 2615 1604
rect 2563 1588 2627 1590
rect 2670 1588 2685 1604
rect 2734 1601 2764 1604
rect 2734 1598 2770 1601
rect 2700 1590 2716 1592
rect 2474 1578 2489 1582
rect 2392 1576 2489 1578
rect 2517 1576 2685 1588
rect 2701 1578 2716 1582
rect 2734 1579 2773 1598
rect 2792 1592 2799 1593
rect 2798 1585 2799 1592
rect 2782 1582 2783 1585
rect 2798 1582 2811 1585
rect 2734 1578 2764 1579
rect 2773 1578 2779 1579
rect 2782 1578 2811 1582
rect 2701 1577 2811 1578
rect 2701 1576 2817 1577
rect 2376 1568 2427 1576
rect 2376 1556 2401 1568
rect 2408 1556 2427 1568
rect 2458 1568 2508 1576
rect 2458 1560 2474 1568
rect 2481 1566 2508 1568
rect 2517 1566 2738 1576
rect 2481 1556 2738 1566
rect 2767 1568 2817 1576
rect 2767 1559 2783 1568
rect 2376 1548 2427 1556
rect 2474 1548 2738 1556
rect 2764 1556 2783 1559
rect 2790 1556 2817 1568
rect 2764 1548 2817 1556
rect 2392 1540 2393 1548
rect 2408 1540 2421 1548
rect 2392 1534 2408 1540
rect 2393 1532 2408 1534
rect 2389 1525 2408 1528
rect 2389 1516 2411 1525
rect 2362 1506 2411 1516
rect 2362 1500 2392 1506
rect 2411 1501 2416 1506
rect 2334 1484 2408 1500
rect 2426 1492 2456 1548
rect 2491 1538 2699 1548
rect 2734 1544 2779 1548
rect 2782 1547 2783 1548
rect 2798 1547 2811 1548
rect 2517 1508 2706 1538
rect 2532 1505 2706 1508
rect 2525 1502 2706 1505
rect 2334 1482 2347 1484
rect 2362 1482 2396 1484
rect 2334 1466 2408 1482
rect 2435 1478 2448 1492
rect 2463 1478 2479 1494
rect 2525 1489 2536 1502
rect 2318 1444 2319 1460
rect 2334 1444 2347 1466
rect 2362 1444 2392 1466
rect 2435 1462 2497 1478
rect 2525 1471 2536 1487
rect 2541 1482 2551 1502
rect 2561 1482 2575 1502
rect 2578 1489 2587 1502
rect 2603 1489 2612 1502
rect 2541 1471 2575 1482
rect 2578 1471 2587 1487
rect 2603 1471 2612 1487
rect 2619 1482 2629 1502
rect 2639 1482 2653 1502
rect 2654 1489 2665 1502
rect 2619 1471 2653 1482
rect 2654 1471 2665 1487
rect 2711 1478 2727 1494
rect 2734 1492 2764 1544
rect 2798 1540 2799 1547
rect 2783 1532 2799 1540
rect 2770 1500 2783 1519
rect 2798 1500 2828 1516
rect 2770 1484 2844 1500
rect 2770 1482 2783 1484
rect 2798 1482 2832 1484
rect 2435 1460 2448 1462
rect 2463 1460 2497 1462
rect 2435 1444 2497 1460
rect 2541 1455 2557 1458
rect 2619 1455 2649 1466
rect 2697 1462 2743 1478
rect 2770 1466 2844 1482
rect 2697 1460 2731 1462
rect 2696 1444 2743 1460
rect 2770 1444 2783 1466
rect 2798 1444 2828 1466
rect 2855 1444 2856 1460
rect 2871 1444 2884 1604
rect 2914 1500 2927 1604
rect 2972 1582 2973 1592
rect 2988 1582 3001 1592
rect 2972 1578 3001 1582
rect 3006 1578 3036 1604
rect 3054 1590 3070 1592
rect 3142 1590 3195 1604
rect 3143 1588 3205 1590
rect 3250 1588 3265 1604
rect 3314 1601 3344 1604
rect 3314 1598 3350 1601
rect 3280 1590 3296 1592
rect 3054 1578 3069 1582
rect 2972 1576 3069 1578
rect 3097 1576 3265 1588
rect 3281 1578 3296 1582
rect 3314 1579 3353 1598
rect 3372 1592 3379 1593
rect 3378 1585 3379 1592
rect 3362 1582 3363 1585
rect 3378 1582 3391 1585
rect 3314 1578 3344 1579
rect 3353 1578 3359 1579
rect 3362 1578 3391 1582
rect 3281 1577 3391 1578
rect 3281 1576 3397 1577
rect 2956 1568 3007 1576
rect 2956 1556 2981 1568
rect 2988 1556 3007 1568
rect 3038 1568 3088 1576
rect 3038 1560 3054 1568
rect 3061 1566 3088 1568
rect 3097 1566 3318 1576
rect 3061 1556 3318 1566
rect 3347 1568 3397 1576
rect 3347 1559 3363 1568
rect 2956 1548 3007 1556
rect 3054 1548 3318 1556
rect 3344 1556 3363 1559
rect 3370 1556 3397 1568
rect 3344 1548 3397 1556
rect 2972 1540 2973 1548
rect 2988 1540 3001 1548
rect 2972 1532 2988 1540
rect 2969 1525 2988 1528
rect 2969 1516 2991 1525
rect 2942 1506 2991 1516
rect 2942 1500 2972 1506
rect 2991 1501 2996 1506
rect 2914 1484 2988 1500
rect 3006 1492 3036 1548
rect 3071 1538 3279 1548
rect 3314 1544 3359 1548
rect 3362 1547 3363 1548
rect 3378 1547 3391 1548
rect 3097 1508 3286 1538
rect 3112 1505 3286 1508
rect 3105 1502 3286 1505
rect 2914 1482 2927 1484
rect 2942 1482 2976 1484
rect 2914 1466 2988 1482
rect 3015 1478 3028 1492
rect 3043 1478 3059 1494
rect 3105 1489 3116 1502
rect 2898 1444 2899 1460
rect 2914 1444 2927 1466
rect 2942 1444 2972 1466
rect 3015 1462 3077 1478
rect 3105 1471 3116 1487
rect 3121 1482 3131 1502
rect 3141 1482 3155 1502
rect 3158 1489 3167 1502
rect 3183 1489 3192 1502
rect 3121 1471 3155 1482
rect 3158 1471 3167 1487
rect 3183 1471 3192 1487
rect 3199 1482 3209 1502
rect 3219 1482 3233 1502
rect 3234 1489 3245 1502
rect 3199 1471 3233 1482
rect 3234 1471 3245 1487
rect 3291 1478 3307 1494
rect 3314 1492 3344 1544
rect 3378 1540 3379 1547
rect 3363 1532 3379 1540
rect 3350 1500 3363 1519
rect 3378 1500 3408 1516
rect 3350 1484 3424 1500
rect 3350 1482 3363 1484
rect 3378 1482 3412 1484
rect 3015 1460 3028 1462
rect 3043 1460 3077 1462
rect 3015 1444 3077 1460
rect 3121 1455 3137 1458
rect 3199 1455 3229 1466
rect 3277 1462 3323 1478
rect 3350 1466 3424 1482
rect 3277 1460 3311 1462
rect 3276 1444 3323 1460
rect 3350 1444 3363 1466
rect 3378 1444 3408 1466
rect 3435 1444 3436 1460
rect 3451 1444 3464 1604
rect 3494 1500 3507 1604
rect 3552 1582 3553 1592
rect 3568 1582 3581 1592
rect 3552 1578 3581 1582
rect 3586 1578 3616 1604
rect 3634 1590 3650 1592
rect 3722 1590 3775 1604
rect 3723 1588 3787 1590
rect 3830 1588 3845 1604
rect 3894 1601 3924 1604
rect 3894 1598 3930 1601
rect 3860 1590 3876 1592
rect 3634 1578 3649 1582
rect 3552 1576 3649 1578
rect 3677 1576 3845 1588
rect 3861 1578 3876 1582
rect 3894 1579 3933 1598
rect 3952 1592 3959 1593
rect 3958 1585 3959 1592
rect 3942 1582 3943 1585
rect 3958 1582 3971 1585
rect 3894 1578 3924 1579
rect 3933 1578 3939 1579
rect 3942 1578 3971 1582
rect 3861 1577 3971 1578
rect 3861 1576 3977 1577
rect 3536 1568 3587 1576
rect 3536 1556 3561 1568
rect 3568 1556 3587 1568
rect 3618 1568 3668 1576
rect 3618 1560 3634 1568
rect 3641 1566 3668 1568
rect 3677 1566 3898 1576
rect 3641 1556 3898 1566
rect 3927 1568 3977 1576
rect 3927 1559 3943 1568
rect 3536 1548 3587 1556
rect 3634 1548 3898 1556
rect 3924 1556 3943 1559
rect 3950 1556 3977 1568
rect 3924 1548 3977 1556
rect 3552 1540 3553 1548
rect 3568 1540 3581 1548
rect 3552 1532 3568 1540
rect 3549 1525 3568 1528
rect 3549 1516 3571 1525
rect 3522 1506 3571 1516
rect 3522 1500 3552 1506
rect 3571 1501 3576 1506
rect 3494 1484 3568 1500
rect 3586 1492 3616 1548
rect 3651 1538 3859 1548
rect 3894 1544 3939 1548
rect 3942 1547 3943 1548
rect 3958 1547 3971 1548
rect 3677 1508 3866 1538
rect 3692 1505 3866 1508
rect 3685 1502 3866 1505
rect 3494 1482 3507 1484
rect 3522 1482 3556 1484
rect 3494 1466 3568 1482
rect 3595 1478 3608 1492
rect 3623 1478 3639 1494
rect 3685 1489 3696 1502
rect 3478 1444 3479 1460
rect 3494 1444 3507 1466
rect 3522 1444 3552 1466
rect 3595 1462 3657 1478
rect 3685 1471 3696 1487
rect 3701 1482 3711 1502
rect 3721 1482 3735 1502
rect 3738 1489 3747 1502
rect 3763 1489 3772 1502
rect 3701 1471 3735 1482
rect 3738 1471 3747 1487
rect 3763 1471 3772 1487
rect 3779 1482 3789 1502
rect 3799 1482 3813 1502
rect 3814 1489 3825 1502
rect 3779 1471 3813 1482
rect 3814 1471 3825 1487
rect 3871 1478 3887 1494
rect 3894 1492 3924 1544
rect 3958 1540 3959 1547
rect 3943 1532 3959 1540
rect 3930 1500 3943 1519
rect 3958 1500 3988 1516
rect 3930 1484 4004 1500
rect 3930 1482 3943 1484
rect 3958 1482 3992 1484
rect 3595 1460 3608 1462
rect 3623 1460 3657 1462
rect 3595 1444 3657 1460
rect 3701 1455 3717 1458
rect 3779 1455 3809 1466
rect 3857 1462 3903 1478
rect 3930 1466 4004 1482
rect 3857 1460 3891 1462
rect 3856 1444 3903 1460
rect 3930 1444 3943 1466
rect 3958 1444 3988 1466
rect 4015 1444 4016 1460
rect 4031 1444 4044 1604
rect 4074 1500 4087 1604
rect 4132 1582 4133 1592
rect 4148 1582 4161 1592
rect 4132 1578 4161 1582
rect 4166 1578 4196 1604
rect 4214 1590 4230 1592
rect 4302 1590 4355 1604
rect 4303 1588 4367 1590
rect 4410 1588 4425 1604
rect 4474 1601 4504 1604
rect 4474 1598 4510 1601
rect 4440 1590 4456 1592
rect 4214 1578 4229 1582
rect 4132 1576 4229 1578
rect 4257 1576 4425 1588
rect 4441 1578 4456 1582
rect 4474 1579 4513 1598
rect 4532 1592 4539 1593
rect 4538 1585 4539 1592
rect 4522 1582 4523 1585
rect 4538 1582 4551 1585
rect 4474 1578 4504 1579
rect 4513 1578 4519 1579
rect 4522 1578 4551 1582
rect 4441 1577 4551 1578
rect 4441 1576 4557 1577
rect 4116 1568 4167 1576
rect 4116 1556 4141 1568
rect 4148 1556 4167 1568
rect 4198 1568 4248 1576
rect 4198 1560 4214 1568
rect 4221 1566 4248 1568
rect 4257 1566 4478 1576
rect 4221 1556 4478 1566
rect 4507 1568 4557 1576
rect 4507 1559 4523 1568
rect 4116 1548 4167 1556
rect 4214 1548 4478 1556
rect 4504 1556 4523 1559
rect 4530 1556 4557 1568
rect 4504 1548 4557 1556
rect 4132 1540 4133 1548
rect 4148 1540 4161 1548
rect 4132 1532 4148 1540
rect 4129 1525 4148 1528
rect 4129 1516 4151 1525
rect 4102 1506 4151 1516
rect 4102 1500 4132 1506
rect 4151 1501 4156 1506
rect 4074 1484 4148 1500
rect 4166 1492 4196 1548
rect 4231 1538 4439 1548
rect 4474 1544 4519 1548
rect 4522 1547 4523 1548
rect 4538 1547 4551 1548
rect 4257 1508 4446 1538
rect 4272 1505 4446 1508
rect 4265 1502 4446 1505
rect 4074 1482 4087 1484
rect 4102 1482 4136 1484
rect 4074 1466 4148 1482
rect 4175 1478 4188 1492
rect 4203 1478 4219 1494
rect 4265 1489 4276 1502
rect 4058 1444 4059 1460
rect 4074 1444 4087 1466
rect 4102 1444 4132 1466
rect 4175 1462 4237 1478
rect 4265 1471 4276 1487
rect 4281 1482 4291 1502
rect 4301 1482 4315 1502
rect 4318 1489 4327 1502
rect 4343 1489 4352 1502
rect 4281 1471 4315 1482
rect 4318 1471 4327 1487
rect 4343 1471 4352 1487
rect 4359 1482 4369 1502
rect 4379 1482 4393 1502
rect 4394 1489 4405 1502
rect 4359 1471 4393 1482
rect 4394 1471 4405 1487
rect 4451 1478 4467 1494
rect 4474 1492 4504 1544
rect 4538 1540 4539 1547
rect 4523 1532 4539 1540
rect 4510 1500 4523 1519
rect 4538 1500 4568 1516
rect 4510 1484 4584 1500
rect 4510 1482 4523 1484
rect 4538 1482 4572 1484
rect 4175 1460 4188 1462
rect 4203 1460 4237 1462
rect 4175 1444 4237 1460
rect 4281 1455 4297 1458
rect 4359 1455 4389 1466
rect 4437 1462 4483 1478
rect 4510 1466 4584 1482
rect 4437 1460 4471 1462
rect 4436 1444 4483 1460
rect 4510 1444 4523 1466
rect 4538 1444 4568 1466
rect 4595 1444 4596 1460
rect 4611 1444 4624 1604
rect 4654 1500 4667 1604
rect 4712 1582 4713 1592
rect 4733 1590 4741 1592
rect 4731 1588 4741 1590
rect 4729 1586 4741 1588
rect 4728 1582 4741 1586
rect 4712 1578 4741 1582
rect 4746 1578 4776 1604
rect 4794 1590 4810 1592
rect 4882 1590 4933 1604
rect 4883 1588 4947 1590
rect 4990 1588 5005 1604
rect 5054 1601 5084 1604
rect 5054 1598 5090 1601
rect 5020 1590 5036 1592
rect 4794 1578 4809 1582
rect 4712 1576 4809 1578
rect 4837 1576 5005 1588
rect 5021 1578 5036 1582
rect 5054 1579 5093 1598
rect 5112 1592 5119 1593
rect 5118 1585 5119 1592
rect 5102 1582 5103 1585
rect 5118 1582 5131 1585
rect 5054 1578 5084 1579
rect 5093 1578 5099 1579
rect 5102 1578 5131 1582
rect 5021 1577 5131 1578
rect 5021 1576 5137 1577
rect 4696 1568 4747 1576
rect 4696 1556 4721 1568
rect 4728 1556 4747 1568
rect 4778 1568 4828 1576
rect 4778 1560 4794 1568
rect 4801 1566 4828 1568
rect 4837 1566 5058 1576
rect 4801 1556 5058 1566
rect 5087 1568 5137 1576
rect 5087 1559 5103 1568
rect 4696 1548 4747 1556
rect 4794 1548 5058 1556
rect 5084 1556 5103 1559
rect 5110 1556 5137 1568
rect 5084 1548 5137 1556
rect 4712 1540 4713 1548
rect 4728 1540 4741 1548
rect 4712 1532 4728 1540
rect 4709 1525 4728 1528
rect 4709 1516 4731 1525
rect 4682 1506 4731 1516
rect 4682 1500 4712 1506
rect 4731 1501 4736 1506
rect 4654 1484 4728 1500
rect 4746 1492 4776 1548
rect 4811 1538 5019 1548
rect 5054 1544 5099 1548
rect 5102 1547 5103 1548
rect 5118 1547 5131 1548
rect 4837 1508 5026 1538
rect 4852 1505 5026 1508
rect 4845 1502 5026 1505
rect 4654 1482 4667 1484
rect 4682 1482 4716 1484
rect 4654 1466 4728 1482
rect 4755 1478 4768 1492
rect 4783 1478 4799 1494
rect 4845 1489 4856 1502
rect 4638 1444 4639 1460
rect 4654 1444 4667 1466
rect 4682 1444 4712 1466
rect 4755 1462 4817 1478
rect 4845 1471 4856 1487
rect 4861 1482 4871 1502
rect 4881 1482 4895 1502
rect 4898 1489 4907 1502
rect 4923 1489 4932 1502
rect 4861 1471 4895 1482
rect 4898 1471 4907 1487
rect 4923 1471 4932 1487
rect 4939 1482 4949 1502
rect 4959 1482 4973 1502
rect 4974 1489 4985 1502
rect 4939 1471 4973 1482
rect 4974 1471 4985 1487
rect 5031 1478 5047 1494
rect 5054 1492 5084 1544
rect 5118 1540 5119 1547
rect 5103 1532 5119 1540
rect 5090 1500 5103 1519
rect 5118 1500 5148 1516
rect 5090 1484 5164 1500
rect 5090 1482 5103 1484
rect 5118 1482 5152 1484
rect 4755 1460 4768 1462
rect 4783 1460 4817 1462
rect 4755 1444 4817 1460
rect 4861 1455 4877 1458
rect 4939 1455 4969 1466
rect 5017 1462 5063 1478
rect 5090 1466 5164 1482
rect 5017 1460 5051 1462
rect 5016 1444 5063 1460
rect 5090 1444 5103 1466
rect 5118 1444 5148 1466
rect 5175 1444 5176 1460
rect 5191 1444 5204 1604
rect 5234 1500 5247 1604
rect 5292 1582 5293 1592
rect 5313 1590 5321 1592
rect 5311 1588 5321 1590
rect 5309 1586 5321 1588
rect 5308 1582 5321 1586
rect 5292 1578 5321 1582
rect 5326 1578 5356 1604
rect 5374 1590 5390 1592
rect 5462 1590 5513 1604
rect 5463 1588 5527 1590
rect 5570 1588 5585 1604
rect 5634 1601 5664 1604
rect 5634 1598 5670 1601
rect 5600 1590 5616 1592
rect 5374 1578 5389 1582
rect 5292 1576 5389 1578
rect 5417 1576 5585 1588
rect 5601 1578 5616 1582
rect 5634 1579 5673 1598
rect 5692 1592 5699 1593
rect 5698 1585 5699 1592
rect 5682 1582 5683 1585
rect 5698 1582 5711 1585
rect 5634 1578 5664 1579
rect 5673 1578 5679 1579
rect 5682 1578 5711 1582
rect 5601 1577 5711 1578
rect 5601 1576 5717 1577
rect 5276 1568 5327 1576
rect 5276 1556 5301 1568
rect 5308 1556 5327 1568
rect 5358 1568 5408 1576
rect 5358 1560 5374 1568
rect 5381 1566 5408 1568
rect 5417 1566 5638 1576
rect 5381 1556 5638 1566
rect 5667 1568 5717 1576
rect 5667 1559 5683 1568
rect 5276 1548 5327 1556
rect 5374 1548 5638 1556
rect 5664 1556 5683 1559
rect 5690 1556 5717 1568
rect 5664 1548 5717 1556
rect 5292 1540 5293 1548
rect 5308 1540 5321 1548
rect 5292 1532 5308 1540
rect 5289 1525 5308 1528
rect 5289 1516 5311 1525
rect 5262 1506 5311 1516
rect 5262 1500 5292 1506
rect 5311 1501 5316 1506
rect 5234 1484 5308 1500
rect 5326 1492 5356 1548
rect 5391 1538 5599 1548
rect 5634 1544 5679 1548
rect 5682 1547 5683 1548
rect 5698 1547 5711 1548
rect 5417 1508 5606 1538
rect 5432 1505 5606 1508
rect 5425 1502 5606 1505
rect 5234 1482 5247 1484
rect 5262 1482 5296 1484
rect 5234 1466 5308 1482
rect 5335 1478 5348 1492
rect 5363 1478 5379 1494
rect 5425 1489 5436 1502
rect 5218 1444 5219 1460
rect 5234 1444 5247 1466
rect 5262 1444 5292 1466
rect 5335 1462 5397 1478
rect 5425 1471 5436 1487
rect 5441 1482 5451 1502
rect 5461 1482 5475 1502
rect 5478 1489 5487 1502
rect 5503 1489 5512 1502
rect 5441 1471 5475 1482
rect 5478 1471 5487 1487
rect 5503 1471 5512 1487
rect 5519 1482 5529 1502
rect 5539 1482 5553 1502
rect 5554 1489 5565 1502
rect 5519 1471 5553 1482
rect 5554 1471 5565 1487
rect 5611 1478 5627 1494
rect 5634 1492 5664 1544
rect 5698 1540 5699 1547
rect 5683 1532 5699 1540
rect 5670 1500 5683 1519
rect 5698 1500 5728 1516
rect 5670 1484 5744 1500
rect 5670 1482 5683 1484
rect 5698 1482 5732 1484
rect 5335 1460 5348 1462
rect 5363 1460 5397 1462
rect 5335 1444 5397 1460
rect 5441 1455 5457 1458
rect 5519 1455 5549 1466
rect 5597 1462 5643 1478
rect 5670 1466 5744 1482
rect 5597 1460 5631 1462
rect 5596 1444 5643 1460
rect 5670 1444 5683 1466
rect 5698 1444 5728 1466
rect 5755 1444 5756 1460
rect 5771 1444 5784 1604
rect 5814 1500 5827 1604
rect 5872 1582 5873 1592
rect 5893 1590 5901 1592
rect 5891 1588 5901 1590
rect 5889 1586 5901 1588
rect 5888 1582 5901 1586
rect 5872 1578 5901 1582
rect 5906 1578 5936 1604
rect 5954 1590 5970 1592
rect 6042 1590 6093 1604
rect 6043 1588 6107 1590
rect 6150 1588 6165 1604
rect 6214 1601 6244 1604
rect 6214 1598 6250 1601
rect 6180 1590 6196 1592
rect 5954 1578 5969 1582
rect 5872 1576 5969 1578
rect 5997 1576 6165 1588
rect 6181 1578 6196 1582
rect 6214 1579 6253 1598
rect 6272 1592 6279 1593
rect 6278 1585 6279 1592
rect 6262 1582 6263 1585
rect 6278 1582 6291 1585
rect 6214 1578 6244 1579
rect 6253 1578 6259 1579
rect 6262 1578 6291 1582
rect 6181 1577 6291 1578
rect 6181 1576 6297 1577
rect 5856 1568 5907 1576
rect 5856 1556 5881 1568
rect 5888 1556 5907 1568
rect 5938 1568 5988 1576
rect 5938 1560 5954 1568
rect 5961 1566 5988 1568
rect 5997 1566 6218 1576
rect 5961 1556 6218 1566
rect 6247 1568 6297 1576
rect 6247 1559 6263 1568
rect 5856 1548 5907 1556
rect 5954 1548 6218 1556
rect 6244 1556 6263 1559
rect 6270 1556 6297 1568
rect 6244 1548 6297 1556
rect 5872 1540 5873 1548
rect 5888 1540 5901 1548
rect 5872 1532 5888 1540
rect 5869 1525 5888 1528
rect 5869 1516 5891 1525
rect 5842 1506 5891 1516
rect 5842 1500 5872 1506
rect 5891 1501 5896 1506
rect 5814 1484 5888 1500
rect 5906 1492 5936 1548
rect 5971 1538 6179 1548
rect 6214 1544 6259 1548
rect 6262 1547 6263 1548
rect 6278 1547 6291 1548
rect 5997 1508 6186 1538
rect 6012 1505 6186 1508
rect 6005 1502 6186 1505
rect 5814 1482 5827 1484
rect 5842 1482 5876 1484
rect 5814 1466 5888 1482
rect 5915 1478 5928 1492
rect 5943 1478 5959 1494
rect 6005 1489 6016 1502
rect 5798 1444 5799 1460
rect 5814 1444 5827 1466
rect 5842 1444 5872 1466
rect 5915 1462 5977 1478
rect 6005 1471 6016 1487
rect 6021 1482 6031 1502
rect 6041 1482 6055 1502
rect 6058 1489 6067 1502
rect 6083 1489 6092 1502
rect 6021 1471 6055 1482
rect 6058 1471 6067 1487
rect 6083 1471 6092 1487
rect 6099 1482 6109 1502
rect 6119 1482 6133 1502
rect 6134 1489 6145 1502
rect 6099 1471 6133 1482
rect 6134 1471 6145 1487
rect 6191 1478 6207 1494
rect 6214 1492 6244 1544
rect 6278 1540 6279 1547
rect 6263 1532 6279 1540
rect 6250 1500 6263 1519
rect 6278 1500 6308 1516
rect 6250 1484 6324 1500
rect 6250 1482 6263 1484
rect 6278 1482 6312 1484
rect 5915 1460 5928 1462
rect 5943 1460 5977 1462
rect 5915 1444 5977 1460
rect 6021 1455 6037 1458
rect 6099 1455 6129 1466
rect 6177 1462 6223 1478
rect 6250 1466 6324 1482
rect 6177 1460 6211 1462
rect 6176 1444 6223 1460
rect 6250 1444 6263 1466
rect 6278 1444 6308 1466
rect 6335 1444 6336 1460
rect 6351 1444 6364 1604
rect 6394 1500 6407 1604
rect 6452 1582 6453 1592
rect 6473 1590 6481 1592
rect 6471 1588 6481 1590
rect 6469 1586 6481 1588
rect 6468 1582 6481 1586
rect 6452 1578 6481 1582
rect 6486 1578 6516 1604
rect 6534 1590 6550 1592
rect 6622 1590 6673 1604
rect 6623 1588 6687 1590
rect 6730 1588 6745 1604
rect 6794 1601 6824 1604
rect 6794 1598 6830 1601
rect 6760 1590 6776 1592
rect 6534 1578 6549 1582
rect 6452 1576 6549 1578
rect 6577 1576 6745 1588
rect 6761 1578 6776 1582
rect 6794 1579 6833 1598
rect 6852 1592 6859 1593
rect 6858 1585 6859 1592
rect 6842 1582 6843 1585
rect 6858 1582 6871 1585
rect 6794 1578 6824 1579
rect 6833 1578 6839 1579
rect 6842 1578 6871 1582
rect 6761 1577 6871 1578
rect 6761 1576 6877 1577
rect 6436 1568 6487 1576
rect 6436 1556 6461 1568
rect 6468 1556 6487 1568
rect 6518 1568 6568 1576
rect 6518 1560 6534 1568
rect 6541 1566 6568 1568
rect 6577 1566 6798 1576
rect 6541 1556 6798 1566
rect 6827 1568 6877 1576
rect 6827 1559 6843 1568
rect 6436 1548 6487 1556
rect 6534 1548 6798 1556
rect 6824 1556 6843 1559
rect 6850 1556 6877 1568
rect 6824 1548 6877 1556
rect 6452 1540 6453 1548
rect 6468 1540 6481 1548
rect 6452 1532 6468 1540
rect 6449 1525 6468 1528
rect 6449 1516 6471 1525
rect 6422 1506 6471 1516
rect 6422 1500 6452 1506
rect 6471 1501 6476 1506
rect 6394 1484 6468 1500
rect 6486 1492 6516 1548
rect 6551 1538 6759 1548
rect 6794 1544 6839 1548
rect 6842 1547 6843 1548
rect 6858 1547 6871 1548
rect 6577 1508 6766 1538
rect 6592 1505 6766 1508
rect 6585 1502 6766 1505
rect 6394 1482 6407 1484
rect 6422 1482 6456 1484
rect 6394 1466 6468 1482
rect 6495 1478 6508 1492
rect 6523 1478 6539 1494
rect 6585 1489 6596 1502
rect 6378 1444 6379 1460
rect 6394 1444 6407 1466
rect 6422 1444 6452 1466
rect 6495 1462 6557 1478
rect 6585 1471 6596 1487
rect 6601 1482 6611 1502
rect 6621 1482 6635 1502
rect 6638 1489 6647 1502
rect 6663 1489 6672 1502
rect 6601 1471 6635 1482
rect 6638 1471 6647 1487
rect 6663 1471 6672 1487
rect 6679 1482 6689 1502
rect 6699 1482 6713 1502
rect 6714 1489 6725 1502
rect 6679 1471 6713 1482
rect 6714 1471 6725 1487
rect 6771 1478 6787 1494
rect 6794 1492 6824 1544
rect 6858 1540 6859 1547
rect 6843 1532 6859 1540
rect 6830 1500 6843 1519
rect 6858 1500 6888 1516
rect 6830 1484 6904 1500
rect 6830 1482 6843 1484
rect 6858 1482 6892 1484
rect 6495 1460 6508 1462
rect 6523 1460 6557 1462
rect 6495 1444 6557 1460
rect 6601 1455 6617 1458
rect 6679 1455 6709 1466
rect 6757 1462 6803 1478
rect 6830 1466 6904 1482
rect 6757 1460 6791 1462
rect 6756 1444 6803 1460
rect 6830 1444 6843 1466
rect 6858 1444 6888 1466
rect 6915 1444 6916 1460
rect 6931 1444 6944 1604
rect 0 1436 33 1444
rect 0 1410 7 1436
rect 14 1410 33 1436
rect 97 1432 159 1444
rect 171 1432 246 1444
rect 304 1432 379 1444
rect 391 1432 422 1444
rect 428 1432 463 1444
rect 97 1430 259 1432
rect 0 1402 33 1410
rect 115 1406 128 1430
rect 143 1428 158 1430
rect 14 1392 27 1402
rect 42 1392 72 1406
rect 115 1392 158 1406
rect 182 1403 189 1410
rect 192 1406 259 1430
rect 291 1430 463 1432
rect 261 1408 289 1412
rect 291 1408 371 1430
rect 392 1428 407 1430
rect 261 1406 371 1408
rect 192 1402 371 1406
rect 165 1392 195 1402
rect 197 1392 350 1402
rect 358 1392 388 1402
rect 392 1392 422 1406
rect 450 1392 463 1430
rect 535 1436 570 1444
rect 535 1410 536 1436
rect 543 1410 570 1436
rect 478 1392 508 1406
rect 535 1402 570 1410
rect 572 1436 613 1444
rect 572 1410 587 1436
rect 594 1410 613 1436
rect 677 1432 739 1444
rect 751 1432 826 1444
rect 884 1432 959 1444
rect 971 1432 1002 1444
rect 1008 1432 1043 1444
rect 677 1430 839 1432
rect 572 1402 613 1410
rect 695 1406 708 1430
rect 723 1428 738 1430
rect 535 1392 536 1402
rect 551 1392 564 1402
rect 578 1392 579 1402
rect 594 1392 607 1402
rect 622 1392 652 1406
rect 695 1392 738 1406
rect 762 1403 769 1410
rect 772 1406 839 1430
rect 871 1430 1043 1432
rect 841 1408 869 1412
rect 871 1408 951 1430
rect 972 1428 987 1430
rect 841 1406 951 1408
rect 772 1402 951 1406
rect 745 1392 775 1402
rect 777 1392 930 1402
rect 938 1392 968 1402
rect 972 1392 1002 1406
rect 1030 1392 1043 1430
rect 1115 1436 1150 1444
rect 1115 1410 1116 1436
rect 1123 1410 1150 1436
rect 1058 1392 1088 1406
rect 1115 1402 1150 1410
rect 1152 1436 1193 1444
rect 1152 1410 1167 1436
rect 1174 1410 1193 1436
rect 1257 1432 1319 1444
rect 1331 1432 1406 1444
rect 1464 1432 1539 1444
rect 1551 1432 1582 1444
rect 1588 1432 1623 1444
rect 1257 1430 1419 1432
rect 1152 1402 1193 1410
rect 1275 1406 1288 1430
rect 1303 1428 1318 1430
rect 1115 1392 1116 1402
rect 1131 1392 1144 1402
rect 1158 1392 1159 1402
rect 1174 1392 1187 1402
rect 1202 1392 1232 1406
rect 1275 1392 1318 1406
rect 1342 1403 1349 1410
rect 1352 1406 1419 1430
rect 1451 1430 1623 1432
rect 1421 1408 1449 1412
rect 1451 1408 1531 1430
rect 1552 1428 1567 1430
rect 1421 1406 1531 1408
rect 1352 1402 1531 1406
rect 1325 1392 1355 1402
rect 1357 1392 1510 1402
rect 1518 1392 1548 1402
rect 1552 1392 1582 1406
rect 1610 1392 1623 1430
rect 1695 1436 1730 1444
rect 1695 1410 1696 1436
rect 1703 1410 1730 1436
rect 1638 1392 1668 1406
rect 1695 1402 1730 1410
rect 1732 1436 1773 1444
rect 1732 1410 1747 1436
rect 1754 1410 1773 1436
rect 1837 1432 1899 1444
rect 1911 1432 1986 1444
rect 2044 1432 2119 1444
rect 2131 1432 2162 1444
rect 2168 1432 2203 1444
rect 1837 1430 1999 1432
rect 1732 1402 1773 1410
rect 1855 1406 1868 1430
rect 1883 1428 1898 1430
rect 1695 1392 1696 1402
rect 1711 1392 1724 1402
rect 1738 1392 1739 1402
rect 1754 1392 1767 1402
rect 1782 1392 1812 1406
rect 1855 1392 1898 1406
rect 1922 1403 1929 1410
rect 1932 1406 1999 1430
rect 2031 1430 2203 1432
rect 2001 1408 2029 1412
rect 2031 1408 2111 1430
rect 2132 1428 2147 1430
rect 2001 1406 2111 1408
rect 1932 1402 2111 1406
rect 1905 1392 1935 1402
rect 1937 1392 2090 1402
rect 2098 1392 2128 1402
rect 2132 1392 2162 1406
rect 2190 1392 2203 1430
rect 2275 1436 2310 1444
rect 2275 1410 2276 1436
rect 2283 1410 2310 1436
rect 2218 1392 2248 1406
rect 2275 1402 2310 1410
rect 2312 1436 2353 1444
rect 2312 1410 2327 1436
rect 2334 1410 2353 1436
rect 2417 1432 2479 1444
rect 2491 1432 2566 1444
rect 2624 1432 2699 1444
rect 2711 1432 2742 1444
rect 2748 1432 2783 1444
rect 2417 1430 2579 1432
rect 2312 1402 2353 1410
rect 2435 1406 2448 1430
rect 2463 1428 2478 1430
rect 2275 1392 2276 1402
rect 2291 1392 2304 1402
rect 2318 1392 2319 1402
rect 2334 1392 2347 1402
rect 2362 1392 2392 1406
rect 2435 1392 2478 1406
rect 2502 1403 2509 1410
rect 2512 1406 2579 1430
rect 2611 1430 2783 1432
rect 2581 1408 2609 1412
rect 2611 1408 2691 1430
rect 2712 1428 2727 1430
rect 2581 1406 2691 1408
rect 2512 1402 2691 1406
rect 2485 1392 2515 1402
rect 2517 1392 2670 1402
rect 2678 1392 2708 1402
rect 2712 1392 2742 1406
rect 2770 1392 2783 1430
rect 2855 1436 2890 1444
rect 2855 1410 2856 1436
rect 2863 1410 2890 1436
rect 2798 1392 2828 1406
rect 2855 1402 2890 1410
rect 2892 1436 2933 1444
rect 2892 1410 2907 1436
rect 2914 1410 2933 1436
rect 2997 1432 3059 1444
rect 3071 1432 3146 1444
rect 3204 1432 3279 1444
rect 3291 1432 3322 1444
rect 3328 1432 3363 1444
rect 2997 1430 3159 1432
rect 2892 1402 2933 1410
rect 3015 1406 3028 1430
rect 3043 1428 3058 1430
rect 2855 1392 2856 1402
rect 2871 1392 2884 1402
rect 2898 1392 2899 1402
rect 2914 1392 2927 1402
rect 2942 1392 2972 1406
rect 3015 1392 3058 1406
rect 3082 1403 3089 1410
rect 3092 1406 3159 1430
rect 3191 1430 3363 1432
rect 3161 1408 3189 1412
rect 3191 1408 3271 1430
rect 3292 1428 3307 1430
rect 3161 1406 3271 1408
rect 3092 1402 3271 1406
rect 3065 1392 3095 1402
rect 3097 1392 3250 1402
rect 3258 1392 3288 1402
rect 3292 1392 3322 1406
rect 3350 1392 3363 1430
rect 3435 1436 3470 1444
rect 3435 1410 3436 1436
rect 3443 1410 3470 1436
rect 3378 1392 3408 1406
rect 3435 1402 3470 1410
rect 3472 1436 3513 1444
rect 3472 1410 3487 1436
rect 3494 1410 3513 1436
rect 3577 1432 3639 1444
rect 3651 1432 3726 1444
rect 3784 1432 3859 1444
rect 3871 1432 3902 1444
rect 3908 1432 3943 1444
rect 3577 1430 3739 1432
rect 3472 1402 3513 1410
rect 3595 1406 3608 1430
rect 3623 1428 3638 1430
rect 3435 1392 3436 1402
rect 3451 1392 3464 1402
rect 3478 1392 3479 1402
rect 3494 1392 3507 1402
rect 3522 1392 3552 1406
rect 3595 1392 3638 1406
rect 3662 1403 3669 1410
rect 3672 1406 3739 1430
rect 3771 1430 3943 1432
rect 3741 1408 3769 1412
rect 3771 1408 3851 1430
rect 3872 1428 3887 1430
rect 3741 1406 3851 1408
rect 3672 1402 3851 1406
rect 3645 1392 3675 1402
rect 3677 1392 3830 1402
rect 3838 1392 3868 1402
rect 3872 1392 3902 1406
rect 3930 1392 3943 1430
rect 4015 1436 4050 1444
rect 4015 1410 4016 1436
rect 4023 1410 4050 1436
rect 3958 1392 3988 1406
rect 4015 1402 4050 1410
rect 4052 1436 4093 1444
rect 4052 1410 4067 1436
rect 4074 1410 4093 1436
rect 4157 1432 4219 1444
rect 4231 1432 4306 1444
rect 4364 1432 4439 1444
rect 4451 1432 4482 1444
rect 4488 1432 4523 1444
rect 4157 1430 4319 1432
rect 4052 1402 4093 1410
rect 4175 1406 4188 1430
rect 4203 1428 4218 1430
rect 4015 1392 4016 1402
rect 4031 1392 4044 1402
rect 4058 1392 4059 1402
rect 4074 1392 4087 1402
rect 4102 1392 4132 1406
rect 4175 1392 4218 1406
rect 4242 1403 4249 1410
rect 4252 1406 4319 1430
rect 4351 1430 4523 1432
rect 4321 1408 4349 1412
rect 4351 1408 4431 1430
rect 4452 1428 4467 1430
rect 4321 1406 4431 1408
rect 4252 1402 4431 1406
rect 4225 1392 4255 1402
rect 4257 1392 4410 1402
rect 4418 1392 4448 1402
rect 4452 1392 4482 1406
rect 4510 1392 4523 1430
rect 4595 1436 4630 1444
rect 4595 1410 4596 1436
rect 4603 1410 4630 1436
rect 4538 1392 4568 1406
rect 4595 1402 4630 1410
rect 4632 1436 4673 1444
rect 4632 1410 4647 1436
rect 4654 1410 4673 1436
rect 4737 1432 4799 1444
rect 4811 1432 4886 1444
rect 4944 1432 5019 1444
rect 5031 1432 5062 1444
rect 5068 1432 5103 1444
rect 4737 1430 4899 1432
rect 4632 1402 4673 1410
rect 4755 1406 4768 1430
rect 4783 1428 4798 1430
rect 4832 1412 4899 1430
rect 4931 1430 5103 1432
rect 4931 1412 5011 1430
rect 5032 1428 5047 1430
rect 4595 1392 4596 1402
rect 4611 1392 4624 1402
rect 4638 1392 4639 1402
rect 4654 1392 4667 1402
rect 4682 1392 4712 1406
rect 4755 1392 4798 1406
rect 4822 1403 4829 1410
rect 4832 1402 5011 1412
rect 4805 1392 4835 1402
rect 4837 1392 4990 1402
rect 4998 1392 5028 1402
rect 5032 1392 5062 1406
rect 5090 1392 5103 1430
rect 5175 1436 5210 1444
rect 5175 1410 5176 1436
rect 5183 1410 5210 1436
rect 5118 1392 5148 1406
rect 5175 1402 5210 1410
rect 5212 1436 5253 1444
rect 5212 1410 5227 1436
rect 5234 1410 5253 1436
rect 5317 1432 5379 1444
rect 5391 1432 5466 1444
rect 5524 1432 5599 1444
rect 5611 1432 5642 1444
rect 5648 1432 5683 1444
rect 5317 1430 5479 1432
rect 5212 1402 5253 1410
rect 5335 1406 5348 1430
rect 5363 1428 5378 1430
rect 5412 1412 5479 1430
rect 5511 1430 5683 1432
rect 5511 1412 5591 1430
rect 5612 1428 5627 1430
rect 5175 1392 5176 1402
rect 5191 1392 5204 1402
rect 5218 1392 5219 1402
rect 5234 1392 5247 1402
rect 5262 1392 5292 1406
rect 5335 1392 5378 1406
rect 5402 1403 5409 1410
rect 5412 1402 5591 1412
rect 5385 1392 5415 1402
rect 5417 1392 5570 1402
rect 5578 1392 5608 1402
rect 5612 1392 5642 1406
rect 5670 1392 5683 1430
rect 5755 1436 5790 1444
rect 5755 1410 5756 1436
rect 5763 1410 5790 1436
rect 5698 1392 5728 1406
rect 5755 1402 5790 1410
rect 5792 1436 5833 1444
rect 5792 1410 5807 1436
rect 5814 1410 5833 1436
rect 5897 1432 5959 1444
rect 5971 1432 6046 1444
rect 6104 1432 6179 1444
rect 6191 1432 6222 1444
rect 6228 1432 6263 1444
rect 5897 1430 6059 1432
rect 5792 1402 5833 1410
rect 5915 1406 5928 1430
rect 5943 1428 5958 1430
rect 5992 1412 6059 1430
rect 6091 1430 6263 1432
rect 6091 1412 6171 1430
rect 6192 1428 6207 1430
rect 5755 1392 5756 1402
rect 5771 1392 5784 1402
rect 5798 1392 5799 1402
rect 5814 1392 5827 1402
rect 5842 1392 5872 1406
rect 5915 1392 5958 1406
rect 5982 1403 5989 1410
rect 5992 1402 6171 1412
rect 5965 1392 5995 1402
rect 5997 1392 6150 1402
rect 6158 1392 6188 1402
rect 6192 1392 6222 1406
rect 6250 1392 6263 1430
rect 6335 1436 6370 1444
rect 6335 1410 6336 1436
rect 6343 1410 6370 1436
rect 6278 1392 6308 1406
rect 6335 1402 6370 1410
rect 6372 1436 6413 1444
rect 6372 1410 6387 1436
rect 6394 1410 6413 1436
rect 6477 1432 6539 1444
rect 6551 1432 6626 1444
rect 6684 1432 6759 1444
rect 6771 1432 6802 1444
rect 6808 1432 6843 1444
rect 6477 1430 6639 1432
rect 6372 1402 6413 1410
rect 6495 1406 6508 1430
rect 6523 1428 6538 1430
rect 6572 1412 6639 1430
rect 6671 1430 6843 1432
rect 6671 1412 6751 1430
rect 6772 1428 6787 1430
rect 6335 1392 6336 1402
rect 6351 1392 6364 1402
rect 6378 1392 6379 1402
rect 6394 1392 6407 1402
rect 6422 1392 6452 1406
rect 6495 1392 6538 1406
rect 6562 1403 6569 1410
rect 6572 1402 6751 1412
rect 6545 1392 6575 1402
rect 6577 1392 6730 1402
rect 6738 1392 6768 1402
rect 6772 1392 6802 1406
rect 6830 1392 6843 1430
rect 6915 1436 6950 1444
rect 6915 1410 6916 1436
rect 6923 1410 6950 1436
rect 6858 1392 6888 1406
rect 6915 1402 6950 1410
rect 6915 1392 6916 1402
rect 6931 1392 6944 1402
rect 0 1378 6944 1392
rect 14 1348 27 1378
rect 42 1360 72 1378
rect 115 1364 129 1378
rect 165 1364 385 1378
rect 116 1362 129 1364
rect 82 1350 97 1362
rect 79 1348 101 1350
rect 106 1348 136 1362
rect 197 1360 350 1364
rect 179 1348 371 1360
rect 414 1348 444 1362
rect 450 1348 463 1378
rect 478 1360 508 1378
rect 551 1348 564 1378
rect 594 1348 607 1378
rect 622 1360 652 1378
rect 695 1364 709 1378
rect 745 1364 965 1378
rect 696 1362 709 1364
rect 662 1350 677 1362
rect 659 1348 681 1350
rect 686 1348 716 1362
rect 777 1360 930 1364
rect 759 1348 951 1360
rect 994 1348 1024 1362
rect 1030 1348 1043 1378
rect 1058 1360 1088 1378
rect 1131 1348 1144 1378
rect 1174 1348 1187 1378
rect 1202 1360 1232 1378
rect 1275 1364 1289 1378
rect 1325 1364 1545 1378
rect 1276 1362 1289 1364
rect 1242 1350 1257 1362
rect 1239 1348 1261 1350
rect 1266 1348 1296 1362
rect 1357 1360 1510 1364
rect 1339 1348 1531 1360
rect 1574 1348 1604 1362
rect 1610 1348 1623 1378
rect 1638 1360 1668 1378
rect 1711 1348 1724 1378
rect 1754 1348 1767 1378
rect 1782 1360 1812 1378
rect 1855 1364 1869 1378
rect 1905 1364 2125 1378
rect 1856 1362 1869 1364
rect 1822 1350 1837 1362
rect 1819 1348 1841 1350
rect 1846 1348 1876 1362
rect 1937 1360 2090 1364
rect 1919 1348 2111 1360
rect 2154 1348 2184 1362
rect 2190 1348 2203 1378
rect 2218 1360 2248 1378
rect 2291 1348 2304 1378
rect 2334 1348 2347 1378
rect 2362 1360 2392 1378
rect 2435 1364 2449 1378
rect 2485 1364 2705 1378
rect 2436 1362 2449 1364
rect 2402 1350 2417 1362
rect 2399 1348 2421 1350
rect 2426 1348 2456 1362
rect 2517 1360 2670 1364
rect 2499 1348 2691 1360
rect 2734 1348 2764 1362
rect 2770 1348 2783 1378
rect 2798 1360 2828 1378
rect 2871 1348 2884 1378
rect 2914 1348 2927 1378
rect 2942 1360 2972 1378
rect 3015 1364 3029 1378
rect 3065 1364 3285 1378
rect 3016 1362 3029 1364
rect 2982 1350 2997 1362
rect 2979 1348 3001 1350
rect 3006 1348 3036 1362
rect 3097 1360 3250 1364
rect 3079 1348 3271 1360
rect 3314 1348 3344 1362
rect 3350 1348 3363 1378
rect 3378 1360 3408 1378
rect 3451 1348 3464 1378
rect 3494 1348 3507 1378
rect 3522 1360 3552 1378
rect 3595 1364 3609 1378
rect 3645 1364 3865 1378
rect 3596 1362 3609 1364
rect 3562 1350 3577 1362
rect 3559 1348 3581 1350
rect 3586 1348 3616 1362
rect 3677 1360 3830 1364
rect 3659 1348 3851 1360
rect 3894 1348 3924 1362
rect 3930 1348 3943 1378
rect 3958 1360 3988 1378
rect 4031 1348 4044 1378
rect 4074 1348 4087 1378
rect 4102 1360 4132 1378
rect 4175 1364 4189 1378
rect 4225 1364 4445 1378
rect 4176 1362 4189 1364
rect 4142 1350 4157 1362
rect 4139 1348 4161 1350
rect 4166 1348 4196 1362
rect 4257 1360 4410 1364
rect 4239 1348 4431 1360
rect 4474 1348 4504 1362
rect 4510 1348 4523 1378
rect 4538 1360 4568 1378
rect 4611 1348 4624 1378
rect 4654 1348 4667 1378
rect 4682 1360 4712 1378
rect 4755 1364 4769 1378
rect 4805 1364 5025 1378
rect 4756 1362 4769 1364
rect 4722 1350 4737 1362
rect 4719 1348 4741 1350
rect 4746 1348 4776 1362
rect 4837 1360 4990 1364
rect 4819 1348 5011 1360
rect 5054 1348 5084 1362
rect 5090 1348 5103 1378
rect 5118 1360 5148 1378
rect 5191 1348 5204 1378
rect 5234 1348 5247 1378
rect 5262 1360 5292 1378
rect 5335 1364 5349 1378
rect 5385 1364 5605 1378
rect 5336 1362 5349 1364
rect 5302 1350 5317 1362
rect 5299 1348 5321 1350
rect 5326 1348 5356 1362
rect 5417 1360 5570 1364
rect 5399 1348 5591 1360
rect 5634 1348 5664 1362
rect 5670 1348 5683 1378
rect 5698 1360 5728 1378
rect 5771 1348 5784 1378
rect 5814 1348 5827 1378
rect 5842 1360 5872 1378
rect 5915 1364 5929 1378
rect 5965 1364 6185 1378
rect 5916 1362 5929 1364
rect 5882 1350 5897 1362
rect 5879 1348 5901 1350
rect 5906 1348 5936 1362
rect 5997 1360 6150 1364
rect 5979 1348 6171 1360
rect 6214 1348 6244 1362
rect 6250 1348 6263 1378
rect 6278 1360 6308 1378
rect 6351 1348 6364 1378
rect 6394 1348 6407 1378
rect 6422 1360 6452 1378
rect 6495 1364 6509 1378
rect 6545 1364 6765 1378
rect 6496 1362 6509 1364
rect 6462 1350 6477 1362
rect 6459 1348 6481 1350
rect 6486 1348 6516 1362
rect 6577 1360 6730 1364
rect 6559 1348 6751 1360
rect 6794 1348 6824 1362
rect 6830 1348 6843 1378
rect 6858 1360 6888 1378
rect 6931 1348 6944 1378
rect 0 1334 6944 1348
rect 14 1230 27 1334
rect 72 1312 73 1322
rect 88 1312 101 1322
rect 72 1308 101 1312
rect 106 1308 136 1334
rect 154 1320 170 1322
rect 242 1320 295 1334
rect 243 1318 307 1320
rect 350 1318 365 1334
rect 414 1331 444 1334
rect 414 1328 450 1331
rect 380 1320 396 1322
rect 154 1308 169 1312
rect 72 1306 169 1308
rect 197 1306 365 1318
rect 381 1308 396 1312
rect 414 1309 453 1328
rect 472 1322 479 1323
rect 478 1315 479 1322
rect 462 1312 463 1315
rect 478 1312 491 1315
rect 414 1308 444 1309
rect 453 1308 459 1309
rect 462 1308 491 1312
rect 381 1307 491 1308
rect 381 1306 497 1307
rect 56 1298 107 1306
rect 56 1286 81 1298
rect 88 1286 107 1298
rect 138 1298 188 1306
rect 138 1290 154 1298
rect 161 1296 188 1298
rect 197 1296 418 1306
rect 161 1286 418 1296
rect 447 1298 497 1306
rect 447 1289 463 1298
rect 56 1278 107 1286
rect 154 1278 418 1286
rect 444 1286 463 1289
rect 470 1286 497 1298
rect 444 1278 497 1286
rect 72 1270 73 1278
rect 88 1270 101 1278
rect 72 1262 88 1270
rect 69 1255 88 1258
rect 69 1246 91 1255
rect 42 1236 91 1246
rect 42 1230 72 1236
rect 91 1231 96 1236
rect 14 1214 88 1230
rect 106 1222 136 1278
rect 171 1268 379 1278
rect 414 1274 459 1278
rect 462 1277 463 1278
rect 478 1277 491 1278
rect 197 1238 386 1268
rect 212 1235 386 1238
rect 205 1232 386 1235
rect 14 1212 27 1214
rect 42 1212 76 1214
rect 14 1196 88 1212
rect 115 1208 128 1222
rect 143 1208 159 1224
rect 205 1219 216 1232
rect -2 1174 -1 1190
rect 14 1174 27 1196
rect 42 1174 72 1196
rect 115 1192 177 1208
rect 205 1201 216 1217
rect 221 1212 231 1232
rect 241 1212 255 1232
rect 258 1219 267 1232
rect 283 1219 292 1232
rect 221 1201 255 1212
rect 258 1201 267 1217
rect 283 1201 292 1217
rect 299 1212 309 1232
rect 319 1212 333 1232
rect 334 1219 345 1232
rect 299 1201 333 1212
rect 334 1201 345 1217
rect 391 1208 407 1224
rect 414 1222 444 1274
rect 478 1270 479 1277
rect 463 1262 479 1270
rect 450 1230 463 1249
rect 478 1230 508 1246
rect 450 1214 524 1230
rect 450 1212 463 1214
rect 478 1212 512 1214
rect 115 1190 128 1192
rect 143 1190 177 1192
rect 115 1174 177 1190
rect 221 1185 237 1188
rect 299 1185 329 1196
rect 377 1192 423 1208
rect 450 1196 524 1212
rect 377 1190 411 1192
rect 376 1174 423 1190
rect 450 1174 463 1196
rect 478 1174 508 1196
rect 535 1174 536 1190
rect 551 1174 564 1334
rect 594 1230 607 1334
rect 652 1312 653 1322
rect 668 1312 681 1322
rect 652 1308 681 1312
rect 686 1308 716 1334
rect 734 1320 750 1322
rect 822 1320 875 1334
rect 823 1318 887 1320
rect 930 1318 945 1334
rect 994 1331 1024 1334
rect 994 1328 1030 1331
rect 960 1320 976 1322
rect 734 1308 749 1312
rect 652 1306 749 1308
rect 777 1306 945 1318
rect 961 1308 976 1312
rect 994 1309 1033 1328
rect 1052 1322 1059 1323
rect 1058 1315 1059 1322
rect 1042 1312 1043 1315
rect 1058 1312 1071 1315
rect 994 1308 1024 1309
rect 1033 1308 1039 1309
rect 1042 1308 1071 1312
rect 961 1307 1071 1308
rect 961 1306 1077 1307
rect 636 1298 687 1306
rect 636 1286 661 1298
rect 668 1286 687 1298
rect 718 1298 768 1306
rect 718 1290 734 1298
rect 741 1296 768 1298
rect 777 1296 998 1306
rect 741 1286 998 1296
rect 1027 1298 1077 1306
rect 1027 1289 1043 1298
rect 636 1278 687 1286
rect 734 1278 998 1286
rect 1024 1286 1043 1289
rect 1050 1286 1077 1298
rect 1024 1278 1077 1286
rect 652 1270 653 1278
rect 668 1270 681 1278
rect 652 1262 668 1270
rect 649 1255 668 1258
rect 649 1246 671 1255
rect 622 1236 671 1246
rect 622 1230 652 1236
rect 671 1231 676 1236
rect 594 1214 668 1230
rect 686 1222 716 1278
rect 751 1268 959 1278
rect 994 1274 1039 1278
rect 1042 1277 1043 1278
rect 1058 1277 1071 1278
rect 777 1238 966 1268
rect 792 1235 966 1238
rect 785 1232 966 1235
rect 594 1212 607 1214
rect 622 1212 656 1214
rect 594 1196 668 1212
rect 695 1208 708 1222
rect 723 1208 739 1224
rect 785 1219 796 1232
rect 578 1174 579 1190
rect 594 1174 607 1196
rect 622 1174 652 1196
rect 695 1192 757 1208
rect 785 1201 796 1217
rect 801 1212 811 1232
rect 821 1212 835 1232
rect 838 1219 847 1232
rect 863 1219 872 1232
rect 801 1201 835 1212
rect 838 1201 847 1217
rect 863 1201 872 1217
rect 879 1212 889 1232
rect 899 1212 913 1232
rect 914 1219 925 1232
rect 879 1201 913 1212
rect 914 1201 925 1217
rect 971 1208 987 1224
rect 994 1222 1024 1274
rect 1058 1270 1059 1277
rect 1043 1262 1059 1270
rect 1030 1230 1043 1249
rect 1058 1230 1088 1246
rect 1030 1214 1104 1230
rect 1030 1212 1043 1214
rect 1058 1212 1092 1214
rect 695 1190 708 1192
rect 723 1190 757 1192
rect 695 1174 757 1190
rect 801 1185 817 1188
rect 879 1185 909 1196
rect 957 1192 1003 1208
rect 1030 1196 1104 1212
rect 957 1190 991 1192
rect 956 1174 1003 1190
rect 1030 1174 1043 1196
rect 1058 1174 1088 1196
rect 1115 1174 1116 1190
rect 1131 1174 1144 1334
rect 1174 1230 1187 1334
rect 1232 1312 1233 1322
rect 1248 1312 1261 1322
rect 1232 1308 1261 1312
rect 1266 1308 1296 1334
rect 1314 1320 1330 1322
rect 1402 1320 1455 1334
rect 1403 1318 1467 1320
rect 1510 1318 1525 1334
rect 1574 1331 1604 1334
rect 1574 1328 1610 1331
rect 1540 1320 1556 1322
rect 1314 1308 1329 1312
rect 1232 1306 1329 1308
rect 1357 1306 1525 1318
rect 1541 1308 1556 1312
rect 1574 1309 1613 1328
rect 1632 1322 1639 1323
rect 1638 1315 1639 1322
rect 1622 1312 1623 1315
rect 1638 1312 1651 1315
rect 1574 1308 1604 1309
rect 1613 1308 1619 1309
rect 1622 1308 1651 1312
rect 1541 1307 1651 1308
rect 1541 1306 1657 1307
rect 1216 1298 1267 1306
rect 1216 1286 1241 1298
rect 1248 1286 1267 1298
rect 1298 1298 1348 1306
rect 1298 1290 1314 1298
rect 1321 1296 1348 1298
rect 1357 1296 1578 1306
rect 1321 1286 1578 1296
rect 1607 1298 1657 1306
rect 1607 1289 1623 1298
rect 1216 1278 1267 1286
rect 1314 1278 1578 1286
rect 1604 1286 1623 1289
rect 1630 1286 1657 1298
rect 1604 1278 1657 1286
rect 1232 1270 1233 1278
rect 1248 1270 1261 1278
rect 1232 1262 1248 1270
rect 1229 1255 1248 1258
rect 1229 1246 1251 1255
rect 1202 1236 1251 1246
rect 1202 1230 1232 1236
rect 1251 1231 1256 1236
rect 1174 1214 1248 1230
rect 1266 1222 1296 1278
rect 1331 1268 1539 1278
rect 1574 1274 1619 1278
rect 1622 1277 1623 1278
rect 1638 1277 1651 1278
rect 1357 1238 1546 1268
rect 1372 1235 1546 1238
rect 1365 1232 1546 1235
rect 1174 1212 1187 1214
rect 1202 1212 1236 1214
rect 1174 1196 1248 1212
rect 1275 1208 1288 1222
rect 1303 1208 1319 1224
rect 1365 1219 1376 1232
rect 1158 1174 1159 1190
rect 1174 1174 1187 1196
rect 1202 1174 1232 1196
rect 1275 1192 1337 1208
rect 1365 1201 1376 1217
rect 1381 1212 1391 1232
rect 1401 1212 1415 1232
rect 1418 1219 1427 1232
rect 1443 1219 1452 1232
rect 1381 1201 1415 1212
rect 1418 1201 1427 1217
rect 1443 1201 1452 1217
rect 1459 1212 1469 1232
rect 1479 1212 1493 1232
rect 1494 1219 1505 1232
rect 1459 1201 1493 1212
rect 1494 1201 1505 1217
rect 1551 1208 1567 1224
rect 1574 1222 1604 1274
rect 1638 1270 1639 1277
rect 1623 1262 1639 1270
rect 1610 1230 1623 1249
rect 1638 1230 1668 1246
rect 1610 1214 1684 1230
rect 1610 1212 1623 1214
rect 1638 1212 1672 1214
rect 1275 1190 1288 1192
rect 1303 1190 1337 1192
rect 1275 1174 1337 1190
rect 1381 1185 1397 1188
rect 1459 1185 1489 1196
rect 1537 1192 1583 1208
rect 1610 1196 1684 1212
rect 1537 1190 1571 1192
rect 1536 1174 1583 1190
rect 1610 1174 1623 1196
rect 1638 1174 1668 1196
rect 1695 1174 1696 1190
rect 1711 1174 1724 1334
rect 1754 1230 1767 1334
rect 1812 1312 1813 1322
rect 1828 1312 1841 1322
rect 1812 1308 1841 1312
rect 1846 1308 1876 1334
rect 1894 1320 1910 1322
rect 1982 1320 2035 1334
rect 1983 1318 2047 1320
rect 2090 1318 2105 1334
rect 2154 1331 2184 1334
rect 2154 1328 2190 1331
rect 2120 1320 2136 1322
rect 1894 1308 1909 1312
rect 1812 1306 1909 1308
rect 1937 1306 2105 1318
rect 2121 1308 2136 1312
rect 2154 1309 2193 1328
rect 2212 1322 2219 1323
rect 2218 1315 2219 1322
rect 2202 1312 2203 1315
rect 2218 1312 2231 1315
rect 2154 1308 2184 1309
rect 2193 1308 2199 1309
rect 2202 1308 2231 1312
rect 2121 1307 2231 1308
rect 2121 1306 2237 1307
rect 1796 1298 1847 1306
rect 1796 1286 1821 1298
rect 1828 1286 1847 1298
rect 1878 1298 1928 1306
rect 1878 1290 1894 1298
rect 1901 1296 1928 1298
rect 1937 1296 2158 1306
rect 1901 1286 2158 1296
rect 2187 1298 2237 1306
rect 2187 1289 2203 1298
rect 1796 1278 1847 1286
rect 1894 1278 2158 1286
rect 2184 1286 2203 1289
rect 2210 1286 2237 1298
rect 2184 1278 2237 1286
rect 1812 1270 1813 1278
rect 1828 1270 1841 1278
rect 1812 1262 1828 1270
rect 1809 1255 1828 1258
rect 1809 1246 1831 1255
rect 1782 1236 1831 1246
rect 1782 1230 1812 1236
rect 1831 1231 1836 1236
rect 1754 1214 1828 1230
rect 1846 1222 1876 1278
rect 1911 1268 2119 1278
rect 2154 1274 2199 1278
rect 2202 1277 2203 1278
rect 2218 1277 2231 1278
rect 1937 1238 2126 1268
rect 1952 1235 2126 1238
rect 1945 1232 2126 1235
rect 1754 1212 1767 1214
rect 1782 1212 1816 1214
rect 1754 1196 1828 1212
rect 1855 1208 1868 1222
rect 1883 1208 1899 1224
rect 1945 1219 1956 1232
rect 1738 1174 1739 1190
rect 1754 1174 1767 1196
rect 1782 1174 1812 1196
rect 1855 1192 1917 1208
rect 1945 1201 1956 1217
rect 1961 1212 1971 1232
rect 1981 1212 1995 1232
rect 1998 1219 2007 1232
rect 2023 1219 2032 1232
rect 1961 1201 1995 1212
rect 1998 1201 2007 1217
rect 2023 1201 2032 1217
rect 2039 1212 2049 1232
rect 2059 1212 2073 1232
rect 2074 1219 2085 1232
rect 2039 1201 2073 1212
rect 2074 1201 2085 1217
rect 2131 1208 2147 1224
rect 2154 1222 2184 1274
rect 2218 1270 2219 1277
rect 2203 1262 2219 1270
rect 2190 1230 2203 1249
rect 2218 1230 2248 1246
rect 2190 1214 2264 1230
rect 2190 1212 2203 1214
rect 2218 1212 2252 1214
rect 1855 1190 1868 1192
rect 1883 1190 1917 1192
rect 1855 1174 1917 1190
rect 1961 1185 1977 1188
rect 2039 1185 2069 1196
rect 2117 1192 2163 1208
rect 2190 1196 2264 1212
rect 2117 1190 2151 1192
rect 2116 1174 2163 1190
rect 2190 1174 2203 1196
rect 2218 1174 2248 1196
rect 2275 1174 2276 1190
rect 2291 1174 2304 1334
rect 2334 1230 2347 1334
rect 2392 1312 2393 1322
rect 2408 1312 2421 1322
rect 2392 1308 2421 1312
rect 2426 1308 2456 1334
rect 2474 1320 2490 1322
rect 2562 1320 2615 1334
rect 2563 1318 2627 1320
rect 2670 1318 2685 1334
rect 2734 1331 2764 1334
rect 2734 1328 2770 1331
rect 2700 1320 2716 1322
rect 2474 1308 2489 1312
rect 2392 1306 2489 1308
rect 2517 1306 2685 1318
rect 2701 1308 2716 1312
rect 2734 1309 2773 1328
rect 2792 1322 2799 1323
rect 2798 1315 2799 1322
rect 2782 1312 2783 1315
rect 2798 1312 2811 1315
rect 2734 1308 2764 1309
rect 2773 1308 2779 1309
rect 2782 1308 2811 1312
rect 2701 1307 2811 1308
rect 2701 1306 2817 1307
rect 2376 1298 2427 1306
rect 2376 1286 2401 1298
rect 2408 1286 2427 1298
rect 2458 1298 2508 1306
rect 2458 1290 2474 1298
rect 2481 1296 2508 1298
rect 2517 1296 2738 1306
rect 2481 1286 2738 1296
rect 2767 1298 2817 1306
rect 2767 1289 2783 1298
rect 2376 1278 2427 1286
rect 2474 1278 2738 1286
rect 2764 1286 2783 1289
rect 2790 1286 2817 1298
rect 2764 1278 2817 1286
rect 2392 1270 2393 1278
rect 2408 1270 2421 1278
rect 2392 1262 2408 1270
rect 2389 1255 2408 1258
rect 2389 1246 2411 1255
rect 2362 1236 2411 1246
rect 2362 1230 2392 1236
rect 2411 1231 2416 1236
rect 2334 1214 2408 1230
rect 2426 1222 2456 1278
rect 2491 1268 2699 1278
rect 2734 1274 2779 1278
rect 2782 1277 2783 1278
rect 2798 1277 2811 1278
rect 2517 1238 2706 1268
rect 2532 1235 2706 1238
rect 2525 1232 2706 1235
rect 2334 1212 2347 1214
rect 2362 1212 2396 1214
rect 2334 1196 2408 1212
rect 2435 1208 2448 1222
rect 2463 1208 2479 1224
rect 2525 1219 2536 1232
rect 2318 1174 2319 1190
rect 2334 1174 2347 1196
rect 2362 1174 2392 1196
rect 2435 1192 2497 1208
rect 2525 1201 2536 1217
rect 2541 1212 2551 1232
rect 2561 1212 2575 1232
rect 2578 1219 2587 1232
rect 2603 1219 2612 1232
rect 2541 1201 2575 1212
rect 2578 1201 2587 1217
rect 2603 1201 2612 1217
rect 2619 1212 2629 1232
rect 2639 1212 2653 1232
rect 2654 1219 2665 1232
rect 2619 1201 2653 1212
rect 2654 1201 2665 1217
rect 2711 1208 2727 1224
rect 2734 1222 2764 1274
rect 2798 1270 2799 1277
rect 2783 1262 2799 1270
rect 2770 1230 2783 1249
rect 2798 1230 2828 1246
rect 2770 1214 2844 1230
rect 2770 1212 2783 1214
rect 2798 1212 2832 1214
rect 2435 1190 2448 1192
rect 2463 1190 2497 1192
rect 2435 1174 2497 1190
rect 2541 1185 2557 1188
rect 2619 1185 2649 1196
rect 2697 1192 2743 1208
rect 2770 1196 2844 1212
rect 2697 1190 2731 1192
rect 2696 1174 2743 1190
rect 2770 1174 2783 1196
rect 2798 1174 2828 1196
rect 2855 1174 2856 1190
rect 2871 1174 2884 1334
rect 2914 1230 2927 1334
rect 2972 1312 2973 1322
rect 2988 1312 3001 1322
rect 2972 1308 3001 1312
rect 3006 1308 3036 1334
rect 3054 1320 3070 1322
rect 3142 1320 3195 1334
rect 3143 1318 3205 1320
rect 3250 1318 3265 1334
rect 3314 1331 3344 1334
rect 3314 1328 3350 1331
rect 3280 1320 3296 1322
rect 3054 1308 3069 1312
rect 2972 1306 3069 1308
rect 3097 1306 3265 1318
rect 3281 1308 3296 1312
rect 3314 1309 3353 1328
rect 3372 1322 3379 1323
rect 3378 1315 3379 1322
rect 3362 1312 3363 1315
rect 3378 1312 3391 1315
rect 3314 1308 3344 1309
rect 3353 1308 3359 1309
rect 3362 1308 3391 1312
rect 3281 1307 3391 1308
rect 3281 1306 3397 1307
rect 2956 1298 3007 1306
rect 2956 1286 2981 1298
rect 2988 1286 3007 1298
rect 3038 1298 3088 1306
rect 3038 1290 3054 1298
rect 3061 1296 3088 1298
rect 3097 1296 3318 1306
rect 3061 1286 3318 1296
rect 3347 1298 3397 1306
rect 3347 1289 3363 1298
rect 2956 1278 3007 1286
rect 3054 1278 3318 1286
rect 3344 1286 3363 1289
rect 3370 1286 3397 1298
rect 3344 1278 3397 1286
rect 2972 1270 2973 1278
rect 2988 1270 3001 1278
rect 2972 1262 2988 1270
rect 2969 1255 2988 1258
rect 2969 1246 2991 1255
rect 2942 1236 2991 1246
rect 2942 1230 2972 1236
rect 2991 1231 2996 1236
rect 2914 1214 2988 1230
rect 3006 1222 3036 1278
rect 3071 1268 3279 1278
rect 3314 1274 3359 1278
rect 3362 1277 3363 1278
rect 3378 1277 3391 1278
rect 3097 1238 3286 1268
rect 3112 1235 3286 1238
rect 3105 1232 3286 1235
rect 2914 1212 2927 1214
rect 2942 1212 2976 1214
rect 2914 1196 2988 1212
rect 3015 1208 3028 1222
rect 3043 1208 3059 1224
rect 3105 1219 3116 1232
rect 2898 1174 2899 1190
rect 2914 1174 2927 1196
rect 2942 1174 2972 1196
rect 3015 1192 3077 1208
rect 3105 1201 3116 1217
rect 3121 1212 3131 1232
rect 3141 1212 3155 1232
rect 3158 1219 3167 1232
rect 3183 1219 3192 1232
rect 3121 1201 3155 1212
rect 3158 1201 3167 1217
rect 3183 1201 3192 1217
rect 3199 1212 3209 1232
rect 3219 1212 3233 1232
rect 3234 1219 3245 1232
rect 3199 1201 3233 1212
rect 3234 1201 3245 1217
rect 3291 1208 3307 1224
rect 3314 1222 3344 1274
rect 3378 1270 3379 1277
rect 3363 1262 3379 1270
rect 3350 1230 3363 1249
rect 3378 1230 3408 1246
rect 3350 1214 3424 1230
rect 3350 1212 3363 1214
rect 3378 1212 3412 1214
rect 3015 1190 3028 1192
rect 3043 1190 3077 1192
rect 3015 1174 3077 1190
rect 3121 1185 3137 1188
rect 3199 1185 3229 1196
rect 3277 1192 3323 1208
rect 3350 1196 3424 1212
rect 3277 1190 3311 1192
rect 3276 1174 3323 1190
rect 3350 1174 3363 1196
rect 3378 1174 3408 1196
rect 3435 1174 3436 1190
rect 3451 1174 3464 1334
rect 3494 1230 3507 1334
rect 3552 1312 3553 1322
rect 3568 1312 3581 1322
rect 3552 1308 3581 1312
rect 3586 1308 3616 1334
rect 3634 1320 3650 1322
rect 3722 1320 3775 1334
rect 3723 1318 3787 1320
rect 3830 1318 3845 1334
rect 3894 1331 3924 1334
rect 3894 1328 3930 1331
rect 3860 1320 3876 1322
rect 3634 1308 3649 1312
rect 3552 1306 3649 1308
rect 3677 1306 3845 1318
rect 3861 1308 3876 1312
rect 3894 1309 3933 1328
rect 3952 1322 3959 1323
rect 3958 1315 3959 1322
rect 3942 1312 3943 1315
rect 3958 1312 3971 1315
rect 3894 1308 3924 1309
rect 3933 1308 3939 1309
rect 3942 1308 3971 1312
rect 3861 1307 3971 1308
rect 3861 1306 3977 1307
rect 3536 1298 3587 1306
rect 3536 1286 3561 1298
rect 3568 1286 3587 1298
rect 3618 1298 3668 1306
rect 3618 1290 3634 1298
rect 3641 1296 3668 1298
rect 3677 1296 3898 1306
rect 3641 1286 3898 1296
rect 3927 1298 3977 1306
rect 3927 1289 3943 1298
rect 3536 1278 3587 1286
rect 3634 1278 3898 1286
rect 3924 1286 3943 1289
rect 3950 1286 3977 1298
rect 3924 1278 3977 1286
rect 3552 1270 3553 1278
rect 3568 1270 3581 1278
rect 3552 1262 3568 1270
rect 3549 1255 3568 1258
rect 3549 1246 3571 1255
rect 3522 1236 3571 1246
rect 3522 1230 3552 1236
rect 3571 1231 3576 1236
rect 3494 1214 3568 1230
rect 3586 1222 3616 1278
rect 3651 1268 3859 1278
rect 3894 1274 3939 1278
rect 3942 1277 3943 1278
rect 3958 1277 3971 1278
rect 3677 1238 3866 1268
rect 3692 1235 3866 1238
rect 3685 1232 3866 1235
rect 3494 1212 3507 1214
rect 3522 1212 3556 1214
rect 3494 1196 3568 1212
rect 3595 1208 3608 1222
rect 3623 1208 3639 1224
rect 3685 1219 3696 1232
rect 3478 1174 3479 1190
rect 3494 1174 3507 1196
rect 3522 1174 3552 1196
rect 3595 1192 3657 1208
rect 3685 1201 3696 1217
rect 3701 1212 3711 1232
rect 3721 1212 3735 1232
rect 3738 1219 3747 1232
rect 3763 1219 3772 1232
rect 3701 1201 3735 1212
rect 3738 1201 3747 1217
rect 3763 1201 3772 1217
rect 3779 1212 3789 1232
rect 3799 1212 3813 1232
rect 3814 1219 3825 1232
rect 3779 1201 3813 1212
rect 3814 1201 3825 1217
rect 3871 1208 3887 1224
rect 3894 1222 3924 1274
rect 3958 1270 3959 1277
rect 3943 1262 3959 1270
rect 3930 1230 3943 1249
rect 3958 1230 3988 1246
rect 3930 1214 4004 1230
rect 3930 1212 3943 1214
rect 3958 1212 3992 1214
rect 3595 1190 3608 1192
rect 3623 1190 3657 1192
rect 3595 1174 3657 1190
rect 3701 1185 3717 1188
rect 3779 1185 3809 1196
rect 3857 1192 3903 1208
rect 3930 1196 4004 1212
rect 3857 1190 3891 1192
rect 3856 1174 3903 1190
rect 3930 1174 3943 1196
rect 3958 1174 3988 1196
rect 4015 1174 4016 1190
rect 4031 1174 4044 1334
rect 4074 1230 4087 1334
rect 4132 1312 4133 1322
rect 4148 1312 4161 1322
rect 4132 1308 4161 1312
rect 4166 1308 4196 1334
rect 4214 1320 4230 1322
rect 4302 1320 4355 1334
rect 4303 1318 4367 1320
rect 4410 1318 4425 1334
rect 4474 1331 4504 1334
rect 4474 1328 4510 1331
rect 4440 1320 4456 1322
rect 4214 1308 4229 1312
rect 4132 1306 4229 1308
rect 4257 1306 4425 1318
rect 4441 1308 4456 1312
rect 4474 1309 4513 1328
rect 4532 1322 4539 1323
rect 4538 1315 4539 1322
rect 4522 1312 4523 1315
rect 4538 1312 4551 1315
rect 4474 1308 4504 1309
rect 4513 1308 4519 1309
rect 4522 1308 4551 1312
rect 4441 1307 4551 1308
rect 4441 1306 4557 1307
rect 4116 1298 4167 1306
rect 4116 1286 4141 1298
rect 4148 1286 4167 1298
rect 4198 1298 4248 1306
rect 4198 1290 4214 1298
rect 4221 1296 4248 1298
rect 4257 1296 4478 1306
rect 4221 1286 4478 1296
rect 4507 1298 4557 1306
rect 4507 1289 4523 1298
rect 4116 1278 4167 1286
rect 4214 1278 4478 1286
rect 4504 1286 4523 1289
rect 4530 1286 4557 1298
rect 4504 1278 4557 1286
rect 4132 1270 4133 1278
rect 4148 1270 4161 1278
rect 4132 1262 4148 1270
rect 4129 1255 4148 1258
rect 4129 1246 4151 1255
rect 4102 1236 4151 1246
rect 4102 1230 4132 1236
rect 4151 1231 4156 1236
rect 4074 1214 4148 1230
rect 4166 1222 4196 1278
rect 4231 1268 4439 1278
rect 4474 1274 4519 1278
rect 4522 1277 4523 1278
rect 4538 1277 4551 1278
rect 4257 1238 4446 1268
rect 4272 1235 4446 1238
rect 4265 1232 4446 1235
rect 4074 1212 4087 1214
rect 4102 1212 4136 1214
rect 4074 1196 4148 1212
rect 4175 1208 4188 1222
rect 4203 1208 4219 1224
rect 4265 1219 4276 1232
rect 4058 1174 4059 1190
rect 4074 1174 4087 1196
rect 4102 1174 4132 1196
rect 4175 1192 4237 1208
rect 4265 1201 4276 1217
rect 4281 1212 4291 1232
rect 4301 1212 4315 1232
rect 4318 1219 4327 1232
rect 4343 1219 4352 1232
rect 4281 1201 4315 1212
rect 4318 1201 4327 1217
rect 4343 1201 4352 1217
rect 4359 1212 4369 1232
rect 4379 1212 4393 1232
rect 4394 1219 4405 1232
rect 4359 1201 4393 1212
rect 4394 1201 4405 1217
rect 4451 1208 4467 1224
rect 4474 1222 4504 1274
rect 4538 1270 4539 1277
rect 4523 1262 4539 1270
rect 4510 1230 4523 1249
rect 4538 1230 4568 1246
rect 4510 1214 4584 1230
rect 4510 1212 4523 1214
rect 4538 1212 4572 1214
rect 4175 1190 4188 1192
rect 4203 1190 4237 1192
rect 4175 1174 4237 1190
rect 4281 1185 4297 1188
rect 4359 1185 4389 1196
rect 4437 1192 4483 1208
rect 4510 1196 4584 1212
rect 4437 1190 4471 1192
rect 4436 1174 4483 1190
rect 4510 1174 4523 1196
rect 4538 1174 4568 1196
rect 4595 1174 4596 1190
rect 4611 1174 4624 1334
rect 4654 1230 4667 1334
rect 4712 1312 4713 1322
rect 4733 1320 4741 1322
rect 4731 1318 4741 1320
rect 4728 1312 4741 1318
rect 4712 1308 4741 1312
rect 4746 1308 4776 1334
rect 4794 1320 4810 1322
rect 4882 1320 4933 1334
rect 4883 1318 4947 1320
rect 4899 1317 4931 1318
rect 4990 1317 5005 1334
rect 5054 1331 5084 1334
rect 5054 1328 5090 1331
rect 5020 1320 5036 1322
rect 4794 1308 4809 1312
rect 4712 1306 4809 1308
rect 4837 1306 5005 1317
rect 5021 1308 5036 1312
rect 5054 1309 5093 1328
rect 5112 1322 5119 1323
rect 5118 1315 5119 1322
rect 5102 1312 5103 1315
rect 5118 1312 5131 1315
rect 5054 1308 5084 1309
rect 5093 1308 5099 1309
rect 5102 1308 5131 1312
rect 5021 1307 5131 1308
rect 5021 1306 5137 1307
rect 4696 1298 4747 1306
rect 4696 1286 4721 1298
rect 4728 1286 4747 1298
rect 4778 1298 4828 1306
rect 4778 1290 4794 1298
rect 4801 1296 4828 1298
rect 4837 1296 5058 1306
rect 4801 1286 5058 1296
rect 5087 1298 5137 1306
rect 5087 1289 5103 1298
rect 4696 1278 4747 1286
rect 4794 1278 5058 1286
rect 5084 1286 5103 1289
rect 5110 1286 5137 1298
rect 5084 1278 5137 1286
rect 4712 1270 4713 1278
rect 4728 1270 4741 1278
rect 4712 1262 4728 1270
rect 4709 1255 4728 1258
rect 4709 1246 4731 1255
rect 4682 1236 4731 1246
rect 4682 1230 4712 1236
rect 4731 1231 4736 1236
rect 4654 1214 4728 1230
rect 4746 1222 4776 1278
rect 4811 1268 5019 1278
rect 5054 1274 5099 1278
rect 5102 1277 5103 1278
rect 5118 1277 5131 1278
rect 4837 1238 5026 1268
rect 4852 1235 5026 1238
rect 4845 1232 5026 1235
rect 4654 1212 4667 1214
rect 4682 1212 4716 1214
rect 4654 1196 4728 1212
rect 4755 1208 4768 1222
rect 4783 1208 4799 1224
rect 4845 1219 4856 1232
rect 4638 1174 4639 1190
rect 4654 1174 4667 1196
rect 4682 1174 4712 1196
rect 4755 1192 4817 1208
rect 4845 1201 4856 1217
rect 4861 1212 4871 1232
rect 4881 1212 4895 1232
rect 4898 1219 4907 1232
rect 4923 1219 4932 1232
rect 4861 1201 4895 1212
rect 4898 1201 4907 1217
rect 4923 1201 4932 1217
rect 4939 1212 4949 1232
rect 4959 1212 4973 1232
rect 4974 1219 4985 1232
rect 4939 1201 4973 1212
rect 4974 1201 4985 1217
rect 5031 1208 5047 1224
rect 5054 1222 5084 1274
rect 5118 1270 5119 1277
rect 5103 1262 5119 1270
rect 5090 1230 5103 1249
rect 5118 1230 5148 1246
rect 5090 1214 5164 1230
rect 5090 1212 5103 1214
rect 5118 1212 5152 1214
rect 4755 1190 4768 1192
rect 4783 1190 4817 1192
rect 4755 1174 4817 1190
rect 4861 1185 4877 1188
rect 4939 1185 4969 1196
rect 5017 1192 5063 1208
rect 5090 1196 5164 1212
rect 5017 1190 5051 1192
rect 5016 1174 5063 1190
rect 5090 1174 5103 1196
rect 5118 1174 5148 1196
rect 5175 1174 5176 1190
rect 5191 1174 5204 1334
rect 5234 1230 5247 1334
rect 5292 1312 5293 1322
rect 5313 1320 5321 1322
rect 5311 1318 5321 1320
rect 5308 1312 5321 1318
rect 5292 1308 5321 1312
rect 5326 1308 5356 1334
rect 5374 1320 5390 1322
rect 5462 1320 5513 1334
rect 5463 1318 5527 1320
rect 5479 1317 5511 1318
rect 5570 1317 5585 1334
rect 5634 1331 5664 1334
rect 5634 1328 5670 1331
rect 5600 1320 5616 1322
rect 5374 1308 5389 1312
rect 5292 1306 5389 1308
rect 5417 1306 5585 1317
rect 5601 1308 5616 1312
rect 5634 1309 5673 1328
rect 5692 1322 5699 1323
rect 5698 1315 5699 1322
rect 5682 1312 5683 1315
rect 5698 1312 5711 1315
rect 5634 1308 5664 1309
rect 5673 1308 5679 1309
rect 5682 1308 5711 1312
rect 5601 1307 5711 1308
rect 5601 1306 5717 1307
rect 5276 1298 5327 1306
rect 5276 1286 5301 1298
rect 5308 1286 5327 1298
rect 5358 1298 5408 1306
rect 5358 1290 5374 1298
rect 5381 1296 5408 1298
rect 5417 1296 5638 1306
rect 5381 1286 5638 1296
rect 5667 1298 5717 1306
rect 5667 1289 5683 1298
rect 5276 1278 5327 1286
rect 5374 1278 5638 1286
rect 5664 1286 5683 1289
rect 5690 1286 5717 1298
rect 5664 1278 5717 1286
rect 5292 1270 5293 1278
rect 5308 1270 5321 1278
rect 5292 1262 5308 1270
rect 5289 1255 5308 1258
rect 5289 1246 5311 1255
rect 5262 1236 5311 1246
rect 5262 1230 5292 1236
rect 5311 1231 5316 1236
rect 5234 1214 5308 1230
rect 5326 1222 5356 1278
rect 5391 1268 5599 1278
rect 5634 1274 5679 1278
rect 5682 1277 5683 1278
rect 5698 1277 5711 1278
rect 5417 1238 5606 1268
rect 5432 1235 5606 1238
rect 5425 1232 5606 1235
rect 5234 1212 5247 1214
rect 5262 1212 5296 1214
rect 5234 1196 5308 1212
rect 5335 1208 5348 1222
rect 5363 1208 5379 1224
rect 5425 1219 5436 1232
rect 5218 1174 5219 1190
rect 5234 1174 5247 1196
rect 5262 1174 5292 1196
rect 5335 1192 5397 1208
rect 5425 1201 5436 1217
rect 5441 1212 5451 1232
rect 5461 1212 5475 1232
rect 5478 1219 5487 1232
rect 5503 1219 5512 1232
rect 5441 1201 5475 1212
rect 5478 1201 5487 1217
rect 5503 1201 5512 1217
rect 5519 1212 5529 1232
rect 5539 1212 5553 1232
rect 5554 1219 5565 1232
rect 5519 1201 5553 1212
rect 5554 1201 5565 1217
rect 5611 1208 5627 1224
rect 5634 1222 5664 1274
rect 5698 1270 5699 1277
rect 5683 1262 5699 1270
rect 5670 1230 5683 1249
rect 5698 1230 5728 1246
rect 5670 1214 5744 1230
rect 5670 1212 5683 1214
rect 5698 1212 5732 1214
rect 5335 1190 5348 1192
rect 5363 1190 5397 1192
rect 5335 1174 5397 1190
rect 5441 1185 5457 1188
rect 5519 1185 5549 1196
rect 5597 1192 5643 1208
rect 5670 1196 5744 1212
rect 5597 1190 5631 1192
rect 5596 1174 5643 1190
rect 5670 1174 5683 1196
rect 5698 1174 5728 1196
rect 5755 1174 5756 1190
rect 5771 1174 5784 1334
rect 5814 1230 5827 1334
rect 5872 1312 5873 1322
rect 5893 1320 5901 1322
rect 5891 1318 5901 1320
rect 5888 1312 5901 1318
rect 5872 1308 5901 1312
rect 5906 1308 5936 1334
rect 5954 1320 5970 1322
rect 6042 1320 6093 1334
rect 6043 1318 6107 1320
rect 6059 1317 6091 1318
rect 6150 1317 6165 1334
rect 6214 1331 6244 1334
rect 6214 1328 6250 1331
rect 6180 1320 6196 1322
rect 5954 1308 5969 1312
rect 5872 1306 5969 1308
rect 5997 1306 6165 1317
rect 6181 1308 6196 1312
rect 6214 1309 6253 1328
rect 6272 1322 6279 1323
rect 6278 1315 6279 1322
rect 6262 1312 6263 1315
rect 6278 1312 6291 1315
rect 6214 1308 6244 1309
rect 6253 1308 6259 1309
rect 6262 1308 6291 1312
rect 6181 1307 6291 1308
rect 6181 1306 6297 1307
rect 5856 1298 5907 1306
rect 5856 1286 5881 1298
rect 5888 1286 5907 1298
rect 5938 1298 5988 1306
rect 5938 1290 5954 1298
rect 5961 1296 5988 1298
rect 5997 1296 6218 1306
rect 5961 1286 6218 1296
rect 6247 1298 6297 1306
rect 6247 1289 6263 1298
rect 5856 1278 5907 1286
rect 5954 1278 6218 1286
rect 6244 1286 6263 1289
rect 6270 1286 6297 1298
rect 6244 1278 6297 1286
rect 5872 1270 5873 1278
rect 5888 1270 5901 1278
rect 5872 1262 5888 1270
rect 5869 1255 5888 1258
rect 5869 1246 5891 1255
rect 5842 1236 5891 1246
rect 5842 1230 5872 1236
rect 5891 1231 5896 1236
rect 5814 1214 5888 1230
rect 5906 1222 5936 1278
rect 5971 1268 6179 1278
rect 6214 1274 6259 1278
rect 6262 1277 6263 1278
rect 6278 1277 6291 1278
rect 5997 1238 6186 1268
rect 6012 1235 6186 1238
rect 6005 1232 6186 1235
rect 5814 1212 5827 1214
rect 5842 1212 5876 1214
rect 5814 1196 5888 1212
rect 5915 1208 5928 1222
rect 5943 1208 5959 1224
rect 6005 1219 6016 1232
rect 5798 1174 5799 1190
rect 5814 1174 5827 1196
rect 5842 1174 5872 1196
rect 5915 1192 5977 1208
rect 6005 1201 6016 1217
rect 6021 1212 6031 1232
rect 6041 1212 6055 1232
rect 6058 1219 6067 1232
rect 6083 1219 6092 1232
rect 6021 1201 6055 1212
rect 6058 1201 6067 1217
rect 6083 1201 6092 1217
rect 6099 1212 6109 1232
rect 6119 1212 6133 1232
rect 6134 1219 6145 1232
rect 6099 1201 6133 1212
rect 6134 1201 6145 1217
rect 6191 1208 6207 1224
rect 6214 1222 6244 1274
rect 6278 1270 6279 1277
rect 6263 1262 6279 1270
rect 6250 1230 6263 1249
rect 6278 1230 6308 1246
rect 6250 1214 6324 1230
rect 6250 1212 6263 1214
rect 6278 1212 6312 1214
rect 5915 1190 5928 1192
rect 5943 1190 5977 1192
rect 5915 1174 5977 1190
rect 6021 1185 6037 1188
rect 6099 1185 6129 1196
rect 6177 1192 6223 1208
rect 6250 1196 6324 1212
rect 6177 1190 6211 1192
rect 6176 1174 6223 1190
rect 6250 1174 6263 1196
rect 6278 1174 6308 1196
rect 6335 1174 6336 1190
rect 6351 1174 6364 1334
rect 6394 1230 6407 1334
rect 6452 1312 6453 1322
rect 6473 1320 6481 1322
rect 6471 1318 6481 1320
rect 6468 1312 6481 1318
rect 6452 1308 6481 1312
rect 6486 1308 6516 1334
rect 6534 1320 6550 1322
rect 6622 1320 6673 1334
rect 6623 1318 6687 1320
rect 6639 1317 6671 1318
rect 6730 1317 6745 1334
rect 6794 1331 6824 1334
rect 6794 1328 6830 1331
rect 6760 1320 6776 1322
rect 6534 1308 6549 1312
rect 6452 1306 6549 1308
rect 6577 1306 6745 1317
rect 6761 1308 6776 1312
rect 6794 1309 6833 1328
rect 6852 1322 6859 1323
rect 6858 1315 6859 1322
rect 6842 1312 6843 1315
rect 6858 1312 6871 1315
rect 6794 1308 6824 1309
rect 6833 1308 6839 1309
rect 6842 1308 6871 1312
rect 6761 1307 6871 1308
rect 6761 1306 6877 1307
rect 6436 1298 6487 1306
rect 6436 1286 6461 1298
rect 6468 1286 6487 1298
rect 6518 1298 6568 1306
rect 6518 1290 6534 1298
rect 6541 1296 6568 1298
rect 6577 1296 6798 1306
rect 6541 1286 6798 1296
rect 6827 1298 6877 1306
rect 6827 1289 6843 1298
rect 6436 1278 6487 1286
rect 6534 1278 6798 1286
rect 6824 1286 6843 1289
rect 6850 1286 6877 1298
rect 6824 1278 6877 1286
rect 6452 1270 6453 1278
rect 6468 1270 6481 1278
rect 6452 1262 6468 1270
rect 6449 1255 6468 1258
rect 6449 1246 6471 1255
rect 6422 1236 6471 1246
rect 6422 1230 6452 1236
rect 6471 1231 6476 1236
rect 6394 1214 6468 1230
rect 6486 1222 6516 1278
rect 6551 1268 6759 1278
rect 6794 1274 6839 1278
rect 6842 1277 6843 1278
rect 6858 1277 6871 1278
rect 6577 1238 6766 1268
rect 6592 1235 6766 1238
rect 6585 1232 6766 1235
rect 6394 1212 6407 1214
rect 6422 1212 6456 1214
rect 6394 1196 6468 1212
rect 6495 1208 6508 1222
rect 6523 1208 6539 1224
rect 6585 1219 6596 1232
rect 6378 1174 6379 1190
rect 6394 1174 6407 1196
rect 6422 1174 6452 1196
rect 6495 1192 6557 1208
rect 6585 1201 6596 1217
rect 6601 1212 6611 1232
rect 6621 1212 6635 1232
rect 6638 1219 6647 1232
rect 6663 1219 6672 1232
rect 6601 1201 6635 1212
rect 6638 1201 6647 1217
rect 6663 1201 6672 1217
rect 6679 1212 6689 1232
rect 6699 1212 6713 1232
rect 6714 1219 6725 1232
rect 6679 1201 6713 1212
rect 6714 1201 6725 1217
rect 6771 1208 6787 1224
rect 6794 1222 6824 1274
rect 6858 1270 6859 1277
rect 6843 1262 6859 1270
rect 6830 1230 6843 1249
rect 6858 1230 6888 1246
rect 6830 1214 6904 1230
rect 6830 1212 6843 1214
rect 6858 1212 6892 1214
rect 6495 1190 6508 1192
rect 6523 1190 6557 1192
rect 6495 1174 6557 1190
rect 6601 1185 6617 1188
rect 6679 1185 6709 1196
rect 6757 1192 6803 1208
rect 6830 1196 6904 1212
rect 6757 1190 6791 1192
rect 6756 1174 6803 1190
rect 6830 1174 6843 1196
rect 6858 1174 6888 1196
rect 6915 1174 6916 1190
rect 6931 1174 6944 1334
rect -8 1166 33 1174
rect -8 1140 7 1166
rect 14 1140 33 1166
rect 97 1162 159 1174
rect 171 1162 246 1174
rect 304 1162 379 1174
rect 391 1162 422 1174
rect 428 1162 463 1174
rect 97 1160 259 1162
rect -8 1132 33 1140
rect 115 1136 128 1160
rect 143 1158 158 1160
rect -2 1122 -1 1132
rect 14 1122 27 1132
rect 42 1122 72 1136
rect 115 1122 158 1136
rect 182 1133 189 1140
rect 192 1136 259 1160
rect 291 1160 463 1162
rect 261 1138 289 1142
rect 291 1138 371 1160
rect 392 1158 407 1160
rect 261 1136 371 1138
rect 192 1132 371 1136
rect 165 1122 195 1132
rect 197 1122 350 1132
rect 358 1122 388 1132
rect 392 1122 422 1136
rect 450 1122 463 1160
rect 535 1166 570 1174
rect 535 1140 536 1166
rect 543 1140 570 1166
rect 478 1122 508 1136
rect 535 1132 570 1140
rect 572 1166 613 1174
rect 572 1140 587 1166
rect 594 1140 613 1166
rect 677 1162 739 1174
rect 751 1162 826 1174
rect 884 1162 959 1174
rect 971 1162 1002 1174
rect 1008 1162 1043 1174
rect 677 1160 839 1162
rect 572 1132 613 1140
rect 695 1136 708 1160
rect 723 1158 738 1160
rect 535 1122 536 1132
rect 551 1122 564 1132
rect 578 1122 579 1132
rect 594 1122 607 1132
rect 622 1122 652 1136
rect 695 1122 738 1136
rect 762 1133 769 1140
rect 772 1136 839 1160
rect 871 1160 1043 1162
rect 841 1138 869 1142
rect 871 1138 951 1160
rect 972 1158 987 1160
rect 841 1136 951 1138
rect 772 1132 951 1136
rect 745 1122 775 1132
rect 777 1122 930 1132
rect 938 1122 968 1132
rect 972 1122 1002 1136
rect 1030 1122 1043 1160
rect 1115 1166 1150 1174
rect 1115 1140 1116 1166
rect 1123 1140 1150 1166
rect 1058 1122 1088 1136
rect 1115 1132 1150 1140
rect 1152 1166 1193 1174
rect 1152 1140 1167 1166
rect 1174 1140 1193 1166
rect 1257 1162 1319 1174
rect 1331 1162 1406 1174
rect 1464 1162 1539 1174
rect 1551 1162 1582 1174
rect 1588 1162 1623 1174
rect 1257 1160 1419 1162
rect 1152 1132 1193 1140
rect 1275 1136 1288 1160
rect 1303 1158 1318 1160
rect 1115 1122 1116 1132
rect 1131 1122 1144 1132
rect 1158 1122 1159 1132
rect 1174 1122 1187 1132
rect 1202 1122 1232 1136
rect 1275 1122 1318 1136
rect 1342 1133 1349 1140
rect 1352 1136 1419 1160
rect 1451 1160 1623 1162
rect 1421 1138 1449 1142
rect 1451 1138 1531 1160
rect 1552 1158 1567 1160
rect 1421 1136 1531 1138
rect 1352 1132 1531 1136
rect 1325 1122 1355 1132
rect 1357 1122 1510 1132
rect 1518 1122 1548 1132
rect 1552 1122 1582 1136
rect 1610 1122 1623 1160
rect 1695 1166 1730 1174
rect 1695 1140 1696 1166
rect 1703 1140 1730 1166
rect 1638 1122 1668 1136
rect 1695 1132 1730 1140
rect 1732 1166 1773 1174
rect 1732 1140 1747 1166
rect 1754 1140 1773 1166
rect 1837 1162 1899 1174
rect 1911 1162 1986 1174
rect 2044 1162 2119 1174
rect 2131 1162 2162 1174
rect 2168 1162 2203 1174
rect 1837 1160 1999 1162
rect 1732 1132 1773 1140
rect 1855 1136 1868 1160
rect 1883 1158 1898 1160
rect 1695 1122 1696 1132
rect 1711 1122 1724 1132
rect 1738 1122 1739 1132
rect 1754 1122 1767 1132
rect 1782 1122 1812 1136
rect 1855 1122 1898 1136
rect 1922 1133 1929 1140
rect 1932 1136 1999 1160
rect 2031 1160 2203 1162
rect 2001 1138 2029 1142
rect 2031 1138 2111 1160
rect 2132 1158 2147 1160
rect 2001 1136 2111 1138
rect 1932 1132 2111 1136
rect 1905 1122 1935 1132
rect 1937 1122 2090 1132
rect 2098 1122 2128 1132
rect 2132 1122 2162 1136
rect 2190 1122 2203 1160
rect 2275 1166 2310 1174
rect 2275 1140 2276 1166
rect 2283 1140 2310 1166
rect 2218 1122 2248 1136
rect 2275 1132 2310 1140
rect 2312 1166 2353 1174
rect 2312 1140 2327 1166
rect 2334 1140 2353 1166
rect 2417 1162 2479 1174
rect 2491 1162 2566 1174
rect 2624 1162 2699 1174
rect 2711 1162 2742 1174
rect 2748 1162 2783 1174
rect 2417 1160 2579 1162
rect 2312 1132 2353 1140
rect 2435 1136 2448 1160
rect 2463 1158 2478 1160
rect 2275 1122 2276 1132
rect 2291 1122 2304 1132
rect 2318 1122 2319 1132
rect 2334 1122 2347 1132
rect 2362 1122 2392 1136
rect 2435 1122 2478 1136
rect 2502 1133 2509 1140
rect 2512 1136 2579 1160
rect 2611 1160 2783 1162
rect 2581 1138 2609 1142
rect 2611 1138 2691 1160
rect 2712 1158 2727 1160
rect 2581 1136 2691 1138
rect 2512 1132 2691 1136
rect 2485 1122 2515 1132
rect 2517 1122 2670 1132
rect 2678 1122 2708 1132
rect 2712 1122 2742 1136
rect 2770 1122 2783 1160
rect 2855 1166 2890 1174
rect 2855 1140 2856 1166
rect 2863 1140 2890 1166
rect 2798 1122 2828 1136
rect 2855 1132 2890 1140
rect 2892 1166 2933 1174
rect 2892 1140 2907 1166
rect 2914 1140 2933 1166
rect 2997 1162 3059 1174
rect 3071 1162 3146 1174
rect 3204 1162 3279 1174
rect 3291 1162 3322 1174
rect 3328 1162 3363 1174
rect 2997 1160 3159 1162
rect 2892 1132 2933 1140
rect 3015 1136 3028 1160
rect 3043 1158 3058 1160
rect 2855 1122 2856 1132
rect 2871 1122 2884 1132
rect 2898 1122 2899 1132
rect 2914 1122 2927 1132
rect 2942 1122 2972 1136
rect 3015 1122 3058 1136
rect 3082 1133 3089 1140
rect 3092 1136 3159 1160
rect 3191 1160 3363 1162
rect 3161 1138 3189 1142
rect 3191 1138 3271 1160
rect 3292 1158 3307 1160
rect 3161 1136 3271 1138
rect 3092 1132 3271 1136
rect 3065 1122 3095 1132
rect 3097 1122 3250 1132
rect 3258 1122 3288 1132
rect 3292 1122 3322 1136
rect 3350 1122 3363 1160
rect 3435 1166 3470 1174
rect 3435 1140 3436 1166
rect 3443 1140 3470 1166
rect 3378 1122 3408 1136
rect 3435 1132 3470 1140
rect 3472 1166 3513 1174
rect 3472 1140 3487 1166
rect 3494 1140 3513 1166
rect 3577 1162 3639 1174
rect 3651 1162 3726 1174
rect 3784 1162 3859 1174
rect 3871 1162 3902 1174
rect 3908 1162 3943 1174
rect 3577 1160 3739 1162
rect 3472 1132 3513 1140
rect 3595 1136 3608 1160
rect 3623 1158 3638 1160
rect 3435 1122 3436 1132
rect 3451 1122 3464 1132
rect 3478 1122 3479 1132
rect 3494 1122 3507 1132
rect 3522 1122 3552 1136
rect 3595 1122 3638 1136
rect 3662 1133 3669 1140
rect 3672 1136 3739 1160
rect 3771 1160 3943 1162
rect 3741 1138 3769 1142
rect 3771 1138 3851 1160
rect 3872 1158 3887 1160
rect 3741 1136 3851 1138
rect 3672 1132 3851 1136
rect 3645 1122 3675 1132
rect 3677 1122 3830 1132
rect 3838 1122 3868 1132
rect 3872 1122 3902 1136
rect 3930 1122 3943 1160
rect 4015 1166 4050 1174
rect 4015 1140 4016 1166
rect 4023 1140 4050 1166
rect 3958 1122 3988 1136
rect 4015 1132 4050 1140
rect 4052 1166 4093 1174
rect 4052 1140 4067 1166
rect 4074 1140 4093 1166
rect 4157 1162 4219 1174
rect 4231 1162 4306 1174
rect 4364 1162 4439 1174
rect 4451 1162 4482 1174
rect 4488 1162 4523 1174
rect 4157 1160 4319 1162
rect 4052 1132 4093 1140
rect 4175 1136 4188 1160
rect 4203 1158 4218 1160
rect 4015 1122 4016 1132
rect 4031 1122 4044 1132
rect 4058 1122 4059 1132
rect 4074 1122 4087 1132
rect 4102 1122 4132 1136
rect 4175 1122 4218 1136
rect 4242 1133 4249 1140
rect 4252 1136 4319 1160
rect 4351 1160 4523 1162
rect 4321 1138 4349 1142
rect 4351 1138 4431 1160
rect 4452 1158 4467 1160
rect 4321 1136 4431 1138
rect 4252 1132 4431 1136
rect 4225 1122 4255 1132
rect 4257 1122 4410 1132
rect 4418 1122 4448 1132
rect 4452 1122 4482 1136
rect 4510 1122 4523 1160
rect 4595 1166 4630 1174
rect 4595 1140 4596 1166
rect 4603 1140 4630 1166
rect 4538 1122 4568 1136
rect 4595 1132 4630 1140
rect 4632 1166 4673 1174
rect 4632 1140 4647 1166
rect 4654 1140 4673 1166
rect 4737 1162 4799 1174
rect 4811 1162 4886 1174
rect 4944 1162 5019 1174
rect 5031 1162 5062 1174
rect 5068 1162 5103 1174
rect 4737 1160 4899 1162
rect 4755 1141 4768 1160
rect 4783 1158 4798 1160
rect 4632 1132 4673 1140
rect 4756 1135 4768 1141
rect 4832 1142 4899 1160
rect 4931 1160 5103 1162
rect 4931 1142 5011 1160
rect 5032 1158 5047 1160
rect 4595 1122 4596 1132
rect 4611 1122 4624 1132
rect 4638 1122 4639 1132
rect 4654 1122 4667 1132
rect 4682 1122 4712 1135
rect 4756 1122 4798 1135
rect 4822 1133 4829 1140
rect 4832 1132 5011 1142
rect 4805 1131 4813 1132
rect 4832 1131 4835 1132
rect 4805 1124 4835 1131
rect 4837 1124 4990 1132
rect 5017 1131 5028 1132
rect 4998 1124 5028 1131
rect 4805 1122 5028 1124
rect 5032 1122 5062 1135
rect 5090 1122 5103 1160
rect 5175 1166 5210 1174
rect 5175 1140 5176 1166
rect 5183 1140 5210 1166
rect 5118 1122 5148 1135
rect 5175 1132 5210 1140
rect 5212 1166 5253 1174
rect 5212 1140 5227 1166
rect 5234 1140 5253 1166
rect 5317 1162 5379 1174
rect 5391 1162 5466 1174
rect 5524 1162 5599 1174
rect 5611 1162 5642 1174
rect 5648 1162 5683 1174
rect 5317 1160 5479 1162
rect 5335 1141 5348 1160
rect 5363 1158 5378 1160
rect 5212 1132 5253 1140
rect 5336 1135 5348 1141
rect 5412 1142 5479 1160
rect 5511 1160 5683 1162
rect 5511 1142 5591 1160
rect 5612 1158 5627 1160
rect 5175 1122 5176 1132
rect 5191 1122 5204 1132
rect 5218 1122 5219 1132
rect 5234 1122 5247 1132
rect 5262 1122 5292 1135
rect 5336 1122 5378 1135
rect 5402 1133 5409 1140
rect 5412 1132 5591 1142
rect 5385 1131 5393 1132
rect 5412 1131 5415 1132
rect 5385 1124 5415 1131
rect 5417 1124 5570 1132
rect 5597 1131 5608 1132
rect 5578 1124 5608 1131
rect 5385 1122 5608 1124
rect 5612 1122 5642 1135
rect 5670 1122 5683 1160
rect 5755 1166 5790 1174
rect 5755 1140 5756 1166
rect 5763 1140 5790 1166
rect 5698 1122 5728 1135
rect 5755 1132 5790 1140
rect 5792 1166 5833 1174
rect 5792 1140 5807 1166
rect 5814 1140 5833 1166
rect 5897 1162 5959 1174
rect 5971 1162 6046 1174
rect 6104 1162 6179 1174
rect 6191 1162 6222 1174
rect 6228 1162 6263 1174
rect 5897 1160 6059 1162
rect 5915 1141 5928 1160
rect 5943 1158 5958 1160
rect 5792 1132 5833 1140
rect 5916 1135 5928 1141
rect 5992 1142 6059 1160
rect 6091 1160 6263 1162
rect 6091 1142 6171 1160
rect 6192 1158 6207 1160
rect 5755 1122 5756 1132
rect 5771 1122 5784 1132
rect 5798 1122 5799 1132
rect 5814 1122 5827 1132
rect 5842 1122 5872 1135
rect 5916 1122 5958 1135
rect 5982 1133 5989 1140
rect 5992 1132 6171 1142
rect 5965 1131 5973 1132
rect 5992 1131 5995 1132
rect 5965 1124 5995 1131
rect 5997 1124 6150 1132
rect 6177 1131 6188 1132
rect 6158 1124 6188 1131
rect 5965 1122 6188 1124
rect 6192 1122 6222 1135
rect 6250 1122 6263 1160
rect 6335 1166 6370 1174
rect 6335 1140 6336 1166
rect 6343 1140 6370 1166
rect 6278 1122 6308 1135
rect 6335 1132 6370 1140
rect 6372 1166 6413 1174
rect 6372 1140 6387 1166
rect 6394 1140 6413 1166
rect 6477 1162 6539 1174
rect 6551 1162 6626 1174
rect 6684 1162 6759 1174
rect 6771 1162 6802 1174
rect 6808 1162 6843 1174
rect 6477 1160 6639 1162
rect 6495 1141 6508 1160
rect 6523 1158 6538 1160
rect 6372 1132 6413 1140
rect 6496 1135 6508 1141
rect 6572 1142 6639 1160
rect 6671 1160 6843 1162
rect 6671 1142 6751 1160
rect 6772 1158 6787 1160
rect 6335 1122 6336 1132
rect 6351 1122 6364 1132
rect 6378 1122 6379 1132
rect 6394 1122 6407 1132
rect 6422 1122 6452 1135
rect 6496 1122 6538 1135
rect 6562 1133 6569 1140
rect 6572 1132 6751 1142
rect 6545 1131 6553 1132
rect 6572 1131 6575 1132
rect 6545 1124 6575 1131
rect 6577 1124 6730 1132
rect 6757 1131 6768 1132
rect 6738 1124 6768 1131
rect 6545 1122 6768 1124
rect 6772 1122 6802 1135
rect 6830 1122 6843 1160
rect 6915 1166 6950 1174
rect 6915 1140 6916 1166
rect 6923 1140 6950 1166
rect 6858 1122 6888 1135
rect 6915 1132 6950 1140
rect 6915 1122 6916 1132
rect 6931 1122 6944 1132
rect -2 1116 6944 1122
rect -1 1108 6944 1116
rect 14 1078 27 1108
rect 42 1090 72 1108
rect 115 1094 129 1108
rect 165 1094 385 1108
rect 116 1092 129 1094
rect 82 1080 97 1092
rect 79 1078 101 1080
rect 106 1078 136 1092
rect 197 1090 350 1094
rect 179 1078 371 1090
rect 414 1078 444 1092
rect 450 1078 463 1108
rect 478 1090 508 1108
rect 551 1078 564 1108
rect 594 1078 607 1108
rect 622 1090 652 1108
rect 695 1094 709 1108
rect 745 1094 965 1108
rect 696 1092 709 1094
rect 662 1080 677 1092
rect 659 1078 681 1080
rect 686 1078 716 1092
rect 777 1090 930 1094
rect 759 1078 951 1090
rect 994 1078 1024 1092
rect 1030 1078 1043 1108
rect 1058 1090 1088 1108
rect 1131 1078 1144 1108
rect 1174 1078 1187 1108
rect 1202 1090 1232 1108
rect 1275 1094 1289 1108
rect 1325 1094 1545 1108
rect 1276 1092 1289 1094
rect 1242 1080 1257 1092
rect 1239 1078 1261 1080
rect 1266 1078 1296 1092
rect 1357 1090 1510 1094
rect 1339 1078 1531 1090
rect 1574 1078 1604 1092
rect 1610 1078 1623 1108
rect 1638 1090 1668 1108
rect 1711 1078 1724 1108
rect 1754 1078 1767 1108
rect 1782 1090 1812 1108
rect 1855 1094 1869 1108
rect 1905 1094 2125 1108
rect 1856 1092 1869 1094
rect 1822 1080 1837 1092
rect 1819 1078 1841 1080
rect 1846 1078 1876 1092
rect 1937 1090 2090 1094
rect 1919 1078 2111 1090
rect 2154 1078 2184 1092
rect 2190 1078 2203 1108
rect 2218 1090 2248 1108
rect 2291 1078 2304 1108
rect 2334 1078 2347 1108
rect 2362 1090 2392 1108
rect 2435 1094 2449 1108
rect 2485 1094 2705 1108
rect 2436 1092 2449 1094
rect 2402 1080 2417 1092
rect 2399 1078 2421 1080
rect 2426 1078 2456 1092
rect 2517 1090 2670 1094
rect 2499 1078 2691 1090
rect 2734 1078 2764 1092
rect 2770 1078 2783 1108
rect 2798 1090 2828 1108
rect 2871 1078 2884 1108
rect 2914 1078 2927 1108
rect 2942 1090 2972 1108
rect 3015 1094 3029 1108
rect 3065 1094 3285 1108
rect 3016 1092 3029 1094
rect 2982 1080 2997 1092
rect 2979 1078 3001 1080
rect 3006 1078 3036 1092
rect 3097 1090 3250 1094
rect 3079 1078 3271 1090
rect 3314 1078 3344 1092
rect 3350 1078 3363 1108
rect 3378 1090 3408 1108
rect 3451 1078 3464 1108
rect 3494 1078 3507 1108
rect 3522 1090 3552 1108
rect 3595 1094 3609 1108
rect 3645 1094 3865 1108
rect 3596 1092 3609 1094
rect 3562 1080 3577 1092
rect 3559 1078 3581 1080
rect 3586 1078 3616 1092
rect 3677 1090 3830 1094
rect 3659 1078 3851 1090
rect 3894 1078 3924 1092
rect 3930 1078 3943 1108
rect 3958 1090 3988 1108
rect 4031 1078 4044 1108
rect 4074 1078 4087 1108
rect 4102 1090 4132 1108
rect 4175 1094 4189 1108
rect 4225 1094 4445 1108
rect 4176 1092 4189 1094
rect 4142 1080 4157 1092
rect 4139 1078 4161 1080
rect 4166 1078 4196 1092
rect 4257 1090 4410 1094
rect 4239 1078 4431 1090
rect 4474 1078 4504 1092
rect 4510 1078 4523 1108
rect 4538 1090 4568 1108
rect 4611 1078 4624 1108
rect -1 1077 4624 1078
rect 4654 1077 4667 1108
rect 4682 1090 4712 1108
rect 4756 1091 4769 1108
rect 4805 1094 5025 1108
rect 4722 1079 4737 1091
rect 4719 1077 4741 1079
rect 4746 1077 4776 1091
rect 4837 1089 4990 1094
rect 4819 1077 5011 1089
rect 5054 1077 5084 1091
rect 5090 1077 5103 1108
rect 5118 1090 5148 1108
rect 5191 1077 5204 1108
rect 5234 1077 5247 1108
rect 5262 1090 5292 1108
rect 5336 1091 5349 1108
rect 5385 1094 5605 1108
rect 5302 1079 5317 1091
rect 5299 1077 5321 1079
rect 5326 1077 5356 1091
rect 5417 1089 5570 1094
rect 5399 1077 5591 1089
rect 5634 1077 5664 1091
rect 5670 1077 5683 1108
rect 5698 1090 5728 1108
rect 5771 1077 5784 1108
rect 5814 1077 5827 1108
rect 5842 1090 5872 1108
rect 5916 1091 5929 1108
rect 5965 1094 6185 1108
rect 5882 1079 5897 1091
rect 5879 1077 5901 1079
rect 5906 1077 5936 1091
rect 5997 1089 6150 1094
rect 5979 1077 6171 1089
rect 6214 1077 6244 1091
rect 6250 1077 6263 1108
rect 6278 1090 6308 1108
rect 6351 1077 6364 1108
rect 6394 1077 6407 1108
rect 6422 1090 6452 1108
rect 6496 1091 6509 1108
rect 6545 1094 6765 1108
rect 6462 1079 6477 1091
rect 6459 1077 6481 1079
rect 6486 1077 6516 1091
rect 6577 1089 6730 1094
rect 6559 1077 6751 1089
rect 6794 1077 6824 1091
rect 6830 1077 6843 1108
rect 6858 1090 6888 1108
rect 6931 1077 6944 1108
rect -1 1064 6944 1077
rect 14 960 27 1064
rect 72 1042 73 1052
rect 88 1042 101 1052
rect 72 1038 101 1042
rect 106 1038 136 1064
rect 154 1050 170 1052
rect 242 1050 295 1064
rect 243 1048 307 1050
rect 350 1048 365 1064
rect 414 1061 444 1064
rect 414 1058 450 1061
rect 380 1050 396 1052
rect 154 1038 169 1042
rect 72 1036 169 1038
rect 197 1036 365 1048
rect 381 1038 396 1042
rect 414 1039 453 1058
rect 472 1052 479 1053
rect 478 1045 479 1052
rect 462 1042 463 1045
rect 478 1042 491 1045
rect 414 1038 444 1039
rect 453 1038 459 1039
rect 462 1038 491 1042
rect 381 1037 491 1038
rect 381 1036 497 1037
rect 56 1028 107 1036
rect 56 1016 81 1028
rect 88 1016 107 1028
rect 138 1028 188 1036
rect 138 1020 154 1028
rect 161 1026 188 1028
rect 197 1026 418 1036
rect 161 1016 418 1026
rect 447 1028 497 1036
rect 447 1019 463 1028
rect 56 1008 107 1016
rect 154 1008 418 1016
rect 444 1016 463 1019
rect 470 1016 497 1028
rect 444 1008 497 1016
rect 72 1000 73 1008
rect 88 1000 101 1008
rect 72 992 88 1000
rect 69 985 88 988
rect 69 976 91 985
rect 42 966 91 976
rect 42 960 72 966
rect 91 961 96 966
rect 14 944 88 960
rect 106 952 136 1008
rect 171 998 379 1008
rect 414 1004 459 1008
rect 462 1007 463 1008
rect 478 1007 491 1008
rect 197 968 386 998
rect 212 965 386 968
rect 205 962 386 965
rect 14 942 27 944
rect 42 942 76 944
rect 14 926 88 942
rect 115 938 128 952
rect 143 938 159 954
rect 205 949 216 962
rect -2 904 -1 920
rect 14 904 27 926
rect 42 904 72 926
rect 115 922 177 938
rect 205 931 216 947
rect 221 942 231 962
rect 241 942 255 962
rect 258 949 267 962
rect 283 949 292 962
rect 221 931 255 942
rect 258 931 267 947
rect 283 931 292 947
rect 299 942 309 962
rect 319 942 333 962
rect 334 949 345 962
rect 299 931 333 942
rect 334 931 345 947
rect 391 938 407 954
rect 414 952 444 1004
rect 478 1000 479 1007
rect 463 992 479 1000
rect 450 960 463 979
rect 478 960 508 976
rect 450 944 524 960
rect 450 942 463 944
rect 478 942 512 944
rect 115 920 128 922
rect 143 920 177 922
rect 115 904 177 920
rect 221 915 237 918
rect 299 915 329 926
rect 377 922 423 938
rect 450 926 524 942
rect 377 920 411 922
rect 376 904 423 920
rect 450 904 463 926
rect 478 904 508 926
rect 535 904 536 920
rect 551 904 564 1064
rect 594 960 607 1064
rect 652 1042 653 1052
rect 668 1042 681 1052
rect 652 1038 681 1042
rect 686 1038 716 1064
rect 734 1050 750 1052
rect 822 1050 875 1064
rect 823 1048 887 1050
rect 930 1048 945 1064
rect 994 1061 1024 1064
rect 994 1058 1030 1061
rect 960 1050 976 1052
rect 734 1038 749 1042
rect 652 1036 749 1038
rect 777 1036 945 1048
rect 961 1038 976 1042
rect 994 1039 1033 1058
rect 1052 1052 1059 1053
rect 1058 1045 1059 1052
rect 1042 1042 1043 1045
rect 1058 1042 1071 1045
rect 994 1038 1024 1039
rect 1033 1038 1039 1039
rect 1042 1038 1071 1042
rect 961 1037 1071 1038
rect 961 1036 1077 1037
rect 636 1028 687 1036
rect 636 1016 661 1028
rect 668 1016 687 1028
rect 718 1028 768 1036
rect 718 1020 734 1028
rect 741 1026 768 1028
rect 777 1026 998 1036
rect 741 1016 998 1026
rect 1027 1028 1077 1036
rect 1027 1019 1043 1028
rect 636 1008 687 1016
rect 734 1008 998 1016
rect 1024 1016 1043 1019
rect 1050 1016 1077 1028
rect 1024 1008 1077 1016
rect 652 1000 653 1008
rect 668 1000 681 1008
rect 652 992 668 1000
rect 649 985 668 988
rect 649 976 671 985
rect 622 966 671 976
rect 622 960 652 966
rect 671 961 676 966
rect 594 944 668 960
rect 686 952 716 1008
rect 751 998 959 1008
rect 994 1004 1039 1008
rect 1042 1007 1043 1008
rect 1058 1007 1071 1008
rect 777 968 966 998
rect 792 965 966 968
rect 785 962 966 965
rect 594 942 607 944
rect 622 942 656 944
rect 594 926 668 942
rect 695 938 708 952
rect 723 938 739 954
rect 785 949 796 962
rect 578 904 579 920
rect 594 904 607 926
rect 622 904 652 926
rect 695 922 757 938
rect 785 931 796 947
rect 801 942 811 962
rect 821 942 835 962
rect 838 949 847 962
rect 863 949 872 962
rect 801 931 835 942
rect 838 931 847 947
rect 863 931 872 947
rect 879 942 889 962
rect 899 942 913 962
rect 914 949 925 962
rect 879 931 913 942
rect 914 931 925 947
rect 971 938 987 954
rect 994 952 1024 1004
rect 1058 1000 1059 1007
rect 1043 992 1059 1000
rect 1030 960 1043 979
rect 1058 960 1088 976
rect 1030 944 1104 960
rect 1030 942 1043 944
rect 1058 942 1092 944
rect 695 920 708 922
rect 723 920 757 922
rect 695 904 757 920
rect 801 915 817 918
rect 879 915 909 926
rect 957 922 1003 938
rect 1030 926 1104 942
rect 957 920 991 922
rect 956 904 1003 920
rect 1030 904 1043 926
rect 1058 904 1088 926
rect 1115 904 1116 920
rect 1131 904 1144 1064
rect 1174 960 1187 1064
rect 1232 1042 1233 1052
rect 1248 1042 1261 1052
rect 1232 1038 1261 1042
rect 1266 1038 1296 1064
rect 1314 1050 1330 1052
rect 1402 1050 1455 1064
rect 1403 1048 1467 1050
rect 1510 1048 1525 1064
rect 1574 1061 1604 1064
rect 1574 1058 1610 1061
rect 1540 1050 1556 1052
rect 1314 1038 1329 1042
rect 1232 1036 1329 1038
rect 1357 1036 1525 1048
rect 1541 1038 1556 1042
rect 1574 1039 1613 1058
rect 1632 1052 1639 1053
rect 1638 1045 1639 1052
rect 1622 1042 1623 1045
rect 1638 1042 1651 1045
rect 1574 1038 1604 1039
rect 1613 1038 1619 1039
rect 1622 1038 1651 1042
rect 1541 1037 1651 1038
rect 1541 1036 1657 1037
rect 1216 1028 1267 1036
rect 1216 1016 1241 1028
rect 1248 1016 1267 1028
rect 1298 1028 1348 1036
rect 1298 1020 1314 1028
rect 1321 1026 1348 1028
rect 1357 1026 1578 1036
rect 1321 1016 1578 1026
rect 1607 1028 1657 1036
rect 1607 1019 1623 1028
rect 1216 1008 1267 1016
rect 1314 1008 1578 1016
rect 1604 1016 1623 1019
rect 1630 1016 1657 1028
rect 1604 1008 1657 1016
rect 1232 1000 1233 1008
rect 1248 1000 1261 1008
rect 1232 992 1248 1000
rect 1229 985 1248 988
rect 1229 976 1251 985
rect 1202 966 1251 976
rect 1202 960 1232 966
rect 1251 961 1256 966
rect 1174 944 1248 960
rect 1266 952 1296 1008
rect 1331 998 1539 1008
rect 1574 1004 1619 1008
rect 1622 1007 1623 1008
rect 1638 1007 1651 1008
rect 1357 968 1546 998
rect 1372 965 1546 968
rect 1365 962 1546 965
rect 1174 942 1187 944
rect 1202 942 1236 944
rect 1174 926 1248 942
rect 1275 938 1288 952
rect 1303 938 1319 954
rect 1365 949 1376 962
rect 1158 904 1159 920
rect 1174 904 1187 926
rect 1202 904 1232 926
rect 1275 922 1337 938
rect 1365 931 1376 947
rect 1381 942 1391 962
rect 1401 942 1415 962
rect 1418 949 1427 962
rect 1443 949 1452 962
rect 1381 931 1415 942
rect 1418 931 1427 947
rect 1443 931 1452 947
rect 1459 942 1469 962
rect 1479 942 1493 962
rect 1494 949 1505 962
rect 1459 931 1493 942
rect 1494 931 1505 947
rect 1551 938 1567 954
rect 1574 952 1604 1004
rect 1638 1000 1639 1007
rect 1623 992 1639 1000
rect 1610 960 1623 979
rect 1638 960 1668 976
rect 1610 944 1684 960
rect 1610 942 1623 944
rect 1638 942 1672 944
rect 1275 920 1288 922
rect 1303 920 1337 922
rect 1275 904 1337 920
rect 1381 915 1397 918
rect 1459 915 1489 926
rect 1537 922 1583 938
rect 1610 926 1684 942
rect 1537 920 1571 922
rect 1536 904 1583 920
rect 1610 904 1623 926
rect 1638 904 1668 926
rect 1695 904 1696 920
rect 1711 904 1724 1064
rect 1754 960 1767 1064
rect 1812 1042 1813 1052
rect 1828 1042 1841 1052
rect 1812 1038 1841 1042
rect 1846 1038 1876 1064
rect 1894 1050 1910 1052
rect 1982 1050 2035 1064
rect 1983 1048 2047 1050
rect 2090 1048 2105 1064
rect 2154 1061 2184 1064
rect 2154 1058 2190 1061
rect 2120 1050 2136 1052
rect 1894 1038 1909 1042
rect 1812 1036 1909 1038
rect 1937 1036 2105 1048
rect 2121 1038 2136 1042
rect 2154 1039 2193 1058
rect 2212 1052 2219 1053
rect 2218 1045 2219 1052
rect 2202 1042 2203 1045
rect 2218 1042 2231 1045
rect 2154 1038 2184 1039
rect 2193 1038 2199 1039
rect 2202 1038 2231 1042
rect 2121 1037 2231 1038
rect 2121 1036 2237 1037
rect 1796 1028 1847 1036
rect 1796 1016 1821 1028
rect 1828 1016 1847 1028
rect 1878 1028 1928 1036
rect 1878 1020 1894 1028
rect 1901 1026 1928 1028
rect 1937 1026 2158 1036
rect 1901 1016 2158 1026
rect 2187 1028 2237 1036
rect 2187 1019 2203 1028
rect 1796 1008 1847 1016
rect 1894 1008 2158 1016
rect 2184 1016 2203 1019
rect 2210 1016 2237 1028
rect 2184 1008 2237 1016
rect 1812 1000 1813 1008
rect 1828 1000 1841 1008
rect 1812 992 1828 1000
rect 1809 985 1828 988
rect 1809 976 1831 985
rect 1782 966 1831 976
rect 1782 960 1812 966
rect 1831 961 1836 966
rect 1754 944 1828 960
rect 1846 952 1876 1008
rect 1911 998 2119 1008
rect 2154 1004 2199 1008
rect 2202 1007 2203 1008
rect 2218 1007 2231 1008
rect 1937 968 2126 998
rect 1952 965 2126 968
rect 1945 962 2126 965
rect 1754 942 1767 944
rect 1782 942 1816 944
rect 1754 926 1828 942
rect 1855 938 1868 952
rect 1883 938 1899 954
rect 1945 949 1956 962
rect 1738 904 1739 920
rect 1754 904 1767 926
rect 1782 904 1812 926
rect 1855 922 1917 938
rect 1945 931 1956 947
rect 1961 942 1971 962
rect 1981 942 1995 962
rect 1998 949 2007 962
rect 2023 949 2032 962
rect 1961 931 1995 942
rect 1998 931 2007 947
rect 2023 931 2032 947
rect 2039 942 2049 962
rect 2059 942 2073 962
rect 2074 949 2085 962
rect 2039 931 2073 942
rect 2074 931 2085 947
rect 2131 938 2147 954
rect 2154 952 2184 1004
rect 2218 1000 2219 1007
rect 2203 992 2219 1000
rect 2190 960 2203 979
rect 2218 960 2248 976
rect 2190 944 2264 960
rect 2190 942 2203 944
rect 2218 942 2252 944
rect 1855 920 1868 922
rect 1883 920 1917 922
rect 1855 904 1917 920
rect 1961 915 1977 918
rect 2039 915 2069 926
rect 2117 922 2163 938
rect 2190 926 2264 942
rect 2117 920 2151 922
rect 2116 904 2163 920
rect 2190 904 2203 926
rect 2218 904 2248 926
rect 2275 904 2276 920
rect 2291 904 2304 1064
rect 2334 960 2347 1064
rect 2392 1042 2393 1052
rect 2408 1042 2421 1052
rect 2392 1038 2421 1042
rect 2426 1038 2456 1064
rect 2474 1050 2490 1052
rect 2562 1050 2615 1064
rect 2563 1048 2627 1050
rect 2670 1048 2685 1064
rect 2734 1061 2764 1064
rect 2734 1058 2770 1061
rect 2700 1050 2716 1052
rect 2474 1038 2489 1042
rect 2392 1036 2489 1038
rect 2517 1036 2685 1048
rect 2701 1038 2716 1042
rect 2734 1039 2773 1058
rect 2792 1052 2799 1053
rect 2798 1045 2799 1052
rect 2782 1042 2783 1045
rect 2798 1042 2811 1045
rect 2734 1038 2764 1039
rect 2773 1038 2779 1039
rect 2782 1038 2811 1042
rect 2701 1037 2811 1038
rect 2701 1036 2817 1037
rect 2376 1028 2427 1036
rect 2376 1016 2401 1028
rect 2408 1016 2427 1028
rect 2458 1028 2508 1036
rect 2458 1020 2474 1028
rect 2481 1026 2508 1028
rect 2517 1026 2738 1036
rect 2481 1016 2738 1026
rect 2767 1028 2817 1036
rect 2767 1019 2783 1028
rect 2376 1008 2427 1016
rect 2474 1008 2738 1016
rect 2764 1016 2783 1019
rect 2790 1016 2817 1028
rect 2764 1008 2817 1016
rect 2392 1000 2393 1008
rect 2408 1000 2421 1008
rect 2392 992 2408 1000
rect 2389 985 2408 988
rect 2389 976 2411 985
rect 2362 966 2411 976
rect 2362 960 2392 966
rect 2411 961 2416 966
rect 2334 944 2408 960
rect 2426 952 2456 1008
rect 2491 998 2699 1008
rect 2734 1004 2779 1008
rect 2782 1007 2783 1008
rect 2798 1007 2811 1008
rect 2517 968 2706 998
rect 2532 965 2706 968
rect 2525 962 2706 965
rect 2334 942 2347 944
rect 2362 942 2396 944
rect 2334 926 2408 942
rect 2435 938 2448 952
rect 2463 938 2479 954
rect 2525 949 2536 962
rect 2318 904 2319 920
rect 2334 904 2347 926
rect 2362 904 2392 926
rect 2435 922 2497 938
rect 2525 931 2536 947
rect 2541 942 2551 962
rect 2561 942 2575 962
rect 2578 949 2587 962
rect 2603 949 2612 962
rect 2541 931 2575 942
rect 2578 931 2587 947
rect 2603 931 2612 947
rect 2619 942 2629 962
rect 2639 942 2653 962
rect 2654 949 2665 962
rect 2619 931 2653 942
rect 2654 931 2665 947
rect 2711 938 2727 954
rect 2734 952 2764 1004
rect 2798 1000 2799 1007
rect 2783 992 2799 1000
rect 2770 960 2783 979
rect 2798 960 2828 976
rect 2770 944 2844 960
rect 2770 942 2783 944
rect 2798 942 2832 944
rect 2435 920 2448 922
rect 2463 920 2497 922
rect 2435 904 2497 920
rect 2541 915 2557 918
rect 2619 915 2649 926
rect 2697 922 2743 938
rect 2770 926 2844 942
rect 2697 920 2731 922
rect 2696 904 2743 920
rect 2770 904 2783 926
rect 2798 904 2828 926
rect 2855 904 2856 920
rect 2871 904 2884 1064
rect 2914 960 2927 1064
rect 2972 1042 2973 1052
rect 2988 1042 3001 1052
rect 2972 1038 3001 1042
rect 3006 1038 3036 1064
rect 3054 1050 3070 1052
rect 3142 1050 3195 1064
rect 3143 1048 3205 1050
rect 3250 1048 3265 1064
rect 3314 1061 3344 1064
rect 3314 1058 3350 1061
rect 3280 1050 3296 1052
rect 3054 1038 3069 1042
rect 2972 1036 3069 1038
rect 3097 1036 3265 1048
rect 3281 1038 3296 1042
rect 3314 1039 3353 1058
rect 3372 1052 3379 1053
rect 3378 1045 3379 1052
rect 3362 1042 3363 1045
rect 3378 1042 3391 1045
rect 3314 1038 3344 1039
rect 3353 1038 3359 1039
rect 3362 1038 3391 1042
rect 3281 1037 3391 1038
rect 3281 1036 3397 1037
rect 2956 1028 3007 1036
rect 2956 1016 2981 1028
rect 2988 1016 3007 1028
rect 3038 1028 3088 1036
rect 3038 1020 3054 1028
rect 3061 1026 3088 1028
rect 3097 1026 3318 1036
rect 3061 1016 3318 1026
rect 3347 1028 3397 1036
rect 3347 1019 3363 1028
rect 2956 1008 3007 1016
rect 3054 1008 3318 1016
rect 3344 1016 3363 1019
rect 3370 1016 3397 1028
rect 3344 1008 3397 1016
rect 2972 1000 2973 1008
rect 2988 1000 3001 1008
rect 2972 992 2988 1000
rect 2969 985 2988 988
rect 2969 976 2991 985
rect 2942 966 2991 976
rect 2942 960 2972 966
rect 2991 961 2996 966
rect 2914 944 2988 960
rect 3006 952 3036 1008
rect 3071 998 3279 1008
rect 3314 1004 3359 1008
rect 3362 1007 3363 1008
rect 3378 1007 3391 1008
rect 3097 968 3286 998
rect 3112 965 3286 968
rect 3105 962 3286 965
rect 2914 942 2927 944
rect 2942 942 2976 944
rect 2914 926 2988 942
rect 3015 938 3028 952
rect 3043 938 3059 954
rect 3105 949 3116 962
rect 2898 904 2899 920
rect 2914 904 2927 926
rect 2942 904 2972 926
rect 3015 922 3077 938
rect 3105 931 3116 947
rect 3121 942 3131 962
rect 3141 942 3155 962
rect 3158 949 3167 962
rect 3183 949 3192 962
rect 3121 931 3155 942
rect 3158 931 3167 947
rect 3183 931 3192 947
rect 3199 942 3209 962
rect 3219 942 3233 962
rect 3234 949 3245 962
rect 3199 931 3233 942
rect 3234 931 3245 947
rect 3291 938 3307 954
rect 3314 952 3344 1004
rect 3378 1000 3379 1007
rect 3363 992 3379 1000
rect 3350 960 3363 979
rect 3378 960 3408 976
rect 3350 944 3424 960
rect 3350 942 3363 944
rect 3378 942 3412 944
rect 3015 920 3028 922
rect 3043 920 3077 922
rect 3015 904 3077 920
rect 3121 915 3137 918
rect 3199 915 3229 926
rect 3277 922 3323 938
rect 3350 926 3424 942
rect 3277 920 3311 922
rect 3276 904 3323 920
rect 3350 904 3363 926
rect 3378 904 3408 926
rect 3435 904 3436 920
rect 3451 904 3464 1064
rect 3494 960 3507 1064
rect 3552 1042 3553 1052
rect 3568 1042 3581 1052
rect 3552 1038 3581 1042
rect 3586 1038 3616 1064
rect 3634 1050 3650 1052
rect 3722 1050 3775 1064
rect 3723 1048 3787 1050
rect 3830 1048 3845 1064
rect 3894 1061 3924 1064
rect 3894 1058 3930 1061
rect 3860 1050 3876 1052
rect 3634 1038 3649 1042
rect 3552 1036 3649 1038
rect 3677 1036 3845 1048
rect 3861 1038 3876 1042
rect 3894 1039 3933 1058
rect 3952 1052 3959 1053
rect 3958 1045 3959 1052
rect 3942 1042 3943 1045
rect 3958 1042 3971 1045
rect 3894 1038 3924 1039
rect 3933 1038 3939 1039
rect 3942 1038 3971 1042
rect 3861 1037 3971 1038
rect 3861 1036 3977 1037
rect 3536 1028 3587 1036
rect 3536 1016 3561 1028
rect 3568 1016 3587 1028
rect 3618 1028 3668 1036
rect 3618 1020 3634 1028
rect 3641 1026 3668 1028
rect 3677 1026 3898 1036
rect 3641 1016 3898 1026
rect 3927 1028 3977 1036
rect 3927 1019 3943 1028
rect 3536 1008 3587 1016
rect 3634 1008 3898 1016
rect 3924 1016 3943 1019
rect 3950 1016 3977 1028
rect 3924 1008 3977 1016
rect 3552 1000 3553 1008
rect 3568 1000 3581 1008
rect 3552 992 3568 1000
rect 3549 985 3568 988
rect 3549 976 3571 985
rect 3522 966 3571 976
rect 3522 960 3552 966
rect 3571 961 3576 966
rect 3494 944 3568 960
rect 3586 952 3616 1008
rect 3651 998 3859 1008
rect 3894 1004 3939 1008
rect 3942 1007 3943 1008
rect 3958 1007 3971 1008
rect 3677 968 3866 998
rect 3692 965 3866 968
rect 3685 962 3866 965
rect 3494 942 3507 944
rect 3522 942 3556 944
rect 3494 926 3568 942
rect 3595 938 3608 952
rect 3623 938 3639 954
rect 3685 949 3696 962
rect 3478 904 3479 920
rect 3494 904 3507 926
rect 3522 904 3552 926
rect 3595 922 3657 938
rect 3685 931 3696 947
rect 3701 942 3711 962
rect 3721 942 3735 962
rect 3738 949 3747 962
rect 3763 949 3772 962
rect 3701 931 3735 942
rect 3738 931 3747 947
rect 3763 931 3772 947
rect 3779 942 3789 962
rect 3799 942 3813 962
rect 3814 949 3825 962
rect 3779 931 3813 942
rect 3814 931 3825 947
rect 3871 938 3887 954
rect 3894 952 3924 1004
rect 3958 1000 3959 1007
rect 3943 992 3959 1000
rect 3930 960 3943 979
rect 3958 960 3988 976
rect 3930 944 4004 960
rect 3930 942 3943 944
rect 3958 942 3992 944
rect 3595 920 3608 922
rect 3623 920 3657 922
rect 3595 904 3657 920
rect 3701 915 3717 918
rect 3779 915 3809 926
rect 3857 922 3903 938
rect 3930 926 4004 942
rect 3857 920 3891 922
rect 3856 904 3903 920
rect 3930 904 3943 926
rect 3958 904 3988 926
rect 4015 904 4016 920
rect 4031 904 4044 1064
rect 4074 960 4087 1064
rect 4132 1042 4133 1052
rect 4148 1042 4161 1052
rect 4132 1038 4161 1042
rect 4166 1038 4196 1064
rect 4214 1050 4230 1052
rect 4302 1050 4355 1064
rect 4303 1048 4367 1050
rect 4410 1048 4425 1064
rect 4474 1061 4504 1064
rect 4611 1063 6944 1064
rect 4474 1058 4510 1061
rect 4440 1050 4456 1052
rect 4214 1038 4229 1042
rect 4132 1036 4229 1038
rect 4257 1036 4425 1048
rect 4441 1038 4456 1042
rect 4474 1039 4513 1058
rect 4532 1052 4539 1053
rect 4538 1045 4539 1052
rect 4522 1042 4523 1045
rect 4538 1042 4551 1045
rect 4474 1038 4504 1039
rect 4513 1038 4519 1039
rect 4522 1038 4551 1042
rect 4441 1037 4551 1038
rect 4441 1036 4557 1037
rect 4116 1028 4167 1036
rect 4116 1016 4141 1028
rect 4148 1016 4167 1028
rect 4198 1028 4248 1036
rect 4198 1020 4214 1028
rect 4221 1026 4248 1028
rect 4257 1026 4478 1036
rect 4221 1016 4478 1026
rect 4507 1028 4557 1036
rect 4507 1019 4523 1028
rect 4116 1008 4167 1016
rect 4214 1008 4478 1016
rect 4504 1016 4523 1019
rect 4530 1016 4557 1028
rect 4504 1008 4557 1016
rect 4132 1000 4133 1008
rect 4148 1000 4161 1008
rect 4132 992 4148 1000
rect 4129 985 4148 988
rect 4129 976 4151 985
rect 4102 966 4151 976
rect 4102 960 4132 966
rect 4151 961 4156 966
rect 4074 944 4148 960
rect 4166 952 4196 1008
rect 4231 998 4439 1008
rect 4474 1004 4519 1008
rect 4522 1007 4523 1008
rect 4538 1007 4551 1008
rect 4257 968 4446 998
rect 4272 965 4446 968
rect 4265 962 4446 965
rect 4074 942 4087 944
rect 4102 942 4136 944
rect 4074 926 4148 942
rect 4175 938 4188 952
rect 4203 938 4219 954
rect 4265 949 4276 962
rect 4058 904 4059 920
rect 4074 904 4087 926
rect 4102 904 4132 926
rect 4175 922 4237 938
rect 4265 931 4276 947
rect 4281 942 4291 962
rect 4301 942 4315 962
rect 4318 949 4327 962
rect 4343 949 4352 962
rect 4281 931 4315 942
rect 4318 931 4327 947
rect 4343 931 4352 947
rect 4359 942 4369 962
rect 4379 942 4393 962
rect 4394 949 4405 962
rect 4359 931 4393 942
rect 4394 931 4405 947
rect 4451 938 4467 954
rect 4474 952 4504 1004
rect 4538 1000 4539 1007
rect 4523 992 4539 1000
rect 4510 960 4523 979
rect 4538 960 4568 976
rect 4510 944 4584 960
rect 4510 942 4523 944
rect 4538 942 4572 944
rect 4175 920 4188 922
rect 4203 920 4237 922
rect 4175 904 4237 920
rect 4281 915 4297 918
rect 4359 915 4389 926
rect 4437 922 4483 938
rect 4510 926 4584 942
rect 4437 920 4471 922
rect 4436 904 4483 920
rect 4510 904 4523 926
rect 4538 904 4568 926
rect 4595 904 4596 920
rect 4611 904 4624 1063
rect 4654 959 4667 1063
rect 4712 1041 4713 1051
rect 4733 1049 4741 1051
rect 4731 1047 4741 1049
rect 4728 1041 4741 1047
rect 4712 1037 4741 1041
rect 4746 1037 4776 1063
rect 4794 1049 4810 1051
rect 4882 1049 4933 1063
rect 4883 1047 4947 1049
rect 4990 1047 5005 1063
rect 5054 1060 5084 1063
rect 5054 1057 5090 1060
rect 5020 1049 5036 1051
rect 4794 1037 4809 1041
rect 4712 1035 4809 1037
rect 4837 1035 5005 1047
rect 5021 1037 5036 1041
rect 5054 1038 5093 1057
rect 5112 1051 5119 1052
rect 5118 1044 5119 1051
rect 5102 1041 5103 1044
rect 5118 1041 5131 1044
rect 5054 1037 5084 1038
rect 5093 1037 5099 1038
rect 5102 1037 5131 1041
rect 5021 1036 5131 1037
rect 5021 1035 5137 1036
rect 4696 1027 4747 1035
rect 4696 1015 4721 1027
rect 4728 1015 4747 1027
rect 4778 1027 4828 1035
rect 4778 1019 4794 1027
rect 4801 1025 4828 1027
rect 4837 1025 5058 1035
rect 4801 1015 5058 1025
rect 5087 1027 5137 1035
rect 5087 1018 5103 1027
rect 4696 1007 4747 1015
rect 4794 1007 5058 1015
rect 5084 1015 5103 1018
rect 5110 1015 5137 1027
rect 5084 1007 5137 1015
rect 4712 999 4713 1007
rect 4728 999 4741 1007
rect 4712 991 4728 999
rect 4709 984 4728 987
rect 4709 975 4731 984
rect 4682 965 4731 975
rect 4682 959 4712 965
rect 4731 960 4736 965
rect 4654 943 4728 959
rect 4746 951 4776 1007
rect 4811 997 5019 1007
rect 5054 1003 5099 1007
rect 5102 1006 5103 1007
rect 5118 1006 5131 1007
rect 4837 967 5026 997
rect 4852 964 5026 967
rect 4845 961 5026 964
rect 4654 941 4667 943
rect 4682 941 4716 943
rect 4654 925 4728 941
rect 4755 937 4768 951
rect 4783 937 4799 953
rect 4845 948 4856 961
rect -8 896 33 904
rect -8 870 7 896
rect 14 870 33 896
rect 97 892 159 904
rect 171 892 246 904
rect 304 892 379 904
rect 391 892 422 904
rect 428 892 463 904
rect 97 890 259 892
rect -8 862 33 870
rect 115 866 128 890
rect 143 888 158 890
rect -2 852 -1 862
rect 14 852 27 862
rect 42 852 72 866
rect 115 852 158 866
rect 182 863 189 870
rect 192 866 259 890
rect 291 890 463 892
rect 261 868 289 872
rect 291 868 371 890
rect 392 888 407 890
rect 261 866 371 868
rect 192 862 371 866
rect 165 852 195 862
rect 197 852 350 862
rect 358 852 388 862
rect 392 852 422 866
rect 450 852 463 890
rect 535 896 570 904
rect 535 870 536 896
rect 543 870 570 896
rect 478 852 508 866
rect 535 862 570 870
rect 572 896 613 904
rect 572 870 587 896
rect 594 870 613 896
rect 677 892 739 904
rect 751 892 826 904
rect 884 892 959 904
rect 971 892 1002 904
rect 1008 892 1043 904
rect 677 890 839 892
rect 572 862 613 870
rect 695 866 708 890
rect 723 888 738 890
rect 535 852 536 862
rect 551 852 564 862
rect 578 852 579 862
rect 594 852 607 862
rect 622 852 652 866
rect 695 852 738 866
rect 762 863 769 870
rect 772 866 839 890
rect 871 890 1043 892
rect 841 868 869 872
rect 871 868 951 890
rect 972 888 987 890
rect 841 866 951 868
rect 772 862 951 866
rect 745 852 775 862
rect 777 852 930 862
rect 938 852 968 862
rect 972 852 1002 866
rect 1030 852 1043 890
rect 1115 896 1150 904
rect 1115 870 1116 896
rect 1123 870 1150 896
rect 1058 852 1088 866
rect 1115 862 1150 870
rect 1152 896 1193 904
rect 1152 870 1167 896
rect 1174 870 1193 896
rect 1257 892 1319 904
rect 1331 892 1406 904
rect 1464 892 1539 904
rect 1551 892 1582 904
rect 1588 892 1623 904
rect 1257 890 1419 892
rect 1152 862 1193 870
rect 1275 866 1288 890
rect 1303 888 1318 890
rect 1115 852 1116 862
rect 1131 852 1144 862
rect 1158 852 1159 862
rect 1174 852 1187 862
rect 1202 852 1232 866
rect 1275 852 1318 866
rect 1342 863 1349 870
rect 1352 866 1419 890
rect 1451 890 1623 892
rect 1421 868 1449 872
rect 1451 868 1531 890
rect 1552 888 1567 890
rect 1421 866 1531 868
rect 1352 862 1531 866
rect 1325 852 1355 862
rect 1357 852 1510 862
rect 1518 852 1548 862
rect 1552 852 1582 866
rect 1610 852 1623 890
rect 1695 896 1730 904
rect 1695 870 1696 896
rect 1703 870 1730 896
rect 1638 852 1668 866
rect 1695 862 1730 870
rect 1732 896 1773 904
rect 1732 870 1747 896
rect 1754 870 1773 896
rect 1837 892 1899 904
rect 1911 892 1986 904
rect 2044 892 2119 904
rect 2131 892 2162 904
rect 2168 892 2203 904
rect 1837 890 1999 892
rect 1732 862 1773 870
rect 1855 866 1868 890
rect 1883 888 1898 890
rect 1695 852 1696 862
rect 1711 852 1724 862
rect 1738 852 1739 862
rect 1754 852 1767 862
rect 1782 852 1812 866
rect 1855 852 1898 866
rect 1922 863 1929 870
rect 1932 866 1999 890
rect 2031 890 2203 892
rect 2001 868 2029 872
rect 2031 868 2111 890
rect 2132 888 2147 890
rect 2001 866 2111 868
rect 1932 862 2111 866
rect 1905 852 1935 862
rect 1937 852 2090 862
rect 2098 852 2128 862
rect 2132 852 2162 866
rect 2190 852 2203 890
rect 2275 896 2310 904
rect 2275 870 2276 896
rect 2283 870 2310 896
rect 2218 852 2248 866
rect 2275 862 2310 870
rect 2312 896 2353 904
rect 2312 870 2327 896
rect 2334 870 2353 896
rect 2417 892 2479 904
rect 2491 892 2566 904
rect 2624 892 2699 904
rect 2711 892 2742 904
rect 2748 892 2783 904
rect 2417 890 2579 892
rect 2312 862 2353 870
rect 2435 866 2448 890
rect 2463 888 2478 890
rect 2275 852 2276 862
rect 2291 852 2304 862
rect 2318 852 2319 862
rect 2334 852 2347 862
rect 2362 852 2392 866
rect 2435 852 2478 866
rect 2502 863 2509 870
rect 2512 866 2579 890
rect 2611 890 2783 892
rect 2581 868 2609 872
rect 2611 868 2691 890
rect 2712 888 2727 890
rect 2581 866 2691 868
rect 2512 862 2691 866
rect 2485 852 2515 862
rect 2517 852 2670 862
rect 2678 852 2708 862
rect 2712 852 2742 866
rect 2770 852 2783 890
rect 2855 896 2890 904
rect 2855 870 2856 896
rect 2863 870 2890 896
rect 2798 852 2828 866
rect 2855 862 2890 870
rect 2892 896 2933 904
rect 2892 870 2907 896
rect 2914 870 2933 896
rect 2997 892 3059 904
rect 3071 892 3146 904
rect 3204 892 3279 904
rect 3291 892 3322 904
rect 3328 892 3363 904
rect 2997 890 3159 892
rect 2892 862 2933 870
rect 3015 866 3028 890
rect 3043 888 3058 890
rect 2855 852 2856 862
rect 2871 852 2884 862
rect 2898 852 2899 862
rect 2914 852 2927 862
rect 2942 852 2972 866
rect 3015 852 3058 866
rect 3082 863 3089 870
rect 3092 866 3159 890
rect 3191 890 3363 892
rect 3161 868 3189 872
rect 3191 868 3271 890
rect 3292 888 3307 890
rect 3161 866 3271 868
rect 3092 862 3271 866
rect 3065 852 3095 862
rect 3097 852 3250 862
rect 3258 852 3288 862
rect 3292 852 3322 866
rect 3350 852 3363 890
rect 3435 896 3470 904
rect 3435 870 3436 896
rect 3443 870 3470 896
rect 3378 852 3408 866
rect 3435 862 3470 870
rect 3472 896 3513 904
rect 3472 870 3487 896
rect 3494 870 3513 896
rect 3577 892 3639 904
rect 3651 892 3726 904
rect 3784 892 3859 904
rect 3871 892 3902 904
rect 3908 892 3943 904
rect 3577 890 3739 892
rect 3472 862 3513 870
rect 3595 866 3608 890
rect 3623 888 3638 890
rect 3435 852 3436 862
rect 3451 852 3464 862
rect 3478 852 3479 862
rect 3494 852 3507 862
rect 3522 852 3552 866
rect 3595 852 3638 866
rect 3662 863 3669 870
rect 3672 866 3739 890
rect 3771 890 3943 892
rect 3741 868 3769 872
rect 3771 868 3851 890
rect 3872 888 3887 890
rect 3741 866 3851 868
rect 3672 862 3851 866
rect 3645 852 3675 862
rect 3677 852 3830 862
rect 3838 852 3868 862
rect 3872 852 3902 866
rect 3930 852 3943 890
rect 4015 896 4050 904
rect 4015 870 4016 896
rect 4023 870 4050 896
rect 3958 852 3988 866
rect 4015 862 4050 870
rect 4052 896 4093 904
rect 4052 870 4067 896
rect 4074 870 4093 896
rect 4157 892 4219 904
rect 4231 892 4306 904
rect 4364 892 4439 904
rect 4451 892 4482 904
rect 4488 892 4523 904
rect 4157 890 4319 892
rect 4052 862 4093 870
rect 4175 866 4188 890
rect 4203 888 4218 890
rect 4015 852 4016 862
rect 4031 852 4044 862
rect 4058 852 4059 862
rect 4074 852 4087 862
rect 4102 852 4132 866
rect 4175 852 4218 866
rect 4242 863 4249 870
rect 4252 866 4319 890
rect 4351 890 4523 892
rect 4321 868 4349 872
rect 4351 868 4431 890
rect 4452 888 4467 890
rect 4321 866 4431 868
rect 4252 862 4431 866
rect 4225 852 4255 862
rect 4257 852 4410 862
rect 4418 852 4448 862
rect 4452 852 4482 866
rect 4510 852 4523 890
rect 4595 896 4630 904
rect 4638 903 4639 919
rect 4654 903 4667 925
rect 4682 903 4712 925
rect 4755 921 4817 937
rect 4845 930 4856 946
rect 4861 941 4871 961
rect 4881 941 4895 961
rect 4898 948 4907 961
rect 4923 948 4932 961
rect 4861 930 4895 941
rect 4898 930 4907 946
rect 4923 930 4932 946
rect 4939 941 4949 961
rect 4959 941 4973 961
rect 4974 948 4985 961
rect 4939 930 4973 941
rect 4974 930 4985 946
rect 5031 937 5047 953
rect 5054 951 5084 1003
rect 5118 999 5119 1006
rect 5103 991 5119 999
rect 5090 959 5103 978
rect 5118 959 5148 975
rect 5090 943 5164 959
rect 5090 941 5103 943
rect 5118 941 5152 943
rect 4755 919 4768 921
rect 4783 919 4817 921
rect 4755 903 4817 919
rect 4861 914 4877 917
rect 4939 914 4969 925
rect 5017 921 5063 937
rect 5090 925 5164 941
rect 5017 919 5051 921
rect 5016 903 5063 919
rect 5090 903 5103 925
rect 5118 903 5148 925
rect 5175 903 5176 919
rect 5191 903 5204 1063
rect 5234 959 5247 1063
rect 5292 1041 5293 1051
rect 5313 1049 5321 1051
rect 5311 1047 5321 1049
rect 5308 1041 5321 1047
rect 5292 1037 5321 1041
rect 5326 1037 5356 1063
rect 5374 1049 5390 1051
rect 5462 1049 5513 1063
rect 5463 1047 5527 1049
rect 5570 1047 5585 1063
rect 5634 1060 5664 1063
rect 5634 1057 5670 1060
rect 5600 1049 5616 1051
rect 5374 1037 5389 1041
rect 5292 1035 5389 1037
rect 5417 1035 5585 1047
rect 5601 1037 5616 1041
rect 5634 1038 5673 1057
rect 5692 1051 5699 1052
rect 5698 1044 5699 1051
rect 5682 1041 5683 1044
rect 5698 1041 5711 1044
rect 5634 1037 5664 1038
rect 5673 1037 5679 1038
rect 5682 1037 5711 1041
rect 5601 1036 5711 1037
rect 5601 1035 5717 1036
rect 5276 1027 5327 1035
rect 5276 1015 5301 1027
rect 5308 1015 5327 1027
rect 5358 1027 5408 1035
rect 5358 1019 5374 1027
rect 5381 1025 5408 1027
rect 5417 1025 5638 1035
rect 5381 1015 5638 1025
rect 5667 1027 5717 1035
rect 5667 1018 5683 1027
rect 5276 1007 5327 1015
rect 5374 1007 5638 1015
rect 5664 1015 5683 1018
rect 5690 1015 5717 1027
rect 5664 1007 5717 1015
rect 5292 999 5293 1007
rect 5308 999 5321 1007
rect 5292 991 5308 999
rect 5289 984 5308 987
rect 5289 975 5311 984
rect 5262 965 5311 975
rect 5262 959 5292 965
rect 5311 960 5316 965
rect 5234 943 5308 959
rect 5326 951 5356 1007
rect 5391 997 5599 1007
rect 5634 1003 5679 1007
rect 5682 1006 5683 1007
rect 5698 1006 5711 1007
rect 5417 967 5606 997
rect 5432 964 5606 967
rect 5425 961 5606 964
rect 5234 941 5247 943
rect 5262 941 5296 943
rect 5234 925 5308 941
rect 5335 937 5348 951
rect 5363 937 5379 953
rect 5425 948 5436 961
rect 5218 903 5219 919
rect 5234 903 5247 925
rect 5262 903 5292 925
rect 5335 921 5397 937
rect 5425 930 5436 946
rect 5441 941 5451 961
rect 5461 941 5475 961
rect 5478 948 5487 961
rect 5503 948 5512 961
rect 5441 930 5475 941
rect 5478 930 5487 946
rect 5503 930 5512 946
rect 5519 941 5529 961
rect 5539 941 5553 961
rect 5554 948 5565 961
rect 5519 930 5553 941
rect 5554 930 5565 946
rect 5611 937 5627 953
rect 5634 951 5664 1003
rect 5698 999 5699 1006
rect 5683 991 5699 999
rect 5670 959 5683 978
rect 5698 959 5728 975
rect 5670 943 5744 959
rect 5670 941 5683 943
rect 5698 941 5732 943
rect 5335 919 5348 921
rect 5363 919 5397 921
rect 5335 903 5397 919
rect 5441 914 5457 917
rect 5519 914 5549 925
rect 5597 921 5643 937
rect 5670 925 5744 941
rect 5597 919 5631 921
rect 5596 903 5643 919
rect 5670 903 5683 925
rect 5698 903 5728 925
rect 5755 903 5756 919
rect 5771 903 5784 1063
rect 5814 959 5827 1063
rect 5872 1041 5873 1051
rect 5893 1049 5901 1051
rect 5891 1047 5901 1049
rect 5888 1041 5901 1047
rect 5872 1037 5901 1041
rect 5906 1037 5936 1063
rect 5954 1049 5970 1051
rect 6042 1049 6093 1063
rect 6043 1047 6107 1049
rect 6150 1047 6165 1063
rect 6214 1060 6244 1063
rect 6214 1057 6250 1060
rect 6180 1049 6196 1051
rect 5954 1037 5969 1041
rect 5872 1035 5969 1037
rect 5997 1035 6165 1047
rect 6181 1037 6196 1041
rect 6214 1038 6253 1057
rect 6272 1051 6279 1052
rect 6278 1044 6279 1051
rect 6262 1041 6263 1044
rect 6278 1041 6291 1044
rect 6214 1037 6244 1038
rect 6253 1037 6259 1038
rect 6262 1037 6291 1041
rect 6181 1036 6291 1037
rect 6181 1035 6297 1036
rect 5856 1027 5907 1035
rect 5856 1015 5881 1027
rect 5888 1015 5907 1027
rect 5938 1027 5988 1035
rect 5938 1019 5954 1027
rect 5961 1025 5988 1027
rect 5997 1025 6218 1035
rect 5961 1015 6218 1025
rect 6247 1027 6297 1035
rect 6247 1018 6263 1027
rect 5856 1007 5907 1015
rect 5954 1007 6218 1015
rect 6244 1015 6263 1018
rect 6270 1015 6297 1027
rect 6244 1007 6297 1015
rect 5872 999 5873 1007
rect 5888 999 5901 1007
rect 5872 991 5888 999
rect 5869 984 5888 987
rect 5869 975 5891 984
rect 5842 965 5891 975
rect 5842 959 5872 965
rect 5891 960 5896 965
rect 5814 943 5888 959
rect 5906 951 5936 1007
rect 5971 997 6179 1007
rect 6214 1003 6259 1007
rect 6262 1006 6263 1007
rect 6278 1006 6291 1007
rect 5997 967 6186 997
rect 6012 964 6186 967
rect 6005 961 6186 964
rect 5814 941 5827 943
rect 5842 941 5876 943
rect 5814 925 5888 941
rect 5915 937 5928 951
rect 5943 937 5959 953
rect 6005 948 6016 961
rect 5798 903 5799 919
rect 5814 903 5827 925
rect 5842 903 5872 925
rect 5915 921 5977 937
rect 6005 930 6016 946
rect 6021 941 6031 961
rect 6041 941 6055 961
rect 6058 948 6067 961
rect 6083 948 6092 961
rect 6021 930 6055 941
rect 6058 930 6067 946
rect 6083 930 6092 946
rect 6099 941 6109 961
rect 6119 941 6133 961
rect 6134 948 6145 961
rect 6099 930 6133 941
rect 6134 930 6145 946
rect 6191 937 6207 953
rect 6214 951 6244 1003
rect 6278 999 6279 1006
rect 6263 991 6279 999
rect 6250 959 6263 978
rect 6278 959 6308 975
rect 6250 943 6324 959
rect 6250 941 6263 943
rect 6278 941 6312 943
rect 5915 919 5928 921
rect 5943 919 5977 921
rect 5915 903 5977 919
rect 6021 914 6037 917
rect 6099 914 6129 925
rect 6177 921 6223 937
rect 6250 925 6324 941
rect 6177 919 6211 921
rect 6176 903 6223 919
rect 6250 903 6263 925
rect 6278 903 6308 925
rect 6335 903 6336 919
rect 6351 903 6364 1063
rect 6394 959 6407 1063
rect 6452 1041 6453 1051
rect 6473 1049 6481 1051
rect 6471 1047 6481 1049
rect 6468 1041 6481 1047
rect 6452 1037 6481 1041
rect 6486 1037 6516 1063
rect 6534 1049 6550 1051
rect 6622 1049 6673 1063
rect 6623 1047 6687 1049
rect 6730 1047 6745 1063
rect 6794 1060 6824 1063
rect 6794 1057 6830 1060
rect 6760 1049 6776 1051
rect 6534 1037 6549 1041
rect 6452 1035 6549 1037
rect 6577 1035 6745 1047
rect 6761 1037 6776 1041
rect 6794 1038 6833 1057
rect 6852 1051 6859 1052
rect 6858 1044 6859 1051
rect 6842 1041 6843 1044
rect 6858 1041 6871 1044
rect 6794 1037 6824 1038
rect 6833 1037 6839 1038
rect 6842 1037 6871 1041
rect 6761 1036 6871 1037
rect 6761 1035 6877 1036
rect 6436 1027 6487 1035
rect 6436 1015 6461 1027
rect 6468 1015 6487 1027
rect 6518 1027 6568 1035
rect 6518 1019 6534 1027
rect 6541 1025 6568 1027
rect 6577 1025 6798 1035
rect 6541 1015 6798 1025
rect 6827 1027 6877 1035
rect 6827 1018 6843 1027
rect 6436 1007 6487 1015
rect 6534 1007 6798 1015
rect 6824 1015 6843 1018
rect 6850 1015 6877 1027
rect 6824 1007 6877 1015
rect 6452 999 6453 1007
rect 6468 999 6481 1007
rect 6452 991 6468 999
rect 6449 984 6468 987
rect 6449 975 6471 984
rect 6422 965 6471 975
rect 6422 959 6452 965
rect 6471 960 6476 965
rect 6394 943 6468 959
rect 6486 951 6516 1007
rect 6551 997 6759 1007
rect 6794 1003 6839 1007
rect 6842 1006 6843 1007
rect 6858 1006 6871 1007
rect 6577 967 6766 997
rect 6592 964 6766 967
rect 6585 961 6766 964
rect 6394 941 6407 943
rect 6422 941 6456 943
rect 6394 925 6468 941
rect 6495 937 6508 951
rect 6523 937 6539 953
rect 6585 948 6596 961
rect 6378 903 6379 919
rect 6394 903 6407 925
rect 6422 903 6452 925
rect 6495 921 6557 937
rect 6585 930 6596 946
rect 6601 941 6611 961
rect 6621 941 6635 961
rect 6638 948 6647 961
rect 6663 948 6672 961
rect 6601 930 6635 941
rect 6638 930 6647 946
rect 6663 930 6672 946
rect 6679 941 6689 961
rect 6699 941 6713 961
rect 6714 948 6725 961
rect 6679 930 6713 941
rect 6714 930 6725 946
rect 6771 937 6787 953
rect 6794 951 6824 1003
rect 6858 999 6859 1006
rect 6843 991 6859 999
rect 6830 959 6843 978
rect 6858 959 6888 975
rect 6830 943 6904 959
rect 6830 941 6843 943
rect 6858 941 6892 943
rect 6495 919 6508 921
rect 6523 919 6557 921
rect 6495 903 6557 919
rect 6601 914 6617 917
rect 6679 914 6709 925
rect 6757 921 6803 937
rect 6830 925 6904 941
rect 6757 919 6791 921
rect 6756 903 6803 919
rect 6830 903 6843 925
rect 6858 903 6888 925
rect 6915 903 6916 919
rect 6931 903 6944 1063
rect 4595 870 4596 896
rect 4603 870 4630 896
rect 4538 852 4568 866
rect 4595 862 4630 870
rect 4632 895 4673 903
rect 4632 869 4647 895
rect 4654 869 4673 895
rect 4737 891 4799 903
rect 4811 891 4886 903
rect 4944 891 5019 903
rect 5031 891 5062 903
rect 5068 891 5103 903
rect 4737 889 4899 891
rect 4595 852 4596 862
rect 4611 852 4624 862
rect 4632 861 4673 869
rect 4755 865 4768 889
rect 4783 887 4798 889
rect 4832 871 4899 889
rect 4931 889 5103 891
rect 4931 871 5011 889
rect 5032 887 5047 889
rect -2 851 4624 852
rect 4638 851 4639 861
rect 4654 851 4667 861
rect 4682 851 4712 865
rect 4755 851 4798 865
rect 4822 862 4829 869
rect 4832 861 5011 871
rect 4805 851 4835 861
rect 4837 851 4990 861
rect 4998 851 5028 861
rect 5032 851 5062 865
rect 5090 851 5103 889
rect 5175 895 5210 903
rect 5175 869 5176 895
rect 5183 869 5210 895
rect 5118 851 5148 865
rect 5175 861 5210 869
rect 5212 895 5253 903
rect 5212 869 5227 895
rect 5234 869 5253 895
rect 5317 891 5379 903
rect 5391 891 5466 903
rect 5524 891 5599 903
rect 5611 891 5642 903
rect 5648 891 5683 903
rect 5317 889 5479 891
rect 5212 861 5253 869
rect 5335 865 5348 889
rect 5363 887 5378 889
rect 5412 871 5479 889
rect 5511 889 5683 891
rect 5511 871 5591 889
rect 5612 887 5627 889
rect 5175 851 5176 861
rect 5191 851 5204 861
rect 5218 851 5219 861
rect 5234 851 5247 861
rect 5262 851 5292 865
rect 5335 851 5378 865
rect 5402 862 5409 869
rect 5412 861 5591 871
rect 5385 851 5415 861
rect 5417 851 5570 861
rect 5578 851 5608 861
rect 5612 851 5642 865
rect 5670 851 5683 889
rect 5755 895 5790 903
rect 5755 869 5756 895
rect 5763 869 5790 895
rect 5698 851 5728 865
rect 5755 861 5790 869
rect 5792 895 5833 903
rect 5792 869 5807 895
rect 5814 869 5833 895
rect 5897 891 5959 903
rect 5971 891 6046 903
rect 6104 891 6179 903
rect 6191 891 6222 903
rect 6228 891 6263 903
rect 5897 889 6059 891
rect 5792 861 5833 869
rect 5915 865 5928 889
rect 5943 887 5958 889
rect 5992 871 6059 889
rect 6091 889 6263 891
rect 6091 871 6171 889
rect 6192 887 6207 889
rect 5755 851 5756 861
rect 5771 851 5784 861
rect 5798 851 5799 861
rect 5814 851 5827 861
rect 5842 851 5872 865
rect 5915 851 5958 865
rect 5982 862 5989 869
rect 5992 861 6171 871
rect 5965 851 5995 861
rect 5997 851 6150 861
rect 6158 851 6188 861
rect 6192 851 6222 865
rect 6250 851 6263 889
rect 6335 895 6370 903
rect 6335 869 6336 895
rect 6343 869 6370 895
rect 6278 851 6308 865
rect 6335 861 6370 869
rect 6372 895 6413 903
rect 6372 869 6387 895
rect 6394 869 6413 895
rect 6477 891 6539 903
rect 6551 891 6626 903
rect 6684 891 6759 903
rect 6771 891 6802 903
rect 6808 891 6843 903
rect 6477 889 6639 891
rect 6372 861 6413 869
rect 6495 865 6508 889
rect 6523 887 6538 889
rect 6572 871 6639 889
rect 6671 889 6843 891
rect 6671 871 6751 889
rect 6772 887 6787 889
rect 6335 851 6336 861
rect 6351 851 6364 861
rect 6378 851 6379 861
rect 6394 851 6407 861
rect 6422 851 6452 865
rect 6495 851 6538 865
rect 6562 862 6569 869
rect 6572 861 6751 871
rect 6545 851 6575 861
rect 6577 851 6730 861
rect 6738 851 6768 861
rect 6772 851 6802 865
rect 6830 851 6843 889
rect 6915 895 6950 903
rect 6915 869 6916 895
rect 6923 869 6950 895
rect 6858 851 6888 865
rect 6915 861 6950 869
rect 6915 851 6916 861
rect 6931 851 6944 861
rect -2 846 6944 851
rect -1 838 6944 846
rect 14 808 27 838
rect 42 820 72 838
rect 115 824 129 838
rect 165 824 385 838
rect 116 822 129 824
rect 82 810 97 822
rect 79 808 101 810
rect 106 808 136 822
rect 197 820 350 824
rect 179 808 371 820
rect 414 808 444 822
rect 450 808 463 838
rect 478 820 508 838
rect 551 808 564 838
rect 594 808 607 838
rect 622 820 652 838
rect 695 824 709 838
rect 745 824 965 838
rect 696 822 709 824
rect 662 810 677 822
rect 659 808 681 810
rect 686 808 716 822
rect 777 820 930 824
rect 759 808 951 820
rect 994 808 1024 822
rect 1030 808 1043 838
rect 1058 820 1088 838
rect 1131 808 1144 838
rect 1174 808 1187 838
rect 1202 820 1232 838
rect 1275 824 1289 838
rect 1325 824 1545 838
rect 1276 822 1289 824
rect 1242 810 1257 822
rect 1239 808 1261 810
rect 1266 808 1296 822
rect 1357 820 1510 824
rect 1339 808 1531 820
rect 1574 808 1604 822
rect 1610 808 1623 838
rect 1638 820 1668 838
rect 1711 808 1724 838
rect 1754 808 1767 838
rect 1782 820 1812 838
rect 1855 824 1869 838
rect 1905 824 2125 838
rect 1856 822 1869 824
rect 1822 810 1837 822
rect 1819 808 1841 810
rect 1846 808 1876 822
rect 1937 820 2090 824
rect 1919 808 2111 820
rect 2154 808 2184 822
rect 2190 808 2203 838
rect 2218 820 2248 838
rect 2291 808 2304 838
rect 2334 808 2347 838
rect 2362 820 2392 838
rect 2435 824 2449 838
rect 2485 824 2705 838
rect 2436 822 2449 824
rect 2402 810 2417 822
rect 2399 808 2421 810
rect 2426 808 2456 822
rect 2517 820 2670 824
rect 2499 808 2691 820
rect 2734 808 2764 822
rect 2770 808 2783 838
rect 2798 820 2828 838
rect 2871 808 2884 838
rect 2914 808 2927 838
rect 2942 820 2972 838
rect 3015 824 3029 838
rect 3065 824 3285 838
rect 3016 822 3029 824
rect 2982 810 2997 822
rect 2979 808 3001 810
rect 3006 808 3036 822
rect 3097 820 3250 824
rect 3079 808 3271 820
rect 3314 808 3344 822
rect 3350 808 3363 838
rect 3378 820 3408 838
rect 3451 808 3464 838
rect 3494 808 3507 838
rect 3522 820 3552 838
rect 3595 824 3609 838
rect 3645 824 3865 838
rect 3596 822 3609 824
rect 3562 810 3577 822
rect 3559 808 3581 810
rect 3586 808 3616 822
rect 3677 820 3830 824
rect 3659 808 3851 820
rect 3894 808 3924 822
rect 3930 808 3943 838
rect 3958 820 3988 838
rect 4031 808 4044 838
rect 4074 808 4087 838
rect 4102 820 4132 838
rect 4175 824 4189 838
rect 4225 824 4445 838
rect 4176 822 4189 824
rect 4142 810 4157 822
rect 4139 808 4161 810
rect 4166 808 4196 822
rect 4257 820 4410 824
rect 4239 808 4431 820
rect 4474 808 4504 822
rect 4510 808 4523 838
rect 4538 820 4568 838
rect 4611 837 6944 838
rect 4611 808 4624 837
rect -1 807 4624 808
rect 4654 807 4667 837
rect 4682 819 4712 837
rect 4755 823 4769 837
rect 4805 823 5025 837
rect 4756 821 4769 823
rect 4722 809 4737 821
rect 4719 807 4741 809
rect 4746 807 4776 821
rect 4837 819 4990 823
rect 4819 807 5011 819
rect 5054 807 5084 821
rect 5090 807 5103 837
rect 5118 819 5148 837
rect 5191 807 5204 837
rect 5234 807 5247 837
rect 5262 819 5292 837
rect 5335 823 5349 837
rect 5385 823 5605 837
rect 5336 821 5349 823
rect 5302 809 5317 821
rect 5299 807 5321 809
rect 5326 807 5356 821
rect 5417 819 5570 823
rect 5399 807 5591 819
rect 5634 807 5664 821
rect 5670 807 5683 837
rect 5698 819 5728 837
rect 5771 807 5784 837
rect 5814 807 5827 837
rect 5842 819 5872 837
rect 5915 823 5929 837
rect 5965 823 6185 837
rect 5916 821 5929 823
rect 5882 809 5897 821
rect 5879 807 5901 809
rect 5906 807 5936 821
rect 5997 819 6150 823
rect 5979 807 6171 819
rect 6214 807 6244 821
rect 6250 807 6263 837
rect 6278 819 6308 837
rect 6351 807 6364 837
rect 6394 807 6407 837
rect 6422 819 6452 837
rect 6495 823 6509 837
rect 6545 823 6765 837
rect 6496 821 6509 823
rect 6462 809 6477 821
rect 6459 807 6481 809
rect 6486 807 6516 821
rect 6577 819 6730 823
rect 6559 807 6751 819
rect 6794 807 6824 821
rect 6830 807 6843 837
rect 6858 819 6888 837
rect 6931 807 6944 837
rect -1 794 6944 807
rect 14 690 27 794
rect 72 772 73 782
rect 88 772 101 782
rect 72 768 101 772
rect 106 768 136 794
rect 154 780 170 782
rect 242 780 295 794
rect 243 778 307 780
rect 350 778 365 794
rect 414 791 444 794
rect 414 788 450 791
rect 380 780 396 782
rect 154 768 169 772
rect 72 766 169 768
rect 197 766 365 778
rect 381 768 396 772
rect 414 769 453 788
rect 472 782 479 783
rect 478 775 479 782
rect 462 772 463 775
rect 478 772 491 775
rect 414 768 444 769
rect 453 768 459 769
rect 462 768 491 772
rect 381 767 491 768
rect 381 766 497 767
rect 56 758 107 766
rect 56 746 81 758
rect 88 746 107 758
rect 138 758 188 766
rect 138 750 154 758
rect 161 756 188 758
rect 197 756 418 766
rect 161 746 418 756
rect 447 758 497 766
rect 447 749 463 758
rect 56 738 107 746
rect 154 738 418 746
rect 444 746 463 749
rect 470 746 497 758
rect 444 738 497 746
rect 72 730 73 738
rect 88 730 101 738
rect 72 722 88 730
rect 69 715 88 718
rect 69 706 91 715
rect 42 696 91 706
rect 42 690 72 696
rect 91 691 96 696
rect 14 674 88 690
rect 106 682 136 738
rect 171 728 379 738
rect 414 734 459 738
rect 462 737 463 738
rect 478 737 491 738
rect 197 698 386 728
rect 212 695 386 698
rect 205 692 386 695
rect 14 672 27 674
rect 42 672 76 674
rect 14 656 88 672
rect 115 668 128 682
rect 143 668 159 684
rect 205 679 216 692
rect -2 634 -1 650
rect 14 634 27 656
rect 42 634 72 656
rect 115 652 177 668
rect 205 661 216 677
rect 221 672 231 692
rect 241 672 255 692
rect 258 679 267 692
rect 283 679 292 692
rect 221 661 255 672
rect 258 661 267 677
rect 283 661 292 677
rect 299 672 309 692
rect 319 672 333 692
rect 334 679 345 692
rect 299 661 333 672
rect 334 661 345 677
rect 391 668 407 684
rect 414 682 444 734
rect 478 730 479 737
rect 463 722 479 730
rect 450 690 463 709
rect 478 690 508 706
rect 450 674 524 690
rect 450 672 463 674
rect 478 672 512 674
rect 115 650 128 652
rect 143 650 177 652
rect 115 634 177 650
rect 221 645 237 648
rect 299 645 329 656
rect 377 652 423 668
rect 450 656 524 672
rect 377 650 411 652
rect 376 634 423 650
rect 450 634 463 656
rect 478 634 508 656
rect 535 634 536 650
rect 551 634 564 794
rect 594 690 607 794
rect 652 772 653 782
rect 668 772 681 782
rect 652 768 681 772
rect 686 768 716 794
rect 734 780 750 782
rect 822 780 875 794
rect 823 778 887 780
rect 930 778 945 794
rect 994 791 1024 794
rect 994 788 1030 791
rect 960 780 976 782
rect 734 768 749 772
rect 652 766 749 768
rect 777 766 945 778
rect 961 768 976 772
rect 994 769 1033 788
rect 1052 782 1059 783
rect 1058 775 1059 782
rect 1042 772 1043 775
rect 1058 772 1071 775
rect 994 768 1024 769
rect 1033 768 1039 769
rect 1042 768 1071 772
rect 961 767 1071 768
rect 961 766 1077 767
rect 636 758 687 766
rect 636 746 661 758
rect 668 746 687 758
rect 718 758 768 766
rect 718 750 734 758
rect 741 756 768 758
rect 777 756 998 766
rect 741 746 998 756
rect 1027 758 1077 766
rect 1027 749 1043 758
rect 636 738 687 746
rect 734 738 998 746
rect 1024 746 1043 749
rect 1050 746 1077 758
rect 1024 738 1077 746
rect 652 730 653 738
rect 668 730 681 738
rect 652 722 668 730
rect 649 715 668 718
rect 649 706 671 715
rect 622 696 671 706
rect 622 690 652 696
rect 671 691 676 696
rect 594 674 668 690
rect 686 682 716 738
rect 751 728 959 738
rect 994 734 1039 738
rect 1042 737 1043 738
rect 1058 737 1071 738
rect 777 698 966 728
rect 792 695 966 698
rect 785 692 966 695
rect 594 672 607 674
rect 622 672 656 674
rect 594 656 668 672
rect 695 668 708 682
rect 723 668 739 684
rect 785 679 796 692
rect 578 634 579 650
rect 594 634 607 656
rect 622 634 652 656
rect 695 652 757 668
rect 785 661 796 677
rect 801 672 811 692
rect 821 672 835 692
rect 838 679 847 692
rect 863 679 872 692
rect 801 661 835 672
rect 838 661 847 677
rect 863 661 872 677
rect 879 672 889 692
rect 899 672 913 692
rect 914 679 925 692
rect 879 661 913 672
rect 914 661 925 677
rect 971 668 987 684
rect 994 682 1024 734
rect 1058 730 1059 737
rect 1043 722 1059 730
rect 1030 690 1043 709
rect 1058 690 1088 706
rect 1030 674 1104 690
rect 1030 672 1043 674
rect 1058 672 1092 674
rect 695 650 708 652
rect 723 650 757 652
rect 695 634 757 650
rect 801 645 817 648
rect 879 645 909 656
rect 957 652 1003 668
rect 1030 656 1104 672
rect 957 650 991 652
rect 956 634 1003 650
rect 1030 634 1043 656
rect 1058 634 1088 656
rect 1115 634 1116 650
rect 1131 634 1144 794
rect 1174 690 1187 794
rect 1232 772 1233 782
rect 1248 772 1261 782
rect 1232 768 1261 772
rect 1266 768 1296 794
rect 1314 780 1330 782
rect 1402 780 1455 794
rect 1403 778 1467 780
rect 1510 778 1525 794
rect 1574 791 1604 794
rect 1574 788 1610 791
rect 1540 780 1556 782
rect 1314 768 1329 772
rect 1232 766 1329 768
rect 1357 766 1525 778
rect 1541 768 1556 772
rect 1574 769 1613 788
rect 1632 782 1639 783
rect 1638 775 1639 782
rect 1622 772 1623 775
rect 1638 772 1651 775
rect 1574 768 1604 769
rect 1613 768 1619 769
rect 1622 768 1651 772
rect 1541 767 1651 768
rect 1541 766 1657 767
rect 1216 758 1267 766
rect 1216 746 1241 758
rect 1248 746 1267 758
rect 1298 758 1348 766
rect 1298 750 1314 758
rect 1321 756 1348 758
rect 1357 756 1578 766
rect 1321 746 1578 756
rect 1607 758 1657 766
rect 1607 749 1623 758
rect 1216 738 1267 746
rect 1314 738 1578 746
rect 1604 746 1623 749
rect 1630 746 1657 758
rect 1604 738 1657 746
rect 1232 730 1233 738
rect 1248 730 1261 738
rect 1232 722 1248 730
rect 1229 715 1248 718
rect 1229 706 1251 715
rect 1202 696 1251 706
rect 1202 690 1232 696
rect 1251 691 1256 696
rect 1174 674 1248 690
rect 1266 682 1296 738
rect 1331 728 1539 738
rect 1574 734 1619 738
rect 1622 737 1623 738
rect 1638 737 1651 738
rect 1357 698 1546 728
rect 1372 695 1546 698
rect 1365 692 1546 695
rect 1174 672 1187 674
rect 1202 672 1236 674
rect 1174 656 1248 672
rect 1275 668 1288 682
rect 1303 668 1319 684
rect 1365 679 1376 692
rect 1158 634 1159 650
rect 1174 634 1187 656
rect 1202 634 1232 656
rect 1275 652 1337 668
rect 1365 661 1376 677
rect 1381 672 1391 692
rect 1401 672 1415 692
rect 1418 679 1427 692
rect 1443 679 1452 692
rect 1381 661 1415 672
rect 1418 661 1427 677
rect 1443 661 1452 677
rect 1459 672 1469 692
rect 1479 672 1493 692
rect 1494 679 1505 692
rect 1459 661 1493 672
rect 1494 661 1505 677
rect 1551 668 1567 684
rect 1574 682 1604 734
rect 1638 730 1639 737
rect 1623 722 1639 730
rect 1610 690 1623 709
rect 1638 690 1668 706
rect 1610 674 1684 690
rect 1610 672 1623 674
rect 1638 672 1672 674
rect 1275 650 1288 652
rect 1303 650 1337 652
rect 1275 634 1337 650
rect 1381 645 1397 648
rect 1459 645 1489 656
rect 1537 652 1583 668
rect 1610 656 1684 672
rect 1537 650 1571 652
rect 1536 634 1583 650
rect 1610 634 1623 656
rect 1638 634 1668 656
rect 1695 634 1696 650
rect 1711 634 1724 794
rect 1754 690 1767 794
rect 1812 772 1813 782
rect 1828 772 1841 782
rect 1812 768 1841 772
rect 1846 768 1876 794
rect 1894 780 1910 782
rect 1982 780 2035 794
rect 1983 778 2047 780
rect 2090 778 2105 794
rect 2154 791 2184 794
rect 2154 788 2190 791
rect 2120 780 2136 782
rect 1894 768 1909 772
rect 1812 766 1909 768
rect 1937 766 2105 778
rect 2121 768 2136 772
rect 2154 769 2193 788
rect 2212 782 2219 783
rect 2218 775 2219 782
rect 2202 772 2203 775
rect 2218 772 2231 775
rect 2154 768 2184 769
rect 2193 768 2199 769
rect 2202 768 2231 772
rect 2121 767 2231 768
rect 2121 766 2237 767
rect 1796 758 1847 766
rect 1796 746 1821 758
rect 1828 746 1847 758
rect 1878 758 1928 766
rect 1878 750 1894 758
rect 1901 756 1928 758
rect 1937 756 2158 766
rect 1901 746 2158 756
rect 2187 758 2237 766
rect 2187 749 2203 758
rect 1796 738 1847 746
rect 1894 738 2158 746
rect 2184 746 2203 749
rect 2210 746 2237 758
rect 2184 738 2237 746
rect 1812 730 1813 738
rect 1828 730 1841 738
rect 1812 722 1828 730
rect 1809 715 1828 718
rect 1809 706 1831 715
rect 1782 696 1831 706
rect 1782 690 1812 696
rect 1831 691 1836 696
rect 1754 674 1828 690
rect 1846 682 1876 738
rect 1911 728 2119 738
rect 2154 734 2199 738
rect 2202 737 2203 738
rect 2218 737 2231 738
rect 1937 698 2126 728
rect 1952 695 2126 698
rect 1945 692 2126 695
rect 1754 672 1767 674
rect 1782 672 1816 674
rect 1754 656 1828 672
rect 1855 668 1868 682
rect 1883 668 1899 684
rect 1945 679 1956 692
rect 1738 634 1739 650
rect 1754 634 1767 656
rect 1782 634 1812 656
rect 1855 652 1917 668
rect 1945 661 1956 677
rect 1961 672 1971 692
rect 1981 672 1995 692
rect 1998 679 2007 692
rect 2023 679 2032 692
rect 1961 661 1995 672
rect 1998 661 2007 677
rect 2023 661 2032 677
rect 2039 672 2049 692
rect 2059 672 2073 692
rect 2074 679 2085 692
rect 2039 661 2073 672
rect 2074 661 2085 677
rect 2131 668 2147 684
rect 2154 682 2184 734
rect 2218 730 2219 737
rect 2203 722 2219 730
rect 2190 690 2203 709
rect 2218 690 2248 706
rect 2190 674 2264 690
rect 2190 672 2203 674
rect 2218 672 2252 674
rect 1855 650 1868 652
rect 1883 650 1917 652
rect 1855 634 1917 650
rect 1961 645 1977 648
rect 2039 645 2069 656
rect 2117 652 2163 668
rect 2190 656 2264 672
rect 2117 650 2151 652
rect 2116 634 2163 650
rect 2190 634 2203 656
rect 2218 634 2248 656
rect 2275 634 2276 650
rect 2291 634 2304 794
rect 2334 690 2347 794
rect 2392 772 2393 782
rect 2408 772 2421 782
rect 2392 768 2421 772
rect 2426 768 2456 794
rect 2474 780 2490 782
rect 2562 780 2615 794
rect 2563 778 2627 780
rect 2670 778 2685 794
rect 2734 791 2764 794
rect 2734 788 2770 791
rect 2700 780 2716 782
rect 2474 768 2489 772
rect 2392 766 2489 768
rect 2517 766 2685 778
rect 2701 768 2716 772
rect 2734 769 2773 788
rect 2792 782 2799 783
rect 2798 775 2799 782
rect 2782 772 2783 775
rect 2798 772 2811 775
rect 2734 768 2764 769
rect 2773 768 2779 769
rect 2782 768 2811 772
rect 2701 767 2811 768
rect 2701 766 2817 767
rect 2376 758 2427 766
rect 2376 746 2401 758
rect 2408 746 2427 758
rect 2458 758 2508 766
rect 2458 750 2474 758
rect 2481 756 2508 758
rect 2517 756 2738 766
rect 2481 746 2738 756
rect 2767 758 2817 766
rect 2767 749 2783 758
rect 2376 738 2427 746
rect 2474 738 2738 746
rect 2764 746 2783 749
rect 2790 746 2817 758
rect 2764 738 2817 746
rect 2392 730 2393 738
rect 2408 730 2421 738
rect 2392 722 2408 730
rect 2389 715 2408 718
rect 2389 706 2411 715
rect 2362 696 2411 706
rect 2362 690 2392 696
rect 2411 691 2416 696
rect 2334 674 2408 690
rect 2426 682 2456 738
rect 2491 728 2699 738
rect 2734 734 2779 738
rect 2782 737 2783 738
rect 2798 737 2811 738
rect 2517 698 2706 728
rect 2532 695 2706 698
rect 2525 692 2706 695
rect 2334 672 2347 674
rect 2362 672 2396 674
rect 2334 656 2408 672
rect 2435 668 2448 682
rect 2463 668 2479 684
rect 2525 679 2536 692
rect 2318 634 2319 650
rect 2334 634 2347 656
rect 2362 634 2392 656
rect 2435 652 2497 668
rect 2525 661 2536 677
rect 2541 672 2551 692
rect 2561 672 2575 692
rect 2578 679 2587 692
rect 2603 679 2612 692
rect 2541 661 2575 672
rect 2578 661 2587 677
rect 2603 661 2612 677
rect 2619 672 2629 692
rect 2639 672 2653 692
rect 2654 679 2665 692
rect 2619 661 2653 672
rect 2654 661 2665 677
rect 2711 668 2727 684
rect 2734 682 2764 734
rect 2798 730 2799 737
rect 2783 722 2799 730
rect 2770 690 2783 709
rect 2798 690 2828 706
rect 2770 674 2844 690
rect 2770 672 2783 674
rect 2798 672 2832 674
rect 2435 650 2448 652
rect 2463 650 2497 652
rect 2435 634 2497 650
rect 2541 645 2557 648
rect 2619 645 2649 656
rect 2697 652 2743 668
rect 2770 656 2844 672
rect 2697 650 2731 652
rect 2696 634 2743 650
rect 2770 634 2783 656
rect 2798 634 2828 656
rect 2855 634 2856 650
rect 2871 634 2884 794
rect 2914 690 2927 794
rect 2972 772 2973 782
rect 2988 772 3001 782
rect 2972 768 3001 772
rect 3006 768 3036 794
rect 3054 780 3070 782
rect 3142 780 3195 794
rect 3143 778 3205 780
rect 3250 778 3265 794
rect 3314 791 3344 794
rect 3314 788 3350 791
rect 3280 780 3296 782
rect 3054 768 3069 772
rect 2972 766 3069 768
rect 3097 766 3265 778
rect 3281 768 3296 772
rect 3314 769 3353 788
rect 3372 782 3379 783
rect 3378 775 3379 782
rect 3362 772 3363 775
rect 3378 772 3391 775
rect 3314 768 3344 769
rect 3353 768 3359 769
rect 3362 768 3391 772
rect 3281 767 3391 768
rect 3281 766 3397 767
rect 2956 758 3007 766
rect 2956 746 2981 758
rect 2988 746 3007 758
rect 3038 758 3088 766
rect 3038 750 3054 758
rect 3061 756 3088 758
rect 3097 756 3318 766
rect 3061 746 3318 756
rect 3347 758 3397 766
rect 3347 749 3363 758
rect 2956 738 3007 746
rect 3054 738 3318 746
rect 3344 746 3363 749
rect 3370 746 3397 758
rect 3344 738 3397 746
rect 2972 730 2973 738
rect 2988 730 3001 738
rect 2972 722 2988 730
rect 2969 715 2988 718
rect 2969 706 2991 715
rect 2942 696 2991 706
rect 2942 690 2972 696
rect 2991 691 2996 696
rect 2914 674 2988 690
rect 3006 682 3036 738
rect 3071 728 3279 738
rect 3314 734 3359 738
rect 3362 737 3363 738
rect 3378 737 3391 738
rect 3097 698 3286 728
rect 3112 695 3286 698
rect 3105 692 3286 695
rect 2914 672 2927 674
rect 2942 672 2976 674
rect 2914 656 2988 672
rect 3015 668 3028 682
rect 3043 668 3059 684
rect 3105 679 3116 692
rect 2898 634 2899 650
rect 2914 634 2927 656
rect 2942 634 2972 656
rect 3015 652 3077 668
rect 3105 661 3116 677
rect 3121 672 3131 692
rect 3141 672 3155 692
rect 3158 679 3167 692
rect 3183 679 3192 692
rect 3121 661 3155 672
rect 3158 661 3167 677
rect 3183 661 3192 677
rect 3199 672 3209 692
rect 3219 672 3233 692
rect 3234 679 3245 692
rect 3199 661 3233 672
rect 3234 661 3245 677
rect 3291 668 3307 684
rect 3314 682 3344 734
rect 3378 730 3379 737
rect 3363 722 3379 730
rect 3350 690 3363 709
rect 3378 690 3408 706
rect 3350 674 3424 690
rect 3350 672 3363 674
rect 3378 672 3412 674
rect 3015 650 3028 652
rect 3043 650 3077 652
rect 3015 634 3077 650
rect 3121 645 3137 648
rect 3199 645 3229 656
rect 3277 652 3323 668
rect 3350 656 3424 672
rect 3277 650 3311 652
rect 3276 634 3323 650
rect 3350 634 3363 656
rect 3378 634 3408 656
rect 3435 634 3436 650
rect 3451 634 3464 794
rect 3494 690 3507 794
rect 3552 772 3553 782
rect 3568 772 3581 782
rect 3552 768 3581 772
rect 3586 768 3616 794
rect 3634 780 3650 782
rect 3722 780 3775 794
rect 3723 778 3787 780
rect 3830 778 3845 794
rect 3894 791 3924 794
rect 3894 788 3930 791
rect 3860 780 3876 782
rect 3634 768 3649 772
rect 3552 766 3649 768
rect 3677 766 3845 778
rect 3861 768 3876 772
rect 3894 769 3933 788
rect 3952 782 3959 783
rect 3958 775 3959 782
rect 3942 772 3943 775
rect 3958 772 3971 775
rect 3894 768 3924 769
rect 3933 768 3939 769
rect 3942 768 3971 772
rect 3861 767 3971 768
rect 3861 766 3977 767
rect 3536 758 3587 766
rect 3536 746 3561 758
rect 3568 746 3587 758
rect 3618 758 3668 766
rect 3618 750 3634 758
rect 3641 756 3668 758
rect 3677 756 3898 766
rect 3641 746 3898 756
rect 3927 758 3977 766
rect 3927 749 3943 758
rect 3536 738 3587 746
rect 3634 738 3898 746
rect 3924 746 3943 749
rect 3950 746 3977 758
rect 3924 738 3977 746
rect 3552 730 3553 738
rect 3568 730 3581 738
rect 3552 722 3568 730
rect 3549 715 3568 718
rect 3549 706 3571 715
rect 3522 696 3571 706
rect 3522 690 3552 696
rect 3571 691 3576 696
rect 3494 674 3568 690
rect 3586 682 3616 738
rect 3651 728 3859 738
rect 3894 734 3939 738
rect 3942 737 3943 738
rect 3958 737 3971 738
rect 3677 698 3866 728
rect 3692 695 3866 698
rect 3685 692 3866 695
rect 3494 672 3507 674
rect 3522 672 3556 674
rect 3494 656 3568 672
rect 3595 668 3608 682
rect 3623 668 3639 684
rect 3685 679 3696 692
rect 3478 634 3479 650
rect 3494 634 3507 656
rect 3522 634 3552 656
rect 3595 652 3657 668
rect 3685 661 3696 677
rect 3701 672 3711 692
rect 3721 672 3735 692
rect 3738 679 3747 692
rect 3763 679 3772 692
rect 3701 661 3735 672
rect 3738 661 3747 677
rect 3763 661 3772 677
rect 3779 672 3789 692
rect 3799 672 3813 692
rect 3814 679 3825 692
rect 3779 661 3813 672
rect 3814 661 3825 677
rect 3871 668 3887 684
rect 3894 682 3924 734
rect 3958 730 3959 737
rect 3943 722 3959 730
rect 3930 690 3943 709
rect 3958 690 3988 706
rect 3930 674 4004 690
rect 3930 672 3943 674
rect 3958 672 3992 674
rect 3595 650 3608 652
rect 3623 650 3657 652
rect 3595 634 3657 650
rect 3701 645 3717 648
rect 3779 645 3809 656
rect 3857 652 3903 668
rect 3930 656 4004 672
rect 3857 650 3891 652
rect 3856 634 3903 650
rect 3930 634 3943 656
rect 3958 634 3988 656
rect 4015 634 4016 650
rect 4031 634 4044 794
rect 4074 690 4087 794
rect 4132 772 4133 782
rect 4148 772 4161 782
rect 4132 768 4161 772
rect 4166 768 4196 794
rect 4214 780 4230 782
rect 4302 780 4355 794
rect 4303 778 4367 780
rect 4410 778 4425 794
rect 4474 791 4504 794
rect 4611 793 6944 794
rect 4474 788 4510 791
rect 4440 780 4456 782
rect 4214 768 4229 772
rect 4132 766 4229 768
rect 4257 766 4425 778
rect 4441 768 4456 772
rect 4474 769 4513 788
rect 4532 782 4539 783
rect 4538 775 4539 782
rect 4522 772 4523 775
rect 4538 772 4551 775
rect 4474 768 4504 769
rect 4513 768 4519 769
rect 4522 768 4551 772
rect 4441 767 4551 768
rect 4441 766 4557 767
rect 4116 758 4167 766
rect 4116 746 4141 758
rect 4148 746 4167 758
rect 4198 758 4248 766
rect 4198 750 4214 758
rect 4221 756 4248 758
rect 4257 756 4478 766
rect 4221 746 4478 756
rect 4507 758 4557 766
rect 4507 749 4523 758
rect 4116 738 4167 746
rect 4214 738 4478 746
rect 4504 746 4523 749
rect 4530 746 4557 758
rect 4504 738 4557 746
rect 4132 730 4133 738
rect 4148 730 4161 738
rect 4132 722 4148 730
rect 4129 715 4148 718
rect 4129 706 4151 715
rect 4102 696 4151 706
rect 4102 690 4132 696
rect 4151 691 4156 696
rect 4074 674 4148 690
rect 4166 682 4196 738
rect 4231 728 4439 738
rect 4474 734 4519 738
rect 4522 737 4523 738
rect 4538 737 4551 738
rect 4257 698 4446 728
rect 4272 695 4446 698
rect 4265 692 4446 695
rect 4074 672 4087 674
rect 4102 672 4136 674
rect 4074 656 4148 672
rect 4175 668 4188 682
rect 4203 668 4219 684
rect 4265 679 4276 692
rect 4058 634 4059 650
rect 4074 634 4087 656
rect 4102 634 4132 656
rect 4175 652 4237 668
rect 4265 661 4276 677
rect 4281 672 4291 692
rect 4301 672 4315 692
rect 4318 679 4327 692
rect 4343 679 4352 692
rect 4281 661 4315 672
rect 4318 661 4327 677
rect 4343 661 4352 677
rect 4359 672 4369 692
rect 4379 672 4393 692
rect 4394 679 4405 692
rect 4359 661 4393 672
rect 4394 661 4405 677
rect 4451 668 4467 684
rect 4474 682 4504 734
rect 4538 730 4539 737
rect 4523 722 4539 730
rect 4510 690 4523 709
rect 4538 690 4568 706
rect 4510 674 4584 690
rect 4510 672 4523 674
rect 4538 672 4572 674
rect 4175 650 4188 652
rect 4203 650 4237 652
rect 4175 634 4237 650
rect 4281 645 4297 648
rect 4359 645 4389 656
rect 4437 652 4483 668
rect 4510 656 4584 672
rect 4437 650 4471 652
rect 4436 634 4483 650
rect 4510 634 4523 656
rect 4538 634 4568 656
rect 4595 634 4596 650
rect 4611 634 4624 793
rect 4654 689 4667 793
rect 4712 771 4713 781
rect 4733 779 4741 781
rect 4731 777 4741 779
rect 4728 771 4741 777
rect 4712 767 4741 771
rect 4746 767 4776 793
rect 4794 779 4810 781
rect 4882 779 4933 793
rect 4883 777 4947 779
rect 4990 777 5005 793
rect 5054 790 5084 793
rect 5054 787 5090 790
rect 5020 779 5036 781
rect 4794 767 4809 771
rect 4712 765 4809 767
rect 4837 765 5005 777
rect 5021 767 5036 771
rect 5054 768 5093 787
rect 5112 781 5119 782
rect 5118 774 5119 781
rect 5102 771 5103 774
rect 5118 771 5131 774
rect 5054 767 5084 768
rect 5093 767 5099 768
rect 5102 767 5131 771
rect 5021 766 5131 767
rect 5021 765 5137 766
rect 4696 757 4747 765
rect 4696 745 4721 757
rect 4728 745 4747 757
rect 4778 757 4828 765
rect 4778 749 4794 757
rect 4801 755 4828 757
rect 4837 755 5058 765
rect 4801 745 5058 755
rect 5087 757 5137 765
rect 5087 748 5103 757
rect 4696 737 4747 745
rect 4794 737 5058 745
rect 5084 745 5103 748
rect 5110 745 5137 757
rect 5084 737 5137 745
rect 4712 729 4713 737
rect 4728 729 4741 737
rect 4712 721 4728 729
rect 4709 714 4728 717
rect 4709 705 4731 714
rect 4682 695 4731 705
rect 4682 689 4712 695
rect 4731 690 4736 695
rect 4654 673 4728 689
rect 4746 681 4776 737
rect 4811 727 5019 737
rect 5054 733 5099 737
rect 5102 736 5103 737
rect 5118 736 5131 737
rect 4837 697 5026 727
rect 4852 694 5026 697
rect 4845 691 5026 694
rect 4654 671 4667 673
rect 4682 671 4716 673
rect 4654 655 4728 671
rect 4755 667 4768 681
rect 4783 667 4799 683
rect 4845 678 4856 691
rect -8 626 33 634
rect -8 600 7 626
rect 14 600 33 626
rect 97 622 159 634
rect 171 622 246 634
rect 304 622 379 634
rect 391 622 422 634
rect 428 622 463 634
rect 97 620 259 622
rect -8 592 33 600
rect 115 596 128 620
rect 143 618 158 620
rect -2 582 -1 592
rect 14 582 27 592
rect 42 582 72 596
rect 115 582 158 596
rect 182 593 189 600
rect 192 596 259 620
rect 291 620 463 622
rect 261 598 289 602
rect 291 598 371 620
rect 392 618 407 620
rect 261 596 371 598
rect 192 592 371 596
rect 165 582 195 592
rect 197 582 350 592
rect 358 582 388 592
rect 392 582 422 596
rect 450 582 463 620
rect 535 626 570 634
rect 535 600 536 626
rect 543 600 570 626
rect 478 582 508 596
rect 535 592 570 600
rect 572 626 613 634
rect 572 600 587 626
rect 594 600 613 626
rect 677 622 739 634
rect 751 622 826 634
rect 884 622 959 634
rect 971 622 1002 634
rect 1008 622 1043 634
rect 677 620 839 622
rect 572 592 613 600
rect 695 596 708 620
rect 723 618 738 620
rect 535 582 536 592
rect 551 582 564 592
rect 578 582 579 592
rect 594 582 607 592
rect 622 582 652 596
rect 695 582 738 596
rect 762 593 769 600
rect 772 596 839 620
rect 871 620 1043 622
rect 841 598 869 602
rect 871 598 951 620
rect 972 618 987 620
rect 841 596 951 598
rect 772 592 951 596
rect 745 582 775 592
rect 777 582 930 592
rect 938 582 968 592
rect 972 582 1002 596
rect 1030 582 1043 620
rect 1115 626 1150 634
rect 1115 600 1116 626
rect 1123 600 1150 626
rect 1058 582 1088 596
rect 1115 592 1150 600
rect 1152 626 1193 634
rect 1152 600 1167 626
rect 1174 600 1193 626
rect 1257 622 1319 634
rect 1331 622 1406 634
rect 1464 622 1539 634
rect 1551 622 1582 634
rect 1588 622 1623 634
rect 1257 620 1419 622
rect 1152 592 1193 600
rect 1275 596 1288 620
rect 1303 618 1318 620
rect 1115 582 1116 592
rect 1131 582 1144 592
rect 1158 582 1159 592
rect 1174 582 1187 592
rect 1202 582 1232 596
rect 1275 582 1318 596
rect 1342 593 1349 600
rect 1352 596 1419 620
rect 1451 620 1623 622
rect 1421 598 1449 602
rect 1451 598 1531 620
rect 1552 618 1567 620
rect 1421 596 1531 598
rect 1352 592 1531 596
rect 1325 582 1355 592
rect 1357 582 1510 592
rect 1518 582 1548 592
rect 1552 582 1582 596
rect 1610 582 1623 620
rect 1695 626 1730 634
rect 1695 600 1696 626
rect 1703 600 1730 626
rect 1638 582 1668 596
rect 1695 592 1730 600
rect 1732 626 1773 634
rect 1732 600 1747 626
rect 1754 600 1773 626
rect 1837 622 1899 634
rect 1911 622 1986 634
rect 2044 622 2119 634
rect 2131 622 2162 634
rect 2168 622 2203 634
rect 1837 620 1999 622
rect 1732 592 1773 600
rect 1855 596 1868 620
rect 1883 618 1898 620
rect 1695 582 1696 592
rect 1711 582 1724 592
rect 1738 582 1739 592
rect 1754 582 1767 592
rect 1782 582 1812 596
rect 1855 582 1898 596
rect 1922 593 1929 600
rect 1932 596 1999 620
rect 2031 620 2203 622
rect 2001 598 2029 602
rect 2031 598 2111 620
rect 2132 618 2147 620
rect 2001 596 2111 598
rect 1932 592 2111 596
rect 1905 582 1935 592
rect 1937 582 2090 592
rect 2098 582 2128 592
rect 2132 582 2162 596
rect 2190 582 2203 620
rect 2275 626 2310 634
rect 2275 600 2276 626
rect 2283 600 2310 626
rect 2218 582 2248 596
rect 2275 592 2310 600
rect 2312 626 2353 634
rect 2312 600 2327 626
rect 2334 600 2353 626
rect 2417 622 2479 634
rect 2491 622 2566 634
rect 2624 622 2699 634
rect 2711 622 2742 634
rect 2748 622 2783 634
rect 2417 620 2579 622
rect 2312 592 2353 600
rect 2435 596 2448 620
rect 2463 618 2478 620
rect 2275 582 2276 592
rect 2291 582 2304 592
rect 2318 582 2319 592
rect 2334 582 2347 592
rect 2362 582 2392 596
rect 2435 582 2478 596
rect 2502 593 2509 600
rect 2512 596 2579 620
rect 2611 620 2783 622
rect 2581 598 2609 602
rect 2611 598 2691 620
rect 2712 618 2727 620
rect 2581 596 2691 598
rect 2512 592 2691 596
rect 2485 582 2515 592
rect 2517 582 2670 592
rect 2678 582 2708 592
rect 2712 582 2742 596
rect 2770 582 2783 620
rect 2855 626 2890 634
rect 2855 600 2856 626
rect 2863 600 2890 626
rect 2798 582 2828 596
rect 2855 592 2890 600
rect 2892 626 2933 634
rect 2892 600 2907 626
rect 2914 600 2933 626
rect 2997 622 3059 634
rect 3071 622 3146 634
rect 3204 622 3279 634
rect 3291 622 3322 634
rect 3328 622 3363 634
rect 2997 620 3159 622
rect 2892 592 2933 600
rect 3015 596 3028 620
rect 3043 618 3058 620
rect 2855 582 2856 592
rect 2871 582 2884 592
rect 2898 582 2899 592
rect 2914 582 2927 592
rect 2942 582 2972 596
rect 3015 582 3058 596
rect 3082 593 3089 600
rect 3092 596 3159 620
rect 3191 620 3363 622
rect 3161 598 3189 602
rect 3191 598 3271 620
rect 3292 618 3307 620
rect 3161 596 3271 598
rect 3092 592 3271 596
rect 3065 582 3095 592
rect 3097 582 3250 592
rect 3258 582 3288 592
rect 3292 582 3322 596
rect 3350 582 3363 620
rect 3435 626 3470 634
rect 3435 600 3436 626
rect 3443 600 3470 626
rect 3378 582 3408 596
rect 3435 592 3470 600
rect 3472 626 3513 634
rect 3472 600 3487 626
rect 3494 600 3513 626
rect 3577 622 3639 634
rect 3651 622 3726 634
rect 3784 622 3859 634
rect 3871 622 3902 634
rect 3908 622 3943 634
rect 3577 620 3739 622
rect 3472 592 3513 600
rect 3595 596 3608 620
rect 3623 618 3638 620
rect 3435 582 3436 592
rect 3451 582 3464 592
rect 3478 582 3479 592
rect 3494 582 3507 592
rect 3522 582 3552 596
rect 3595 582 3638 596
rect 3662 593 3669 600
rect 3672 596 3739 620
rect 3771 620 3943 622
rect 3741 598 3769 602
rect 3771 598 3851 620
rect 3872 618 3887 620
rect 3741 596 3851 598
rect 3672 592 3851 596
rect 3645 582 3675 592
rect 3677 582 3830 592
rect 3838 582 3868 592
rect 3872 582 3902 596
rect 3930 582 3943 620
rect 4015 626 4050 634
rect 4015 600 4016 626
rect 4023 600 4050 626
rect 3958 582 3988 596
rect 4015 592 4050 600
rect 4052 626 4093 634
rect 4052 600 4067 626
rect 4074 600 4093 626
rect 4157 622 4219 634
rect 4231 622 4306 634
rect 4364 622 4439 634
rect 4451 622 4482 634
rect 4488 622 4523 634
rect 4157 620 4319 622
rect 4052 592 4093 600
rect 4175 596 4188 620
rect 4203 618 4218 620
rect 4015 582 4016 592
rect 4031 582 4044 592
rect 4058 582 4059 592
rect 4074 582 4087 592
rect 4102 582 4132 596
rect 4175 582 4218 596
rect 4242 593 4249 600
rect 4252 596 4319 620
rect 4351 620 4523 622
rect 4321 598 4349 602
rect 4351 598 4431 620
rect 4452 618 4467 620
rect 4321 596 4431 598
rect 4252 592 4431 596
rect 4225 582 4255 592
rect 4257 582 4410 592
rect 4418 582 4448 592
rect 4452 582 4482 596
rect 4510 582 4523 620
rect 4595 626 4630 634
rect 4638 633 4639 649
rect 4654 633 4667 655
rect 4682 633 4712 655
rect 4755 651 4817 667
rect 4845 660 4856 676
rect 4861 671 4871 691
rect 4881 671 4895 691
rect 4898 678 4907 691
rect 4923 678 4932 691
rect 4861 660 4895 671
rect 4898 660 4907 676
rect 4923 660 4932 676
rect 4939 671 4949 691
rect 4959 671 4973 691
rect 4974 678 4985 691
rect 4939 660 4973 671
rect 4974 660 4985 676
rect 5031 667 5047 683
rect 5054 681 5084 733
rect 5118 729 5119 736
rect 5103 721 5119 729
rect 5090 689 5103 708
rect 5118 689 5148 705
rect 5090 673 5164 689
rect 5090 671 5103 673
rect 5118 671 5152 673
rect 4755 649 4768 651
rect 4783 649 4817 651
rect 4755 633 4817 649
rect 4861 644 4877 647
rect 4939 644 4969 655
rect 5017 651 5063 667
rect 5090 655 5164 671
rect 5017 649 5051 651
rect 5016 633 5063 649
rect 5090 633 5103 655
rect 5118 633 5148 655
rect 5175 633 5176 649
rect 5191 633 5204 793
rect 5234 689 5247 793
rect 5292 771 5293 781
rect 5313 779 5321 781
rect 5311 777 5321 779
rect 5308 771 5321 777
rect 5292 767 5321 771
rect 5326 767 5356 793
rect 5374 779 5390 781
rect 5462 779 5513 793
rect 5463 777 5527 779
rect 5570 777 5585 793
rect 5634 790 5664 793
rect 5634 787 5670 790
rect 5600 779 5616 781
rect 5374 767 5389 771
rect 5292 765 5389 767
rect 5417 765 5585 777
rect 5601 767 5616 771
rect 5634 768 5673 787
rect 5692 781 5699 782
rect 5698 774 5699 781
rect 5682 771 5683 774
rect 5698 771 5711 774
rect 5634 767 5664 768
rect 5673 767 5679 768
rect 5682 767 5711 771
rect 5601 766 5711 767
rect 5601 765 5717 766
rect 5276 757 5327 765
rect 5276 745 5301 757
rect 5308 745 5327 757
rect 5358 757 5408 765
rect 5358 749 5374 757
rect 5381 755 5408 757
rect 5417 755 5638 765
rect 5381 745 5638 755
rect 5667 757 5717 765
rect 5667 748 5683 757
rect 5276 737 5327 745
rect 5374 737 5638 745
rect 5664 745 5683 748
rect 5690 745 5717 757
rect 5664 737 5717 745
rect 5292 729 5293 737
rect 5308 729 5321 737
rect 5292 721 5308 729
rect 5289 714 5308 717
rect 5289 705 5311 714
rect 5262 695 5311 705
rect 5262 689 5292 695
rect 5311 690 5316 695
rect 5234 673 5308 689
rect 5326 681 5356 737
rect 5391 727 5599 737
rect 5634 733 5679 737
rect 5682 736 5683 737
rect 5698 736 5711 737
rect 5417 697 5606 727
rect 5432 694 5606 697
rect 5425 691 5606 694
rect 5234 671 5247 673
rect 5262 671 5296 673
rect 5234 655 5308 671
rect 5335 667 5348 681
rect 5363 667 5379 683
rect 5425 678 5436 691
rect 5218 633 5219 649
rect 5234 633 5247 655
rect 5262 633 5292 655
rect 5335 651 5397 667
rect 5425 660 5436 676
rect 5441 671 5451 691
rect 5461 671 5475 691
rect 5478 678 5487 691
rect 5503 678 5512 691
rect 5441 660 5475 671
rect 5478 660 5487 676
rect 5503 660 5512 676
rect 5519 671 5529 691
rect 5539 671 5553 691
rect 5554 678 5565 691
rect 5519 660 5553 671
rect 5554 660 5565 676
rect 5611 667 5627 683
rect 5634 681 5664 733
rect 5698 729 5699 736
rect 5683 721 5699 729
rect 5670 689 5683 708
rect 5698 689 5728 705
rect 5670 673 5744 689
rect 5670 671 5683 673
rect 5698 671 5732 673
rect 5335 649 5348 651
rect 5363 649 5397 651
rect 5335 633 5397 649
rect 5441 644 5457 647
rect 5519 644 5549 655
rect 5597 651 5643 667
rect 5670 655 5744 671
rect 5597 649 5631 651
rect 5596 633 5643 649
rect 5670 633 5683 655
rect 5698 633 5728 655
rect 5755 633 5756 649
rect 5771 633 5784 793
rect 5814 689 5827 793
rect 5872 771 5873 781
rect 5893 779 5901 781
rect 5891 777 5901 779
rect 5888 771 5901 777
rect 5872 767 5901 771
rect 5906 767 5936 793
rect 5954 779 5970 781
rect 6042 779 6093 793
rect 6043 777 6107 779
rect 6150 777 6165 793
rect 6214 790 6244 793
rect 6214 787 6250 790
rect 6180 779 6196 781
rect 5954 767 5969 771
rect 5872 765 5969 767
rect 5997 765 6165 777
rect 6181 767 6196 771
rect 6214 768 6253 787
rect 6272 781 6279 782
rect 6278 774 6279 781
rect 6262 771 6263 774
rect 6278 771 6291 774
rect 6214 767 6244 768
rect 6253 767 6259 768
rect 6262 767 6291 771
rect 6181 766 6291 767
rect 6181 765 6297 766
rect 5856 757 5907 765
rect 5856 745 5881 757
rect 5888 745 5907 757
rect 5938 757 5988 765
rect 5938 749 5954 757
rect 5961 755 5988 757
rect 5997 755 6218 765
rect 5961 745 6218 755
rect 6247 757 6297 765
rect 6247 748 6263 757
rect 5856 737 5907 745
rect 5954 737 6218 745
rect 6244 745 6263 748
rect 6270 745 6297 757
rect 6244 737 6297 745
rect 5872 729 5873 737
rect 5888 729 5901 737
rect 5872 721 5888 729
rect 5869 714 5888 717
rect 5869 705 5891 714
rect 5842 695 5891 705
rect 5842 689 5872 695
rect 5891 690 5896 695
rect 5814 673 5888 689
rect 5906 681 5936 737
rect 5971 727 6179 737
rect 6214 733 6259 737
rect 6262 736 6263 737
rect 6278 736 6291 737
rect 5997 697 6186 727
rect 6012 694 6186 697
rect 6005 691 6186 694
rect 5814 671 5827 673
rect 5842 671 5876 673
rect 5814 655 5888 671
rect 5915 667 5928 681
rect 5943 667 5959 683
rect 6005 678 6016 691
rect 5798 633 5799 649
rect 5814 633 5827 655
rect 5842 633 5872 655
rect 5915 651 5977 667
rect 6005 660 6016 676
rect 6021 671 6031 691
rect 6041 671 6055 691
rect 6058 678 6067 691
rect 6083 678 6092 691
rect 6021 660 6055 671
rect 6058 660 6067 676
rect 6083 660 6092 676
rect 6099 671 6109 691
rect 6119 671 6133 691
rect 6134 678 6145 691
rect 6099 660 6133 671
rect 6134 660 6145 676
rect 6191 667 6207 683
rect 6214 681 6244 733
rect 6278 729 6279 736
rect 6263 721 6279 729
rect 6250 689 6263 708
rect 6278 689 6308 705
rect 6250 673 6324 689
rect 6250 671 6263 673
rect 6278 671 6312 673
rect 5915 649 5928 651
rect 5943 649 5977 651
rect 5915 633 5977 649
rect 6021 644 6037 647
rect 6099 644 6129 655
rect 6177 651 6223 667
rect 6250 655 6324 671
rect 6177 649 6211 651
rect 6176 633 6223 649
rect 6250 633 6263 655
rect 6278 633 6308 655
rect 6335 633 6336 649
rect 6351 633 6364 793
rect 6394 689 6407 793
rect 6452 771 6453 781
rect 6473 779 6481 781
rect 6471 777 6481 779
rect 6468 771 6481 777
rect 6452 767 6481 771
rect 6486 767 6516 793
rect 6534 779 6550 781
rect 6622 779 6673 793
rect 6623 777 6687 779
rect 6730 777 6745 793
rect 6794 790 6824 793
rect 6794 787 6830 790
rect 6760 779 6776 781
rect 6534 767 6549 771
rect 6452 765 6549 767
rect 6577 765 6745 777
rect 6761 767 6776 771
rect 6794 768 6833 787
rect 6852 781 6859 782
rect 6858 774 6859 781
rect 6842 771 6843 774
rect 6858 771 6871 774
rect 6794 767 6824 768
rect 6833 767 6839 768
rect 6842 767 6871 771
rect 6761 766 6871 767
rect 6761 765 6877 766
rect 6436 757 6487 765
rect 6436 745 6461 757
rect 6468 745 6487 757
rect 6518 757 6568 765
rect 6518 749 6534 757
rect 6541 755 6568 757
rect 6577 755 6798 765
rect 6541 745 6798 755
rect 6827 757 6877 765
rect 6827 748 6843 757
rect 6436 737 6487 745
rect 6534 737 6798 745
rect 6824 745 6843 748
rect 6850 745 6877 757
rect 6824 737 6877 745
rect 6452 729 6453 737
rect 6468 729 6481 737
rect 6452 721 6468 729
rect 6449 714 6468 717
rect 6449 705 6471 714
rect 6422 695 6471 705
rect 6422 689 6452 695
rect 6471 690 6476 695
rect 6394 673 6468 689
rect 6486 681 6516 737
rect 6551 727 6759 737
rect 6794 733 6839 737
rect 6842 736 6843 737
rect 6858 736 6871 737
rect 6577 697 6766 727
rect 6592 694 6766 697
rect 6585 691 6766 694
rect 6394 671 6407 673
rect 6422 671 6456 673
rect 6394 655 6468 671
rect 6495 667 6508 681
rect 6523 667 6539 683
rect 6585 678 6596 691
rect 6378 633 6379 649
rect 6394 633 6407 655
rect 6422 633 6452 655
rect 6495 651 6557 667
rect 6585 660 6596 676
rect 6601 671 6611 691
rect 6621 671 6635 691
rect 6638 678 6647 691
rect 6663 678 6672 691
rect 6601 660 6635 671
rect 6638 660 6647 676
rect 6663 660 6672 676
rect 6679 671 6689 691
rect 6699 671 6713 691
rect 6714 678 6725 691
rect 6679 660 6713 671
rect 6714 660 6725 676
rect 6771 667 6787 683
rect 6794 681 6824 733
rect 6858 729 6859 736
rect 6843 721 6859 729
rect 6830 689 6843 708
rect 6858 689 6888 705
rect 6830 673 6904 689
rect 6830 671 6843 673
rect 6858 671 6892 673
rect 6495 649 6508 651
rect 6523 649 6557 651
rect 6495 633 6557 649
rect 6601 644 6617 647
rect 6679 644 6709 655
rect 6757 651 6803 667
rect 6830 655 6904 671
rect 6757 649 6791 651
rect 6756 633 6803 649
rect 6830 633 6843 655
rect 6858 633 6888 655
rect 6915 633 6916 649
rect 6931 633 6944 793
rect 4595 600 4596 626
rect 4603 600 4630 626
rect 4538 582 4568 596
rect 4595 592 4630 600
rect 4632 625 4673 633
rect 4632 599 4647 625
rect 4654 599 4673 625
rect 4737 621 4799 633
rect 4811 621 4886 633
rect 4944 621 5019 633
rect 5031 621 5062 633
rect 5068 621 5103 633
rect 4737 619 4899 621
rect 4755 601 4768 619
rect 4783 617 4798 619
rect 4595 582 4596 592
rect 4611 582 4624 592
rect 4632 591 4673 599
rect 4756 595 4768 601
rect 4832 601 4899 619
rect 4931 619 5103 621
rect 4931 601 5011 619
rect 5032 617 5047 619
rect -2 581 4624 582
rect 4638 581 4639 591
rect 4654 581 4667 591
rect 4682 581 4712 595
rect 4756 581 4798 595
rect 4822 592 4829 599
rect 4832 591 5011 601
rect 4805 581 4835 591
rect 4837 581 4990 591
rect 4998 581 5028 591
rect 5032 581 5062 595
rect 5090 581 5103 619
rect 5175 625 5210 633
rect 5175 599 5176 625
rect 5183 599 5210 625
rect 5118 581 5148 595
rect 5175 591 5210 599
rect 5212 625 5253 633
rect 5212 599 5227 625
rect 5234 599 5253 625
rect 5317 621 5379 633
rect 5391 621 5466 633
rect 5524 621 5599 633
rect 5611 621 5642 633
rect 5648 621 5683 633
rect 5317 619 5479 621
rect 5335 601 5348 619
rect 5363 617 5378 619
rect 5212 591 5253 599
rect 5336 595 5348 601
rect 5412 601 5479 619
rect 5511 619 5683 621
rect 5511 601 5591 619
rect 5612 617 5627 619
rect 5175 581 5176 591
rect 5191 581 5204 591
rect 5218 581 5219 591
rect 5234 581 5247 591
rect 5262 581 5292 595
rect 5336 581 5378 595
rect 5402 592 5409 599
rect 5412 591 5591 601
rect 5385 581 5415 591
rect 5417 581 5570 591
rect 5578 581 5608 591
rect 5612 581 5642 595
rect 5670 581 5683 619
rect 5755 625 5790 633
rect 5755 599 5756 625
rect 5763 599 5790 625
rect 5698 581 5728 595
rect 5755 591 5790 599
rect 5792 625 5833 633
rect 5792 599 5807 625
rect 5814 599 5833 625
rect 5897 621 5959 633
rect 5971 621 6046 633
rect 6104 621 6179 633
rect 6191 621 6222 633
rect 6228 621 6263 633
rect 5897 619 6059 621
rect 5915 601 5928 619
rect 5943 617 5958 619
rect 5792 591 5833 599
rect 5916 595 5928 601
rect 5992 601 6059 619
rect 6091 619 6263 621
rect 6091 601 6171 619
rect 6192 617 6207 619
rect 5755 581 5756 591
rect 5771 581 5784 591
rect 5798 581 5799 591
rect 5814 581 5827 591
rect 5842 581 5872 595
rect 5916 581 5958 595
rect 5982 592 5989 599
rect 5992 591 6171 601
rect 5965 581 5995 591
rect 5997 581 6150 591
rect 6158 581 6188 591
rect 6192 581 6222 595
rect 6250 581 6263 619
rect 6335 625 6370 633
rect 6335 599 6336 625
rect 6343 599 6370 625
rect 6278 581 6308 595
rect 6335 591 6370 599
rect 6372 625 6413 633
rect 6372 599 6387 625
rect 6394 599 6413 625
rect 6477 621 6539 633
rect 6551 621 6626 633
rect 6684 621 6759 633
rect 6771 621 6802 633
rect 6808 621 6843 633
rect 6477 619 6639 621
rect 6495 601 6508 619
rect 6523 617 6538 619
rect 6372 591 6413 599
rect 6496 595 6508 601
rect 6572 601 6639 619
rect 6671 619 6843 621
rect 6671 601 6751 619
rect 6772 617 6787 619
rect 6335 581 6336 591
rect 6351 581 6364 591
rect 6378 581 6379 591
rect 6394 581 6407 591
rect 6422 581 6452 595
rect 6496 581 6538 595
rect 6562 592 6569 599
rect 6572 591 6751 601
rect 6545 581 6575 591
rect 6577 581 6730 591
rect 6738 581 6768 591
rect 6772 581 6802 595
rect 6830 581 6843 619
rect 6915 625 6950 633
rect 6915 599 6916 625
rect 6923 599 6950 625
rect 6858 581 6888 595
rect 6915 591 6950 599
rect 6915 581 6916 591
rect 6931 581 6944 591
rect -2 576 6944 581
rect -1 568 6944 576
rect 14 538 27 568
rect 42 550 72 568
rect 115 554 129 568
rect 165 554 385 568
rect 116 552 129 554
rect 82 540 97 552
rect 79 538 101 540
rect 106 538 136 552
rect 197 550 350 554
rect 179 538 371 550
rect 414 538 444 552
rect 450 538 463 568
rect 478 550 508 568
rect 551 538 564 568
rect 594 538 607 568
rect 622 550 652 568
rect 695 554 709 568
rect 745 554 965 568
rect 696 552 709 554
rect 662 540 677 552
rect 659 538 681 540
rect 686 538 716 552
rect 777 550 930 554
rect 759 538 951 550
rect 994 538 1024 552
rect 1030 538 1043 568
rect 1058 550 1088 568
rect 1131 538 1144 568
rect 1174 538 1187 568
rect 1202 550 1232 568
rect 1275 554 1289 568
rect 1325 554 1545 568
rect 1276 552 1289 554
rect 1242 540 1257 552
rect 1239 538 1261 540
rect 1266 538 1296 552
rect 1357 550 1510 554
rect 1339 538 1531 550
rect 1574 538 1604 552
rect 1610 538 1623 568
rect 1638 550 1668 568
rect 1711 538 1724 568
rect 1754 538 1767 568
rect 1782 550 1812 568
rect 1855 554 1869 568
rect 1905 554 2125 568
rect 1856 552 1869 554
rect 1822 540 1837 552
rect 1819 538 1841 540
rect 1846 538 1876 552
rect 1937 550 2090 554
rect 1919 538 2111 550
rect 2154 538 2184 552
rect 2190 538 2203 568
rect 2218 550 2248 568
rect 2291 538 2304 568
rect 2334 538 2347 568
rect 2362 550 2392 568
rect 2435 554 2449 568
rect 2485 554 2705 568
rect 2436 552 2449 554
rect 2402 540 2417 552
rect 2399 538 2421 540
rect 2426 538 2456 552
rect 2517 550 2670 554
rect 2499 538 2691 550
rect 2734 538 2764 552
rect 2770 538 2783 568
rect 2798 550 2828 568
rect 2871 538 2884 568
rect 2914 538 2927 568
rect 2942 550 2972 568
rect 3015 554 3029 568
rect 3065 554 3285 568
rect 3016 552 3029 554
rect 2982 540 2997 552
rect 2979 538 3001 540
rect 3006 538 3036 552
rect 3097 550 3250 554
rect 3079 538 3271 550
rect 3314 538 3344 552
rect 3350 538 3363 568
rect 3378 550 3408 568
rect 3451 538 3464 568
rect 3494 538 3507 568
rect 3522 550 3552 568
rect 3595 554 3609 568
rect 3645 554 3865 568
rect 3596 552 3609 554
rect 3562 540 3577 552
rect 3559 538 3581 540
rect 3586 538 3616 552
rect 3677 550 3830 554
rect 3659 538 3851 550
rect 3894 538 3924 552
rect 3930 538 3943 568
rect 3958 550 3988 568
rect 4031 538 4044 568
rect 4074 538 4087 568
rect 4102 550 4132 568
rect 4175 554 4189 568
rect 4225 554 4445 568
rect 4176 552 4189 554
rect 4142 540 4157 552
rect 4139 538 4161 540
rect 4166 538 4196 552
rect 4257 550 4410 554
rect 4239 538 4431 550
rect 4474 538 4504 552
rect 4510 538 4523 568
rect 4538 550 4568 568
rect 4611 567 6944 568
rect 4611 538 4624 567
rect -1 537 4624 538
rect 4654 537 4667 567
rect 4682 549 4712 567
rect 4756 551 4769 567
rect 4805 553 5025 567
rect 4722 539 4737 551
rect 4719 537 4741 539
rect 4746 537 4776 551
rect 4837 549 4990 553
rect 4819 537 5011 549
rect 5054 537 5084 551
rect 5090 537 5103 567
rect 5118 549 5148 567
rect 5191 537 5204 567
rect 5234 537 5247 567
rect 5262 549 5292 567
rect 5336 551 5349 567
rect 5385 553 5605 567
rect 5302 539 5317 551
rect 5299 537 5321 539
rect 5326 537 5356 551
rect 5417 549 5570 553
rect 5399 537 5591 549
rect 5634 537 5664 551
rect 5670 537 5683 567
rect 5698 549 5728 567
rect 5771 537 5784 567
rect 5814 537 5827 567
rect 5842 549 5872 567
rect 5916 551 5929 567
rect 5965 553 6185 567
rect 5882 539 5897 551
rect 5879 537 5901 539
rect 5906 537 5936 551
rect 5997 549 6150 553
rect 5979 537 6171 549
rect 6214 537 6244 551
rect 6250 537 6263 567
rect 6278 549 6308 567
rect 6351 537 6364 567
rect 6394 537 6407 567
rect 6422 549 6452 567
rect 6496 551 6509 567
rect 6545 553 6765 567
rect 6462 539 6477 551
rect 6459 537 6481 539
rect 6486 537 6516 551
rect 6577 549 6730 553
rect 6559 537 6751 549
rect 6794 537 6824 551
rect 6830 537 6843 567
rect 6858 549 6888 567
rect 6931 537 6944 567
rect -1 524 6944 537
rect 14 420 27 524
rect 72 502 73 512
rect 88 502 101 512
rect 72 498 101 502
rect 106 498 136 524
rect 154 510 170 512
rect 242 510 295 524
rect 243 508 307 510
rect 350 508 365 524
rect 414 521 444 524
rect 414 518 450 521
rect 380 510 396 512
rect 154 498 169 502
rect 72 496 169 498
rect 197 496 365 508
rect 381 498 396 502
rect 414 499 453 518
rect 472 512 479 513
rect 478 505 479 512
rect 462 502 463 505
rect 478 502 491 505
rect 414 498 444 499
rect 453 498 459 499
rect 462 498 491 502
rect 381 497 491 498
rect 381 496 497 497
rect 56 488 107 496
rect 56 476 81 488
rect 88 476 107 488
rect 138 488 188 496
rect 138 480 154 488
rect 161 486 188 488
rect 197 486 418 496
rect 161 476 418 486
rect 447 488 497 496
rect 447 479 463 488
rect 56 468 107 476
rect 154 468 418 476
rect 444 476 463 479
rect 470 476 497 488
rect 444 468 497 476
rect 72 460 73 468
rect 88 460 101 468
rect 72 452 88 460
rect 69 445 88 448
rect 69 436 91 445
rect 42 426 91 436
rect 42 420 72 426
rect 91 421 96 426
rect 14 404 88 420
rect 106 412 136 468
rect 171 458 379 468
rect 414 464 459 468
rect 462 467 463 468
rect 478 467 491 468
rect 197 428 386 458
rect 212 425 386 428
rect 205 422 386 425
rect 14 402 27 404
rect 42 402 76 404
rect 14 386 88 402
rect 115 398 128 412
rect 143 398 159 414
rect 205 409 216 422
rect -2 364 -1 380
rect 14 364 27 386
rect 42 364 72 386
rect 115 382 177 398
rect 205 391 216 407
rect 221 402 231 422
rect 241 402 255 422
rect 258 409 267 422
rect 283 409 292 422
rect 221 391 255 402
rect 258 391 267 407
rect 283 391 292 407
rect 299 402 309 422
rect 319 402 333 422
rect 334 409 345 422
rect 299 391 333 402
rect 334 391 345 407
rect 391 398 407 414
rect 414 412 444 464
rect 478 460 479 467
rect 463 452 479 460
rect 450 420 463 439
rect 478 420 508 436
rect 450 404 524 420
rect 450 402 463 404
rect 478 402 512 404
rect 115 380 128 382
rect 143 380 177 382
rect 115 364 177 380
rect 221 375 237 378
rect 299 375 329 386
rect 377 382 423 398
rect 450 386 524 402
rect 377 380 411 382
rect 376 364 423 380
rect 450 364 463 386
rect 478 364 508 386
rect 535 364 536 380
rect 551 364 564 524
rect 594 420 607 524
rect 652 502 653 512
rect 668 502 681 512
rect 652 498 681 502
rect 686 498 716 524
rect 734 510 750 512
rect 822 510 875 524
rect 823 508 887 510
rect 930 508 945 524
rect 994 521 1024 524
rect 994 518 1030 521
rect 960 510 976 512
rect 734 498 749 502
rect 652 496 749 498
rect 777 496 945 508
rect 961 498 976 502
rect 994 499 1033 518
rect 1052 512 1059 513
rect 1058 505 1059 512
rect 1042 502 1043 505
rect 1058 502 1071 505
rect 994 498 1024 499
rect 1033 498 1039 499
rect 1042 498 1071 502
rect 961 497 1071 498
rect 961 496 1077 497
rect 636 488 687 496
rect 636 476 661 488
rect 668 476 687 488
rect 718 488 768 496
rect 718 480 734 488
rect 741 486 768 488
rect 777 486 998 496
rect 741 476 998 486
rect 1027 488 1077 496
rect 1027 479 1043 488
rect 636 468 687 476
rect 734 468 998 476
rect 1024 476 1043 479
rect 1050 476 1077 488
rect 1024 468 1077 476
rect 652 460 653 468
rect 668 460 681 468
rect 652 452 668 460
rect 649 445 668 448
rect 649 436 671 445
rect 622 426 671 436
rect 622 420 652 426
rect 671 421 676 426
rect 594 404 668 420
rect 686 412 716 468
rect 751 458 959 468
rect 994 464 1039 468
rect 1042 467 1043 468
rect 1058 467 1071 468
rect 777 428 966 458
rect 792 425 966 428
rect 785 422 966 425
rect 594 402 607 404
rect 622 402 656 404
rect 594 386 668 402
rect 695 398 708 412
rect 723 398 739 414
rect 785 409 796 422
rect 578 364 579 380
rect 594 364 607 386
rect 622 364 652 386
rect 695 382 757 398
rect 785 391 796 407
rect 801 402 811 422
rect 821 402 835 422
rect 838 409 847 422
rect 863 409 872 422
rect 801 391 835 402
rect 838 391 847 407
rect 863 391 872 407
rect 879 402 889 422
rect 899 402 913 422
rect 914 409 925 422
rect 879 391 913 402
rect 914 391 925 407
rect 971 398 987 414
rect 994 412 1024 464
rect 1058 460 1059 467
rect 1043 452 1059 460
rect 1030 420 1043 439
rect 1058 420 1088 436
rect 1030 404 1104 420
rect 1030 402 1043 404
rect 1058 402 1092 404
rect 695 380 708 382
rect 723 380 757 382
rect 695 364 757 380
rect 801 375 817 378
rect 879 375 909 386
rect 957 382 1003 398
rect 1030 386 1104 402
rect 957 380 991 382
rect 956 364 1003 380
rect 1030 364 1043 386
rect 1058 364 1088 386
rect 1115 364 1116 380
rect 1131 364 1144 524
rect 1174 420 1187 524
rect 1232 502 1233 512
rect 1248 502 1261 512
rect 1232 498 1261 502
rect 1266 498 1296 524
rect 1314 510 1330 512
rect 1402 510 1455 524
rect 1403 508 1467 510
rect 1510 508 1525 524
rect 1574 521 1604 524
rect 1574 518 1610 521
rect 1540 510 1556 512
rect 1314 498 1329 502
rect 1232 496 1329 498
rect 1357 496 1525 508
rect 1541 498 1556 502
rect 1574 499 1613 518
rect 1632 512 1639 513
rect 1638 505 1639 512
rect 1622 502 1623 505
rect 1638 502 1651 505
rect 1574 498 1604 499
rect 1613 498 1619 499
rect 1622 498 1651 502
rect 1541 497 1651 498
rect 1541 496 1657 497
rect 1216 488 1267 496
rect 1216 476 1241 488
rect 1248 476 1267 488
rect 1298 488 1348 496
rect 1298 480 1314 488
rect 1321 486 1348 488
rect 1357 486 1578 496
rect 1321 476 1578 486
rect 1607 488 1657 496
rect 1607 479 1623 488
rect 1216 468 1267 476
rect 1314 468 1578 476
rect 1604 476 1623 479
rect 1630 476 1657 488
rect 1604 468 1657 476
rect 1232 460 1233 468
rect 1248 460 1261 468
rect 1232 452 1248 460
rect 1229 445 1248 448
rect 1229 436 1251 445
rect 1202 426 1251 436
rect 1202 420 1232 426
rect 1251 421 1256 426
rect 1174 404 1248 420
rect 1266 412 1296 468
rect 1331 458 1539 468
rect 1574 464 1619 468
rect 1622 467 1623 468
rect 1638 467 1651 468
rect 1357 428 1546 458
rect 1372 425 1546 428
rect 1365 422 1546 425
rect 1174 402 1187 404
rect 1202 402 1236 404
rect 1174 386 1248 402
rect 1275 398 1288 412
rect 1303 398 1319 414
rect 1365 409 1376 422
rect 1158 364 1159 380
rect 1174 364 1187 386
rect 1202 364 1232 386
rect 1275 382 1337 398
rect 1365 391 1376 407
rect 1381 402 1391 422
rect 1401 402 1415 422
rect 1418 409 1427 422
rect 1443 409 1452 422
rect 1381 391 1415 402
rect 1418 391 1427 407
rect 1443 391 1452 407
rect 1459 402 1469 422
rect 1479 402 1493 422
rect 1494 409 1505 422
rect 1459 391 1493 402
rect 1494 391 1505 407
rect 1551 398 1567 414
rect 1574 412 1604 464
rect 1638 460 1639 467
rect 1623 452 1639 460
rect 1610 420 1623 439
rect 1638 420 1668 436
rect 1610 404 1684 420
rect 1610 402 1623 404
rect 1638 402 1672 404
rect 1275 380 1288 382
rect 1303 380 1337 382
rect 1275 364 1337 380
rect 1381 375 1397 378
rect 1459 375 1489 386
rect 1537 382 1583 398
rect 1610 386 1684 402
rect 1537 380 1571 382
rect 1536 364 1583 380
rect 1610 364 1623 386
rect 1638 364 1668 386
rect 1695 364 1696 380
rect 1711 364 1724 524
rect 1754 420 1767 524
rect 1812 502 1813 512
rect 1828 502 1841 512
rect 1812 498 1841 502
rect 1846 498 1876 524
rect 1894 510 1910 512
rect 1982 510 2035 524
rect 1983 508 2047 510
rect 2090 508 2105 524
rect 2154 521 2184 524
rect 2154 518 2190 521
rect 2120 510 2136 512
rect 1894 498 1909 502
rect 1812 496 1909 498
rect 1937 496 2105 508
rect 2121 498 2136 502
rect 2154 499 2193 518
rect 2212 512 2219 513
rect 2218 505 2219 512
rect 2202 502 2203 505
rect 2218 502 2231 505
rect 2154 498 2184 499
rect 2193 498 2199 499
rect 2202 498 2231 502
rect 2121 497 2231 498
rect 2121 496 2237 497
rect 1796 488 1847 496
rect 1796 476 1821 488
rect 1828 476 1847 488
rect 1878 488 1928 496
rect 1878 480 1894 488
rect 1901 486 1928 488
rect 1937 486 2158 496
rect 1901 476 2158 486
rect 2187 488 2237 496
rect 2187 479 2203 488
rect 1796 468 1847 476
rect 1894 468 2158 476
rect 2184 476 2203 479
rect 2210 476 2237 488
rect 2184 468 2237 476
rect 1812 460 1813 468
rect 1828 460 1841 468
rect 1812 452 1828 460
rect 1809 445 1828 448
rect 1809 436 1831 445
rect 1782 426 1831 436
rect 1782 420 1812 426
rect 1831 421 1836 426
rect 1754 404 1828 420
rect 1846 412 1876 468
rect 1911 458 2119 468
rect 2154 464 2199 468
rect 2202 467 2203 468
rect 2218 467 2231 468
rect 1937 428 2126 458
rect 1952 425 2126 428
rect 1945 422 2126 425
rect 1754 402 1767 404
rect 1782 402 1816 404
rect 1754 386 1828 402
rect 1855 398 1868 412
rect 1883 398 1899 414
rect 1945 409 1956 422
rect 1738 364 1739 380
rect 1754 364 1767 386
rect 1782 364 1812 386
rect 1855 382 1917 398
rect 1945 391 1956 407
rect 1961 402 1971 422
rect 1981 402 1995 422
rect 1998 409 2007 422
rect 2023 409 2032 422
rect 1961 391 1995 402
rect 1998 391 2007 407
rect 2023 391 2032 407
rect 2039 402 2049 422
rect 2059 402 2073 422
rect 2074 409 2085 422
rect 2039 391 2073 402
rect 2074 391 2085 407
rect 2131 398 2147 414
rect 2154 412 2184 464
rect 2218 460 2219 467
rect 2203 452 2219 460
rect 2190 420 2203 439
rect 2218 420 2248 436
rect 2190 404 2264 420
rect 2190 402 2203 404
rect 2218 402 2252 404
rect 1855 380 1868 382
rect 1883 380 1917 382
rect 1855 364 1917 380
rect 1961 375 1977 378
rect 2039 375 2069 386
rect 2117 382 2163 398
rect 2190 386 2264 402
rect 2117 380 2151 382
rect 2116 364 2163 380
rect 2190 364 2203 386
rect 2218 364 2248 386
rect 2275 364 2276 380
rect 2291 364 2304 524
rect 2334 420 2347 524
rect 2392 502 2393 512
rect 2408 502 2421 512
rect 2392 498 2421 502
rect 2426 498 2456 524
rect 2474 510 2490 512
rect 2562 510 2615 524
rect 2563 508 2627 510
rect 2670 508 2685 524
rect 2734 521 2764 524
rect 2734 518 2770 521
rect 2700 510 2716 512
rect 2474 498 2489 502
rect 2392 496 2489 498
rect 2517 496 2685 508
rect 2701 498 2716 502
rect 2734 499 2773 518
rect 2792 512 2799 513
rect 2798 505 2799 512
rect 2782 502 2783 505
rect 2798 502 2811 505
rect 2734 498 2764 499
rect 2773 498 2779 499
rect 2782 498 2811 502
rect 2701 497 2811 498
rect 2701 496 2817 497
rect 2376 488 2427 496
rect 2376 476 2401 488
rect 2408 476 2427 488
rect 2458 488 2508 496
rect 2458 480 2474 488
rect 2481 486 2508 488
rect 2517 486 2738 496
rect 2481 476 2738 486
rect 2767 488 2817 496
rect 2767 479 2783 488
rect 2376 468 2427 476
rect 2474 468 2738 476
rect 2764 476 2783 479
rect 2790 476 2817 488
rect 2764 468 2817 476
rect 2392 460 2393 468
rect 2408 460 2421 468
rect 2392 452 2408 460
rect 2389 445 2408 448
rect 2389 436 2411 445
rect 2362 426 2411 436
rect 2362 420 2392 426
rect 2411 421 2416 426
rect 2334 404 2408 420
rect 2426 412 2456 468
rect 2491 458 2699 468
rect 2734 464 2779 468
rect 2782 467 2783 468
rect 2798 467 2811 468
rect 2517 428 2706 458
rect 2532 425 2706 428
rect 2525 422 2706 425
rect 2334 402 2347 404
rect 2362 402 2396 404
rect 2334 386 2408 402
rect 2435 398 2448 412
rect 2463 398 2479 414
rect 2525 409 2536 422
rect 2318 364 2319 380
rect 2334 364 2347 386
rect 2362 364 2392 386
rect 2435 382 2497 398
rect 2525 391 2536 407
rect 2541 402 2551 422
rect 2561 402 2575 422
rect 2578 409 2587 422
rect 2603 409 2612 422
rect 2541 391 2575 402
rect 2578 391 2587 407
rect 2603 391 2612 407
rect 2619 402 2629 422
rect 2639 402 2653 422
rect 2654 409 2665 422
rect 2619 391 2653 402
rect 2654 391 2665 407
rect 2711 398 2727 414
rect 2734 412 2764 464
rect 2798 460 2799 467
rect 2783 452 2799 460
rect 2770 420 2783 439
rect 2798 420 2828 436
rect 2770 404 2844 420
rect 2770 402 2783 404
rect 2798 402 2832 404
rect 2435 380 2448 382
rect 2463 380 2497 382
rect 2435 364 2497 380
rect 2541 375 2557 378
rect 2619 375 2649 386
rect 2697 382 2743 398
rect 2770 386 2844 402
rect 2697 380 2731 382
rect 2696 364 2743 380
rect 2770 364 2783 386
rect 2798 364 2828 386
rect 2855 364 2856 380
rect 2871 364 2884 524
rect 2914 420 2927 524
rect 2972 502 2973 512
rect 2988 502 3001 512
rect 2972 498 3001 502
rect 3006 498 3036 524
rect 3054 510 3070 512
rect 3142 510 3195 524
rect 3143 508 3205 510
rect 3250 508 3265 524
rect 3314 521 3344 524
rect 3314 518 3350 521
rect 3280 510 3296 512
rect 3054 498 3069 502
rect 2972 496 3069 498
rect 3097 496 3265 508
rect 3281 498 3296 502
rect 3314 499 3353 518
rect 3372 512 3379 513
rect 3378 505 3379 512
rect 3362 502 3363 505
rect 3378 502 3391 505
rect 3314 498 3344 499
rect 3353 498 3359 499
rect 3362 498 3391 502
rect 3281 497 3391 498
rect 3281 496 3397 497
rect 2956 488 3007 496
rect 2956 476 2981 488
rect 2988 476 3007 488
rect 3038 488 3088 496
rect 3038 480 3054 488
rect 3061 486 3088 488
rect 3097 486 3318 496
rect 3061 476 3318 486
rect 3347 488 3397 496
rect 3347 479 3363 488
rect 2956 468 3007 476
rect 3054 468 3318 476
rect 3344 476 3363 479
rect 3370 476 3397 488
rect 3344 468 3397 476
rect 2972 460 2973 468
rect 2988 460 3001 468
rect 2972 452 2988 460
rect 2969 445 2988 448
rect 2969 436 2991 445
rect 2942 426 2991 436
rect 2942 420 2972 426
rect 2991 421 2996 426
rect 2914 404 2988 420
rect 3006 412 3036 468
rect 3071 458 3279 468
rect 3314 464 3359 468
rect 3362 467 3363 468
rect 3378 467 3391 468
rect 3097 428 3286 458
rect 3112 425 3286 428
rect 3105 422 3286 425
rect 2914 402 2927 404
rect 2942 402 2976 404
rect 2914 386 2988 402
rect 3015 398 3028 412
rect 3043 398 3059 414
rect 3105 409 3116 422
rect 2898 364 2899 380
rect 2914 364 2927 386
rect 2942 364 2972 386
rect 3015 382 3077 398
rect 3105 391 3116 407
rect 3121 402 3131 422
rect 3141 402 3155 422
rect 3158 409 3167 422
rect 3183 409 3192 422
rect 3121 391 3155 402
rect 3158 391 3167 407
rect 3183 391 3192 407
rect 3199 402 3209 422
rect 3219 402 3233 422
rect 3234 409 3245 422
rect 3199 391 3233 402
rect 3234 391 3245 407
rect 3291 398 3307 414
rect 3314 412 3344 464
rect 3378 460 3379 467
rect 3363 452 3379 460
rect 3350 420 3363 439
rect 3378 420 3408 436
rect 3350 404 3424 420
rect 3350 402 3363 404
rect 3378 402 3412 404
rect 3015 380 3028 382
rect 3043 380 3077 382
rect 3015 364 3077 380
rect 3121 375 3137 378
rect 3199 375 3229 386
rect 3277 382 3323 398
rect 3350 386 3424 402
rect 3277 380 3311 382
rect 3276 364 3323 380
rect 3350 364 3363 386
rect 3378 364 3408 386
rect 3435 364 3436 380
rect 3451 364 3464 524
rect 3494 420 3507 524
rect 3552 502 3553 512
rect 3568 502 3581 512
rect 3552 498 3581 502
rect 3586 498 3616 524
rect 3634 510 3650 512
rect 3722 510 3775 524
rect 3723 508 3787 510
rect 3830 508 3845 524
rect 3894 521 3924 524
rect 3894 518 3930 521
rect 3860 510 3876 512
rect 3634 498 3649 502
rect 3552 496 3649 498
rect 3677 496 3845 508
rect 3861 498 3876 502
rect 3894 499 3933 518
rect 3952 512 3959 513
rect 3958 505 3959 512
rect 3942 502 3943 505
rect 3958 502 3971 505
rect 3894 498 3924 499
rect 3933 498 3939 499
rect 3942 498 3971 502
rect 3861 497 3971 498
rect 3861 496 3977 497
rect 3536 488 3587 496
rect 3536 476 3561 488
rect 3568 476 3587 488
rect 3618 488 3668 496
rect 3618 480 3634 488
rect 3641 486 3668 488
rect 3677 486 3898 496
rect 3641 476 3898 486
rect 3927 488 3977 496
rect 3927 479 3943 488
rect 3536 468 3587 476
rect 3634 468 3898 476
rect 3924 476 3943 479
rect 3950 476 3977 488
rect 3924 468 3977 476
rect 3552 460 3553 468
rect 3568 460 3581 468
rect 3552 452 3568 460
rect 3549 445 3568 448
rect 3549 436 3571 445
rect 3522 426 3571 436
rect 3522 420 3552 426
rect 3571 421 3576 426
rect 3494 404 3568 420
rect 3586 412 3616 468
rect 3651 458 3859 468
rect 3894 464 3939 468
rect 3942 467 3943 468
rect 3958 467 3971 468
rect 3677 428 3866 458
rect 3692 425 3866 428
rect 3685 422 3866 425
rect 3494 402 3507 404
rect 3522 402 3556 404
rect 3494 386 3568 402
rect 3595 398 3608 412
rect 3623 398 3639 414
rect 3685 409 3696 422
rect 3478 364 3479 380
rect 3494 364 3507 386
rect 3522 364 3552 386
rect 3595 382 3657 398
rect 3685 391 3696 407
rect 3701 402 3711 422
rect 3721 402 3735 422
rect 3738 409 3747 422
rect 3763 409 3772 422
rect 3701 391 3735 402
rect 3738 391 3747 407
rect 3763 391 3772 407
rect 3779 402 3789 422
rect 3799 402 3813 422
rect 3814 409 3825 422
rect 3779 391 3813 402
rect 3814 391 3825 407
rect 3871 398 3887 414
rect 3894 412 3924 464
rect 3958 460 3959 467
rect 3943 452 3959 460
rect 3930 420 3943 439
rect 3958 420 3988 436
rect 3930 404 4004 420
rect 3930 402 3943 404
rect 3958 402 3992 404
rect 3595 380 3608 382
rect 3623 380 3657 382
rect 3595 364 3657 380
rect 3701 375 3717 378
rect 3779 375 3809 386
rect 3857 382 3903 398
rect 3930 386 4004 402
rect 3857 380 3891 382
rect 3856 364 3903 380
rect 3930 364 3943 386
rect 3958 364 3988 386
rect 4015 364 4016 380
rect 4031 364 4044 524
rect 4074 420 4087 524
rect 4132 502 4133 512
rect 4148 502 4161 512
rect 4132 498 4161 502
rect 4166 498 4196 524
rect 4214 510 4230 512
rect 4302 510 4355 524
rect 4303 508 4367 510
rect 4410 508 4425 524
rect 4474 521 4504 524
rect 4611 523 6944 524
rect 4474 518 4510 521
rect 4440 510 4456 512
rect 4214 498 4229 502
rect 4132 496 4229 498
rect 4257 496 4425 508
rect 4441 498 4456 502
rect 4474 499 4513 518
rect 4532 512 4539 513
rect 4538 505 4539 512
rect 4522 502 4523 505
rect 4538 502 4551 505
rect 4474 498 4504 499
rect 4513 498 4519 499
rect 4522 498 4551 502
rect 4441 497 4551 498
rect 4441 496 4557 497
rect 4116 488 4167 496
rect 4116 476 4141 488
rect 4148 476 4167 488
rect 4198 488 4248 496
rect 4198 480 4214 488
rect 4221 486 4248 488
rect 4257 486 4478 496
rect 4221 476 4478 486
rect 4507 488 4557 496
rect 4507 479 4523 488
rect 4116 468 4167 476
rect 4214 468 4478 476
rect 4504 476 4523 479
rect 4530 476 4557 488
rect 4504 468 4557 476
rect 4132 460 4133 468
rect 4148 460 4161 468
rect 4132 452 4148 460
rect 4129 445 4148 448
rect 4129 436 4151 445
rect 4102 426 4151 436
rect 4102 420 4132 426
rect 4151 421 4156 426
rect 4074 404 4148 420
rect 4166 412 4196 468
rect 4231 458 4439 468
rect 4474 464 4519 468
rect 4522 467 4523 468
rect 4538 467 4551 468
rect 4257 428 4446 458
rect 4272 425 4446 428
rect 4265 422 4446 425
rect 4074 402 4087 404
rect 4102 402 4136 404
rect 4074 386 4148 402
rect 4175 398 4188 412
rect 4203 398 4219 414
rect 4265 409 4276 422
rect 4058 364 4059 380
rect 4074 364 4087 386
rect 4102 364 4132 386
rect 4175 382 4237 398
rect 4265 391 4276 407
rect 4281 402 4291 422
rect 4301 402 4315 422
rect 4318 409 4327 422
rect 4343 409 4352 422
rect 4281 391 4315 402
rect 4318 391 4327 407
rect 4343 391 4352 407
rect 4359 402 4369 422
rect 4379 402 4393 422
rect 4394 409 4405 422
rect 4359 391 4393 402
rect 4394 391 4405 407
rect 4451 398 4467 414
rect 4474 412 4504 464
rect 4538 460 4539 467
rect 4523 452 4539 460
rect 4510 420 4523 439
rect 4538 420 4568 436
rect 4510 404 4584 420
rect 4510 402 4523 404
rect 4538 402 4572 404
rect 4175 380 4188 382
rect 4203 380 4237 382
rect 4175 364 4237 380
rect 4281 375 4297 378
rect 4359 375 4389 386
rect 4437 382 4483 398
rect 4510 386 4584 402
rect 4437 380 4471 382
rect 4436 364 4483 380
rect 4510 364 4523 386
rect 4538 364 4568 386
rect 4595 364 4596 380
rect 4611 364 4624 523
rect 4654 419 4667 523
rect 4712 501 4713 511
rect 4733 509 4741 511
rect 4731 507 4741 509
rect 4728 501 4741 507
rect 4712 497 4741 501
rect 4746 497 4776 523
rect 4794 509 4810 511
rect 4882 509 4933 523
rect 4883 507 4947 509
rect 4990 507 5005 523
rect 5054 520 5084 523
rect 5054 517 5090 520
rect 5020 509 5036 511
rect 4794 497 4809 501
rect 4712 495 4809 497
rect 4837 495 5005 507
rect 5021 497 5036 501
rect 5054 498 5093 517
rect 5112 511 5119 512
rect 5118 504 5119 511
rect 5102 501 5103 504
rect 5118 501 5131 504
rect 5054 497 5084 498
rect 5093 497 5099 498
rect 5102 497 5131 501
rect 5021 496 5131 497
rect 5021 495 5137 496
rect 4696 487 4747 495
rect 4696 475 4721 487
rect 4728 475 4747 487
rect 4778 487 4828 495
rect 4778 479 4794 487
rect 4801 485 4828 487
rect 4837 485 5058 495
rect 4801 475 5058 485
rect 5087 487 5137 495
rect 5087 478 5103 487
rect 4696 467 4747 475
rect 4794 467 5058 475
rect 5084 475 5103 478
rect 5110 475 5137 487
rect 5084 467 5137 475
rect 4712 459 4713 467
rect 4728 459 4741 467
rect 4712 451 4728 459
rect 4709 444 4728 447
rect 4709 435 4731 444
rect 4682 425 4731 435
rect 4682 419 4712 425
rect 4731 420 4736 425
rect 4654 403 4728 419
rect 4746 411 4776 467
rect 4811 457 5019 467
rect 5054 463 5099 467
rect 5102 466 5103 467
rect 5118 466 5131 467
rect 4837 427 5026 457
rect 4852 424 5026 427
rect 4845 421 5026 424
rect 4654 401 4667 403
rect 4682 401 4716 403
rect 4654 385 4728 401
rect 4755 397 4768 411
rect 4783 397 4799 413
rect 4845 408 4856 421
rect -8 356 33 364
rect -8 330 7 356
rect 14 330 33 356
rect 97 352 159 364
rect 171 352 246 364
rect 304 352 379 364
rect 391 352 422 364
rect 428 352 463 364
rect 97 350 259 352
rect -8 322 33 330
rect 115 326 128 350
rect 143 348 158 350
rect -2 312 -1 322
rect 14 312 27 322
rect 42 312 72 326
rect 115 312 158 326
rect 182 323 189 330
rect 192 326 259 350
rect 291 350 463 352
rect 261 328 289 332
rect 291 328 371 350
rect 392 348 407 350
rect 261 326 371 328
rect 192 322 371 326
rect 165 312 195 322
rect 197 312 350 322
rect 358 312 388 322
rect 392 312 422 326
rect 450 312 463 350
rect 535 356 570 364
rect 535 330 536 356
rect 543 330 570 356
rect 478 312 508 326
rect 535 322 570 330
rect 572 356 613 364
rect 572 330 587 356
rect 594 330 613 356
rect 677 352 739 364
rect 751 352 826 364
rect 884 352 959 364
rect 971 352 1002 364
rect 1008 352 1043 364
rect 677 350 839 352
rect 572 322 613 330
rect 695 326 708 350
rect 723 348 738 350
rect 535 312 536 322
rect 551 312 564 322
rect 578 312 579 322
rect 594 312 607 322
rect 622 312 652 326
rect 695 312 738 326
rect 762 323 769 330
rect 772 326 839 350
rect 871 350 1043 352
rect 841 328 869 332
rect 871 328 951 350
rect 972 348 987 350
rect 841 326 951 328
rect 772 322 951 326
rect 745 312 775 322
rect 777 312 930 322
rect 938 312 968 322
rect 972 312 1002 326
rect 1030 312 1043 350
rect 1115 356 1150 364
rect 1115 330 1116 356
rect 1123 330 1150 356
rect 1058 312 1088 326
rect 1115 322 1150 330
rect 1152 356 1193 364
rect 1152 330 1167 356
rect 1174 330 1193 356
rect 1257 352 1319 364
rect 1331 352 1406 364
rect 1464 352 1539 364
rect 1551 352 1582 364
rect 1588 352 1623 364
rect 1257 350 1419 352
rect 1152 322 1193 330
rect 1275 326 1288 350
rect 1303 348 1318 350
rect 1115 312 1116 322
rect 1131 312 1144 322
rect 1158 312 1159 322
rect 1174 312 1187 322
rect 1202 312 1232 326
rect 1275 312 1318 326
rect 1342 323 1349 330
rect 1352 326 1419 350
rect 1451 350 1623 352
rect 1421 328 1449 332
rect 1451 328 1531 350
rect 1552 348 1567 350
rect 1421 326 1531 328
rect 1352 322 1531 326
rect 1325 312 1355 322
rect 1357 312 1510 322
rect 1518 312 1548 322
rect 1552 312 1582 326
rect 1610 312 1623 350
rect 1695 356 1730 364
rect 1695 330 1696 356
rect 1703 330 1730 356
rect 1638 312 1668 326
rect 1695 322 1730 330
rect 1732 356 1773 364
rect 1732 330 1747 356
rect 1754 330 1773 356
rect 1837 352 1899 364
rect 1911 352 1986 364
rect 2044 352 2119 364
rect 2131 352 2162 364
rect 2168 352 2203 364
rect 1837 350 1999 352
rect 1732 322 1773 330
rect 1855 326 1868 350
rect 1883 348 1898 350
rect 1695 312 1696 322
rect 1711 312 1724 322
rect 1738 312 1739 322
rect 1754 312 1767 322
rect 1782 312 1812 326
rect 1855 312 1898 326
rect 1922 323 1929 330
rect 1932 326 1999 350
rect 2031 350 2203 352
rect 2001 328 2029 332
rect 2031 328 2111 350
rect 2132 348 2147 350
rect 2001 326 2111 328
rect 1932 322 2111 326
rect 1905 312 1935 322
rect 1937 312 2090 322
rect 2098 312 2128 322
rect 2132 312 2162 326
rect 2190 312 2203 350
rect 2275 356 2310 364
rect 2275 330 2276 356
rect 2283 330 2310 356
rect 2218 312 2248 326
rect 2275 322 2310 330
rect 2312 356 2353 364
rect 2312 330 2327 356
rect 2334 330 2353 356
rect 2417 352 2479 364
rect 2491 352 2566 364
rect 2624 352 2699 364
rect 2711 352 2742 364
rect 2748 352 2783 364
rect 2417 350 2579 352
rect 2312 322 2353 330
rect 2435 326 2448 350
rect 2463 348 2478 350
rect 2275 312 2276 322
rect 2291 312 2304 322
rect 2318 312 2319 322
rect 2334 312 2347 322
rect 2362 312 2392 326
rect 2435 312 2478 326
rect 2502 323 2509 330
rect 2512 326 2579 350
rect 2611 350 2783 352
rect 2581 328 2609 332
rect 2611 328 2691 350
rect 2712 348 2727 350
rect 2581 326 2691 328
rect 2512 322 2691 326
rect 2485 312 2515 322
rect 2517 312 2670 322
rect 2678 312 2708 322
rect 2712 312 2742 326
rect 2770 312 2783 350
rect 2855 356 2890 364
rect 2855 330 2856 356
rect 2863 330 2890 356
rect 2798 312 2828 326
rect 2855 322 2890 330
rect 2892 356 2933 364
rect 2892 330 2907 356
rect 2914 330 2933 356
rect 2997 352 3059 364
rect 3071 352 3146 364
rect 3204 352 3279 364
rect 3291 352 3322 364
rect 3328 352 3363 364
rect 2997 350 3159 352
rect 2892 322 2933 330
rect 3015 326 3028 350
rect 3043 348 3058 350
rect 2855 312 2856 322
rect 2871 312 2884 322
rect 2898 312 2899 322
rect 2914 312 2927 322
rect 2942 312 2972 326
rect 3015 312 3058 326
rect 3082 323 3089 330
rect 3092 326 3159 350
rect 3191 350 3363 352
rect 3161 328 3189 332
rect 3191 328 3271 350
rect 3292 348 3307 350
rect 3161 326 3271 328
rect 3092 322 3271 326
rect 3065 312 3095 322
rect 3097 312 3250 322
rect 3258 312 3288 322
rect 3292 312 3322 326
rect 3350 312 3363 350
rect 3435 356 3470 364
rect 3435 330 3436 356
rect 3443 330 3470 356
rect 3378 312 3408 326
rect 3435 322 3470 330
rect 3472 356 3513 364
rect 3472 330 3487 356
rect 3494 330 3513 356
rect 3577 352 3639 364
rect 3651 352 3726 364
rect 3784 352 3859 364
rect 3871 352 3902 364
rect 3908 352 3943 364
rect 3577 350 3739 352
rect 3472 322 3513 330
rect 3595 326 3608 350
rect 3623 348 3638 350
rect 3435 312 3436 322
rect 3451 312 3464 322
rect 3478 312 3479 322
rect 3494 312 3507 322
rect 3522 312 3552 326
rect 3595 312 3638 326
rect 3662 323 3669 330
rect 3672 326 3739 350
rect 3771 350 3943 352
rect 3741 328 3769 332
rect 3771 328 3851 350
rect 3872 348 3887 350
rect 3741 326 3851 328
rect 3672 322 3851 326
rect 3645 312 3675 322
rect 3677 312 3830 322
rect 3838 312 3868 322
rect 3872 312 3902 326
rect 3930 312 3943 350
rect 4015 356 4050 364
rect 4015 330 4016 356
rect 4023 330 4050 356
rect 3958 312 3988 326
rect 4015 322 4050 330
rect 4052 356 4093 364
rect 4052 330 4067 356
rect 4074 330 4093 356
rect 4157 352 4219 364
rect 4231 352 4306 364
rect 4364 352 4439 364
rect 4451 352 4482 364
rect 4488 352 4523 364
rect 4157 350 4319 352
rect 4052 322 4093 330
rect 4175 326 4188 350
rect 4203 348 4218 350
rect 4015 312 4016 322
rect 4031 312 4044 322
rect 4058 312 4059 322
rect 4074 312 4087 322
rect 4102 312 4132 326
rect 4175 312 4218 326
rect 4242 323 4249 330
rect 4252 326 4319 350
rect 4351 350 4523 352
rect 4321 328 4349 332
rect 4351 328 4431 350
rect 4452 348 4467 350
rect 4321 326 4431 328
rect 4252 322 4431 326
rect 4225 312 4255 322
rect 4257 312 4410 322
rect 4418 312 4448 322
rect 4452 312 4482 326
rect 4510 312 4523 350
rect 4595 356 4630 364
rect 4638 363 4639 379
rect 4654 363 4667 385
rect 4682 363 4712 385
rect 4755 381 4817 397
rect 4845 390 4856 406
rect 4861 401 4871 421
rect 4881 401 4895 421
rect 4898 408 4907 421
rect 4923 408 4932 421
rect 4861 390 4895 401
rect 4898 390 4907 406
rect 4923 390 4932 406
rect 4939 401 4949 421
rect 4959 401 4973 421
rect 4974 408 4985 421
rect 4939 390 4973 401
rect 4974 390 4985 406
rect 5031 397 5047 413
rect 5054 411 5084 463
rect 5118 459 5119 466
rect 5103 451 5119 459
rect 5090 419 5103 438
rect 5118 419 5148 435
rect 5090 403 5164 419
rect 5090 401 5103 403
rect 5118 401 5152 403
rect 4755 379 4768 381
rect 4783 379 4817 381
rect 4755 363 4817 379
rect 4861 374 4877 377
rect 4939 374 4969 385
rect 5017 381 5063 397
rect 5090 385 5164 401
rect 5017 379 5051 381
rect 5016 363 5063 379
rect 5090 363 5103 385
rect 5118 363 5148 385
rect 5175 363 5176 379
rect 5191 363 5204 523
rect 5234 419 5247 523
rect 5292 501 5293 511
rect 5313 509 5321 511
rect 5311 507 5321 509
rect 5308 501 5321 507
rect 5292 497 5321 501
rect 5326 497 5356 523
rect 5374 509 5390 511
rect 5462 509 5513 523
rect 5463 507 5527 509
rect 5570 507 5585 523
rect 5634 520 5664 523
rect 5634 517 5670 520
rect 5600 509 5616 511
rect 5374 497 5389 501
rect 5292 495 5389 497
rect 5417 495 5585 507
rect 5601 497 5616 501
rect 5634 498 5673 517
rect 5692 511 5699 512
rect 5698 504 5699 511
rect 5682 501 5683 504
rect 5698 501 5711 504
rect 5634 497 5664 498
rect 5673 497 5679 498
rect 5682 497 5711 501
rect 5601 496 5711 497
rect 5601 495 5717 496
rect 5276 487 5327 495
rect 5276 475 5301 487
rect 5308 475 5327 487
rect 5358 487 5408 495
rect 5358 479 5374 487
rect 5381 485 5408 487
rect 5417 485 5638 495
rect 5381 475 5638 485
rect 5667 487 5717 495
rect 5667 478 5683 487
rect 5276 467 5327 475
rect 5374 467 5638 475
rect 5664 475 5683 478
rect 5690 475 5717 487
rect 5664 467 5717 475
rect 5292 459 5293 467
rect 5308 459 5321 467
rect 5292 451 5308 459
rect 5289 444 5308 447
rect 5289 435 5311 444
rect 5262 425 5311 435
rect 5262 419 5292 425
rect 5311 420 5316 425
rect 5234 403 5308 419
rect 5326 411 5356 467
rect 5391 457 5599 467
rect 5634 463 5679 467
rect 5682 466 5683 467
rect 5698 466 5711 467
rect 5417 427 5606 457
rect 5432 424 5606 427
rect 5425 421 5606 424
rect 5234 401 5247 403
rect 5262 401 5296 403
rect 5234 385 5308 401
rect 5335 397 5348 411
rect 5363 397 5379 413
rect 5425 408 5436 421
rect 5218 363 5219 379
rect 5234 363 5247 385
rect 5262 363 5292 385
rect 5335 381 5397 397
rect 5425 390 5436 406
rect 5441 401 5451 421
rect 5461 401 5475 421
rect 5478 408 5487 421
rect 5503 408 5512 421
rect 5441 390 5475 401
rect 5478 390 5487 406
rect 5503 390 5512 406
rect 5519 401 5529 421
rect 5539 401 5553 421
rect 5554 408 5565 421
rect 5519 390 5553 401
rect 5554 390 5565 406
rect 5611 397 5627 413
rect 5634 411 5664 463
rect 5698 459 5699 466
rect 5683 451 5699 459
rect 5670 419 5683 438
rect 5698 419 5728 435
rect 5670 403 5744 419
rect 5670 401 5683 403
rect 5698 401 5732 403
rect 5335 379 5348 381
rect 5363 379 5397 381
rect 5335 363 5397 379
rect 5441 374 5457 377
rect 5519 374 5549 385
rect 5597 381 5643 397
rect 5670 385 5744 401
rect 5597 379 5631 381
rect 5596 363 5643 379
rect 5670 363 5683 385
rect 5698 363 5728 385
rect 5755 363 5756 379
rect 5771 363 5784 523
rect 5814 419 5827 523
rect 5872 501 5873 511
rect 5893 509 5901 511
rect 5891 507 5901 509
rect 5888 501 5901 507
rect 5872 497 5901 501
rect 5906 497 5936 523
rect 5954 509 5970 511
rect 6042 509 6093 523
rect 6043 507 6107 509
rect 6150 507 6165 523
rect 6214 520 6244 523
rect 6214 517 6250 520
rect 6180 509 6196 511
rect 5954 497 5969 501
rect 5872 495 5969 497
rect 5997 495 6165 507
rect 6181 497 6196 501
rect 6214 498 6253 517
rect 6272 511 6279 512
rect 6278 504 6279 511
rect 6262 501 6263 504
rect 6278 501 6291 504
rect 6214 497 6244 498
rect 6253 497 6259 498
rect 6262 497 6291 501
rect 6181 496 6291 497
rect 6181 495 6297 496
rect 5856 487 5907 495
rect 5856 475 5881 487
rect 5888 475 5907 487
rect 5938 487 5988 495
rect 5938 479 5954 487
rect 5961 485 5988 487
rect 5997 485 6218 495
rect 5961 475 6218 485
rect 6247 487 6297 495
rect 6247 478 6263 487
rect 5856 467 5907 475
rect 5954 467 6218 475
rect 6244 475 6263 478
rect 6270 475 6297 487
rect 6244 467 6297 475
rect 5872 459 5873 467
rect 5888 459 5901 467
rect 5872 451 5888 459
rect 5869 444 5888 447
rect 5869 435 5891 444
rect 5842 425 5891 435
rect 5842 419 5872 425
rect 5891 420 5896 425
rect 5814 403 5888 419
rect 5906 411 5936 467
rect 5971 457 6179 467
rect 6214 463 6259 467
rect 6262 466 6263 467
rect 6278 466 6291 467
rect 5997 427 6186 457
rect 6012 424 6186 427
rect 6005 421 6186 424
rect 5814 401 5827 403
rect 5842 401 5876 403
rect 5814 385 5888 401
rect 5915 397 5928 411
rect 5943 397 5959 413
rect 6005 408 6016 421
rect 5798 363 5799 379
rect 5814 363 5827 385
rect 5842 363 5872 385
rect 5915 381 5977 397
rect 6005 390 6016 406
rect 6021 401 6031 421
rect 6041 401 6055 421
rect 6058 408 6067 421
rect 6083 408 6092 421
rect 6021 390 6055 401
rect 6058 390 6067 406
rect 6083 390 6092 406
rect 6099 401 6109 421
rect 6119 401 6133 421
rect 6134 408 6145 421
rect 6099 390 6133 401
rect 6134 390 6145 406
rect 6191 397 6207 413
rect 6214 411 6244 463
rect 6278 459 6279 466
rect 6263 451 6279 459
rect 6250 419 6263 438
rect 6278 419 6308 435
rect 6250 403 6324 419
rect 6250 401 6263 403
rect 6278 401 6312 403
rect 5915 379 5928 381
rect 5943 379 5977 381
rect 5915 363 5977 379
rect 6021 374 6037 377
rect 6099 374 6129 385
rect 6177 381 6223 397
rect 6250 385 6324 401
rect 6177 379 6211 381
rect 6176 363 6223 379
rect 6250 363 6263 385
rect 6278 363 6308 385
rect 6335 363 6336 379
rect 6351 363 6364 523
rect 6394 419 6407 523
rect 6452 501 6453 511
rect 6473 509 6481 511
rect 6471 507 6481 509
rect 6468 501 6481 507
rect 6452 497 6481 501
rect 6486 497 6516 523
rect 6534 509 6550 511
rect 6622 509 6673 523
rect 6623 507 6687 509
rect 6730 507 6745 523
rect 6794 520 6824 523
rect 6794 517 6830 520
rect 6760 509 6776 511
rect 6534 497 6549 501
rect 6452 495 6549 497
rect 6577 495 6745 507
rect 6761 497 6776 501
rect 6794 498 6833 517
rect 6852 511 6859 512
rect 6858 504 6859 511
rect 6842 501 6843 504
rect 6858 501 6871 504
rect 6794 497 6824 498
rect 6833 497 6839 498
rect 6842 497 6871 501
rect 6761 496 6871 497
rect 6761 495 6877 496
rect 6436 487 6487 495
rect 6436 475 6461 487
rect 6468 475 6487 487
rect 6518 487 6568 495
rect 6518 479 6534 487
rect 6541 485 6568 487
rect 6577 485 6798 495
rect 6541 475 6798 485
rect 6827 487 6877 495
rect 6827 478 6843 487
rect 6436 467 6487 475
rect 6534 467 6798 475
rect 6824 475 6843 478
rect 6850 475 6877 487
rect 6824 467 6877 475
rect 6452 459 6453 467
rect 6468 459 6481 467
rect 6452 451 6468 459
rect 6449 444 6468 447
rect 6449 435 6471 444
rect 6422 425 6471 435
rect 6422 419 6452 425
rect 6471 420 6476 425
rect 6394 403 6468 419
rect 6486 411 6516 467
rect 6551 457 6759 467
rect 6794 463 6839 467
rect 6842 466 6843 467
rect 6858 466 6871 467
rect 6577 427 6766 457
rect 6592 424 6766 427
rect 6585 421 6766 424
rect 6394 401 6407 403
rect 6422 401 6456 403
rect 6394 385 6468 401
rect 6495 397 6508 411
rect 6523 397 6539 413
rect 6585 408 6596 421
rect 6378 363 6379 379
rect 6394 363 6407 385
rect 6422 363 6452 385
rect 6495 381 6557 397
rect 6585 390 6596 406
rect 6601 401 6611 421
rect 6621 401 6635 421
rect 6638 408 6647 421
rect 6663 408 6672 421
rect 6601 390 6635 401
rect 6638 390 6647 406
rect 6663 390 6672 406
rect 6679 401 6689 421
rect 6699 401 6713 421
rect 6714 408 6725 421
rect 6679 390 6713 401
rect 6714 390 6725 406
rect 6771 397 6787 413
rect 6794 411 6824 463
rect 6858 459 6859 466
rect 6843 451 6859 459
rect 6830 419 6843 438
rect 6858 419 6888 435
rect 6830 403 6904 419
rect 6830 401 6843 403
rect 6858 401 6892 403
rect 6495 379 6508 381
rect 6523 379 6557 381
rect 6495 363 6557 379
rect 6601 374 6617 377
rect 6679 374 6709 385
rect 6757 381 6803 397
rect 6830 385 6904 401
rect 6757 379 6791 381
rect 6756 363 6803 379
rect 6830 363 6843 385
rect 6858 363 6888 385
rect 6915 363 6916 379
rect 6931 363 6944 523
rect 4595 330 4596 356
rect 4603 330 4630 356
rect 4538 312 4568 326
rect 4595 322 4630 330
rect 4632 355 4673 363
rect 4632 329 4647 355
rect 4654 329 4673 355
rect 4737 351 4799 363
rect 4811 351 4886 363
rect 4944 351 5019 363
rect 5031 351 5062 363
rect 5068 351 5103 363
rect 4737 349 4899 351
rect 4595 312 4596 322
rect 4611 312 4624 322
rect 4632 321 4673 329
rect 4755 325 4768 349
rect 4783 347 4798 349
rect 4832 331 4899 349
rect 4931 349 5103 351
rect 4931 331 5011 349
rect 5032 347 5047 349
rect -2 311 4624 312
rect 4638 311 4639 321
rect 4654 311 4667 321
rect 4682 311 4712 325
rect 4755 311 4798 325
rect 4822 322 4829 329
rect 4832 321 5011 331
rect 4805 311 4835 321
rect 4837 311 4990 321
rect 4998 311 5028 321
rect 5032 311 5062 325
rect 5090 311 5103 349
rect 5175 355 5210 363
rect 5175 329 5176 355
rect 5183 329 5210 355
rect 5118 311 5148 325
rect 5175 321 5210 329
rect 5212 355 5253 363
rect 5212 329 5227 355
rect 5234 329 5253 355
rect 5317 351 5379 363
rect 5391 351 5466 363
rect 5524 351 5599 363
rect 5611 351 5642 363
rect 5648 351 5683 363
rect 5317 349 5479 351
rect 5212 321 5253 329
rect 5335 325 5348 349
rect 5363 347 5378 349
rect 5412 331 5479 349
rect 5511 349 5683 351
rect 5511 331 5591 349
rect 5612 347 5627 349
rect 5175 311 5176 321
rect 5191 311 5204 321
rect 5218 311 5219 321
rect 5234 311 5247 321
rect 5262 311 5292 325
rect 5335 311 5378 325
rect 5402 322 5409 329
rect 5412 321 5591 331
rect 5385 311 5415 321
rect 5417 311 5570 321
rect 5578 311 5608 321
rect 5612 311 5642 325
rect 5670 311 5683 349
rect 5755 355 5790 363
rect 5755 329 5756 355
rect 5763 329 5790 355
rect 5698 311 5728 325
rect 5755 321 5790 329
rect 5792 355 5833 363
rect 5792 329 5807 355
rect 5814 329 5833 355
rect 5897 351 5959 363
rect 5971 351 6046 363
rect 6104 351 6179 363
rect 6191 351 6222 363
rect 6228 351 6263 363
rect 5897 349 6059 351
rect 5792 321 5833 329
rect 5915 325 5928 349
rect 5943 347 5958 349
rect 5992 331 6059 349
rect 6091 349 6263 351
rect 6091 331 6171 349
rect 6192 347 6207 349
rect 5755 311 5756 321
rect 5771 311 5784 321
rect 5798 311 5799 321
rect 5814 311 5827 321
rect 5842 311 5872 325
rect 5915 311 5958 325
rect 5982 322 5989 329
rect 5992 321 6171 331
rect 5965 311 5995 321
rect 5997 311 6150 321
rect 6158 311 6188 321
rect 6192 311 6222 325
rect 6250 311 6263 349
rect 6335 355 6370 363
rect 6335 329 6336 355
rect 6343 329 6370 355
rect 6278 311 6308 325
rect 6335 321 6370 329
rect 6372 355 6413 363
rect 6372 329 6387 355
rect 6394 329 6413 355
rect 6477 351 6539 363
rect 6551 351 6626 363
rect 6684 351 6759 363
rect 6771 351 6802 363
rect 6808 351 6843 363
rect 6477 349 6639 351
rect 6372 321 6413 329
rect 6495 325 6508 349
rect 6523 347 6538 349
rect 6572 331 6639 349
rect 6671 349 6843 351
rect 6671 331 6751 349
rect 6772 347 6787 349
rect 6335 311 6336 321
rect 6351 311 6364 321
rect 6378 311 6379 321
rect 6394 311 6407 321
rect 6422 311 6452 325
rect 6495 311 6538 325
rect 6562 322 6569 329
rect 6572 321 6751 331
rect 6545 311 6575 321
rect 6577 311 6730 321
rect 6738 311 6768 321
rect 6772 311 6802 325
rect 6830 311 6843 349
rect 6915 355 6950 363
rect 6915 329 6916 355
rect 6923 329 6950 355
rect 6858 311 6888 325
rect 6915 321 6950 329
rect 6915 311 6916 321
rect 6931 311 6944 321
rect -2 306 6944 311
rect -1 298 6944 306
rect 14 268 27 298
rect 42 280 72 298
rect 115 284 129 298
rect 165 284 385 298
rect 116 282 129 284
rect 82 270 97 282
rect 79 268 101 270
rect 106 268 136 282
rect 197 280 350 284
rect 179 268 371 280
rect 414 268 444 282
rect 450 268 463 298
rect 478 280 508 298
rect 551 268 564 298
rect 594 268 607 298
rect 622 280 652 298
rect 695 284 709 298
rect 745 284 965 298
rect 696 282 709 284
rect 662 270 677 282
rect 659 268 681 270
rect 686 268 716 282
rect 777 280 930 284
rect 759 268 951 280
rect 994 268 1024 282
rect 1030 268 1043 298
rect 1058 280 1088 298
rect 1131 268 1144 298
rect 1174 268 1187 298
rect 1202 280 1232 298
rect 1275 284 1289 298
rect 1325 284 1545 298
rect 1276 282 1289 284
rect 1242 270 1257 282
rect 1239 268 1261 270
rect 1266 268 1296 282
rect 1357 280 1510 284
rect 1339 268 1531 280
rect 1574 268 1604 282
rect 1610 268 1623 298
rect 1638 280 1668 298
rect 1711 268 1724 298
rect 1754 268 1767 298
rect 1782 280 1812 298
rect 1855 284 1869 298
rect 1905 284 2125 298
rect 1856 282 1869 284
rect 1822 270 1837 282
rect 1819 268 1841 270
rect 1846 268 1876 282
rect 1937 280 2090 284
rect 1919 268 2111 280
rect 2154 268 2184 282
rect 2190 268 2203 298
rect 2218 280 2248 298
rect 2291 268 2304 298
rect 2334 268 2347 298
rect 2362 280 2392 298
rect 2435 284 2449 298
rect 2485 284 2705 298
rect 2436 282 2449 284
rect 2402 270 2417 282
rect 2399 268 2421 270
rect 2426 268 2456 282
rect 2517 280 2670 284
rect 2499 268 2691 280
rect 2734 268 2764 282
rect 2770 268 2783 298
rect 2798 280 2828 298
rect 2871 268 2884 298
rect 2914 268 2927 298
rect 2942 280 2972 298
rect 3015 284 3029 298
rect 3065 284 3285 298
rect 3016 282 3029 284
rect 2982 270 2997 282
rect 2979 268 3001 270
rect 3006 268 3036 282
rect 3097 280 3250 284
rect 3079 268 3271 280
rect 3314 268 3344 282
rect 3350 268 3363 298
rect 3378 280 3408 298
rect 3451 268 3464 298
rect 3494 268 3507 298
rect 3522 280 3552 298
rect 3595 284 3609 298
rect 3645 284 3865 298
rect 3596 282 3609 284
rect 3562 270 3577 282
rect 3559 268 3581 270
rect 3586 268 3616 282
rect 3677 280 3830 284
rect 3659 268 3851 280
rect 3894 268 3924 282
rect 3930 268 3943 298
rect 3958 280 3988 298
rect 4031 268 4044 298
rect 4074 268 4087 298
rect 4102 280 4132 298
rect 4175 284 4189 298
rect 4225 284 4445 298
rect 4176 282 4189 284
rect 4142 270 4157 282
rect 4139 268 4161 270
rect 4166 268 4196 282
rect 4257 280 4410 284
rect 4239 268 4431 280
rect 4474 268 4504 282
rect 4510 268 4523 298
rect 4538 280 4568 298
rect 4611 297 6944 298
rect 4611 268 4624 297
rect -1 267 4624 268
rect 4654 267 4667 297
rect 4682 279 4712 297
rect 4755 283 4769 297
rect 4805 283 5025 297
rect 4756 281 4769 283
rect 4722 269 4737 281
rect 4719 267 4741 269
rect 4746 267 4776 281
rect 4837 279 4990 283
rect 4819 267 5011 279
rect 5054 267 5084 281
rect 5090 267 5103 297
rect 5118 279 5148 297
rect 5191 267 5204 297
rect 5234 267 5247 297
rect 5262 279 5292 297
rect 5335 283 5349 297
rect 5385 283 5605 297
rect 5336 281 5349 283
rect 5302 269 5317 281
rect 5299 267 5321 269
rect 5326 267 5356 281
rect 5417 279 5570 283
rect 5399 267 5591 279
rect 5634 267 5664 281
rect 5670 267 5683 297
rect 5698 279 5728 297
rect 5771 267 5784 297
rect 5814 267 5827 297
rect 5842 279 5872 297
rect 5915 283 5929 297
rect 5965 283 6185 297
rect 5916 281 5929 283
rect 5882 269 5897 281
rect 5879 267 5901 269
rect 5906 267 5936 281
rect 5997 279 6150 283
rect 5979 267 6171 279
rect 6214 267 6244 281
rect 6250 267 6263 297
rect 6278 279 6308 297
rect 6351 267 6364 297
rect 6394 267 6407 297
rect 6422 279 6452 297
rect 6495 283 6509 297
rect 6545 283 6765 297
rect 6496 281 6509 283
rect 6462 269 6477 281
rect 6459 267 6481 269
rect 6486 267 6516 281
rect 6577 279 6730 283
rect 6559 267 6751 279
rect 6794 267 6824 281
rect 6830 267 6843 297
rect 6858 279 6888 297
rect 6931 267 6944 297
rect -1 254 6944 267
rect 14 150 27 254
rect 72 232 73 242
rect 88 232 101 242
rect 72 228 101 232
rect 106 228 136 254
rect 154 240 170 242
rect 242 240 295 254
rect 243 238 307 240
rect 350 238 365 254
rect 414 251 444 254
rect 414 248 450 251
rect 380 240 396 242
rect 154 228 169 232
rect 72 226 169 228
rect 197 226 365 238
rect 381 228 396 232
rect 414 229 453 248
rect 472 242 479 243
rect 478 235 479 242
rect 462 232 463 235
rect 478 232 491 235
rect 414 228 444 229
rect 453 228 459 229
rect 462 228 491 232
rect 381 227 491 228
rect 381 226 497 227
rect 56 218 107 226
rect 56 206 81 218
rect 88 206 107 218
rect 138 218 188 226
rect 138 210 154 218
rect 161 216 188 218
rect 197 216 418 226
rect 161 206 418 216
rect 447 218 497 226
rect 447 209 463 218
rect 56 198 107 206
rect 154 198 418 206
rect 444 206 463 209
rect 470 206 497 218
rect 444 198 497 206
rect 72 190 73 198
rect 88 190 101 198
rect 72 182 88 190
rect 69 175 88 178
rect 69 166 91 175
rect 42 156 91 166
rect 42 150 72 156
rect 91 151 96 156
rect 14 134 88 150
rect 106 142 136 198
rect 171 188 379 198
rect 414 194 459 198
rect 462 197 463 198
rect 478 197 491 198
rect 197 158 386 188
rect 212 155 386 158
rect 205 152 386 155
rect 14 132 27 134
rect 42 132 76 134
rect 14 116 88 132
rect 115 128 128 142
rect 143 128 159 144
rect 205 139 216 152
rect -2 94 -1 110
rect 14 94 27 116
rect 42 94 72 116
rect 115 112 177 128
rect 205 121 216 137
rect 221 132 231 152
rect 241 132 255 152
rect 258 139 267 152
rect 283 139 292 152
rect 221 121 255 132
rect 258 121 266 137
rect 283 121 292 137
rect 299 132 309 152
rect 319 132 333 152
rect 334 139 345 152
rect 299 121 333 132
rect 334 121 345 137
rect 391 128 407 144
rect 414 142 444 194
rect 478 190 479 197
rect 463 182 479 190
rect 450 150 463 169
rect 478 150 508 166
rect 450 134 524 150
rect 450 132 463 134
rect 478 132 512 134
rect 115 110 128 112
rect 143 110 177 112
rect 115 94 177 110
rect 221 105 234 108
rect 299 105 329 116
rect 377 112 423 128
rect 450 116 524 132
rect 377 110 411 112
rect 376 94 423 110
rect 450 94 463 116
rect 478 94 508 116
rect 535 94 536 110
rect 551 94 564 254
rect 594 150 607 254
rect 652 232 653 242
rect 668 232 681 242
rect 652 228 681 232
rect 686 228 716 254
rect 734 240 750 242
rect 822 240 875 254
rect 823 238 887 240
rect 930 238 945 254
rect 994 251 1024 254
rect 994 248 1030 251
rect 960 240 976 242
rect 734 228 749 232
rect 652 226 749 228
rect 777 226 945 238
rect 961 228 976 232
rect 994 229 1033 248
rect 1052 242 1059 243
rect 1058 235 1059 242
rect 1042 232 1043 235
rect 1058 232 1071 235
rect 994 228 1024 229
rect 1033 228 1039 229
rect 1042 228 1071 232
rect 961 227 1071 228
rect 961 226 1077 227
rect 636 218 687 226
rect 636 206 661 218
rect 668 206 687 218
rect 718 218 768 226
rect 718 210 734 218
rect 741 216 768 218
rect 777 216 998 226
rect 741 206 998 216
rect 1027 218 1077 226
rect 1027 209 1043 218
rect 636 198 687 206
rect 734 198 998 206
rect 1024 206 1043 209
rect 1050 206 1077 218
rect 1024 198 1077 206
rect 652 190 653 198
rect 668 190 681 198
rect 652 182 668 190
rect 649 175 668 178
rect 649 166 671 175
rect 622 156 671 166
rect 622 150 652 156
rect 671 151 676 156
rect 594 134 668 150
rect 686 142 716 198
rect 751 188 959 198
rect 994 194 1039 198
rect 1042 197 1043 198
rect 1058 197 1071 198
rect 777 158 966 188
rect 792 155 966 158
rect 785 152 966 155
rect 594 132 607 134
rect 622 132 656 134
rect 594 116 668 132
rect 695 128 708 142
rect 723 128 739 144
rect 785 139 796 152
rect 578 94 579 110
rect 594 94 607 116
rect 622 94 652 116
rect 695 112 757 128
rect 785 121 796 137
rect 801 132 811 152
rect 821 132 835 152
rect 838 139 847 152
rect 863 139 872 152
rect 801 121 835 132
rect 838 121 846 137
rect 863 121 872 137
rect 879 132 889 152
rect 899 132 913 152
rect 914 139 925 152
rect 879 121 913 132
rect 914 121 925 137
rect 971 128 987 144
rect 994 142 1024 194
rect 1058 190 1059 197
rect 1043 182 1059 190
rect 1030 150 1043 169
rect 1058 150 1088 166
rect 1030 134 1104 150
rect 1030 132 1043 134
rect 1058 132 1092 134
rect 695 110 708 112
rect 723 110 757 112
rect 695 94 757 110
rect 801 105 814 108
rect 879 105 909 116
rect 957 112 1003 128
rect 1030 116 1104 132
rect 957 110 991 112
rect 956 94 1003 110
rect 1030 94 1043 116
rect 1058 94 1088 116
rect 1115 94 1116 110
rect 1131 94 1144 254
rect 1174 150 1187 254
rect 1232 232 1233 242
rect 1248 232 1261 242
rect 1232 228 1261 232
rect 1266 228 1296 254
rect 1314 240 1330 242
rect 1402 240 1455 254
rect 1403 238 1467 240
rect 1510 238 1525 254
rect 1574 251 1604 254
rect 1574 248 1610 251
rect 1540 240 1556 242
rect 1314 228 1329 232
rect 1232 226 1329 228
rect 1357 226 1525 238
rect 1541 228 1556 232
rect 1574 229 1613 248
rect 1632 242 1639 243
rect 1638 235 1639 242
rect 1622 232 1623 235
rect 1638 232 1651 235
rect 1574 228 1604 229
rect 1613 228 1619 229
rect 1622 228 1651 232
rect 1541 227 1651 228
rect 1541 226 1657 227
rect 1216 218 1267 226
rect 1216 206 1241 218
rect 1248 206 1267 218
rect 1298 218 1348 226
rect 1298 210 1314 218
rect 1321 216 1348 218
rect 1357 216 1578 226
rect 1321 206 1578 216
rect 1607 218 1657 226
rect 1607 209 1623 218
rect 1216 198 1267 206
rect 1314 198 1578 206
rect 1604 206 1623 209
rect 1630 206 1657 218
rect 1604 198 1657 206
rect 1232 190 1233 198
rect 1248 190 1261 198
rect 1232 182 1248 190
rect 1229 175 1248 178
rect 1229 166 1251 175
rect 1202 156 1251 166
rect 1202 150 1232 156
rect 1251 151 1256 156
rect 1174 134 1248 150
rect 1266 142 1296 198
rect 1331 188 1539 198
rect 1574 194 1619 198
rect 1622 197 1623 198
rect 1638 197 1651 198
rect 1357 158 1546 188
rect 1372 155 1546 158
rect 1365 152 1546 155
rect 1174 132 1187 134
rect 1202 132 1236 134
rect 1174 116 1248 132
rect 1275 128 1288 142
rect 1303 128 1319 144
rect 1365 139 1376 152
rect 1158 94 1159 110
rect 1174 94 1187 116
rect 1202 94 1232 116
rect 1275 112 1337 128
rect 1365 121 1376 137
rect 1381 132 1391 152
rect 1401 132 1415 152
rect 1418 139 1427 152
rect 1443 139 1452 152
rect 1381 121 1415 132
rect 1418 121 1426 137
rect 1443 121 1452 137
rect 1459 132 1469 152
rect 1479 132 1493 152
rect 1494 139 1505 152
rect 1459 121 1493 132
rect 1494 121 1505 137
rect 1551 128 1567 144
rect 1574 142 1604 194
rect 1638 190 1639 197
rect 1623 182 1639 190
rect 1610 150 1623 169
rect 1638 150 1668 166
rect 1610 134 1684 150
rect 1610 132 1623 134
rect 1638 132 1672 134
rect 1275 110 1288 112
rect 1303 110 1337 112
rect 1275 94 1337 110
rect 1381 105 1394 108
rect 1459 105 1489 116
rect 1537 112 1583 128
rect 1610 116 1684 132
rect 1537 110 1571 112
rect 1536 94 1583 110
rect 1610 94 1623 116
rect 1638 94 1668 116
rect 1695 94 1696 110
rect 1711 94 1724 254
rect 1754 150 1767 254
rect 1812 232 1813 242
rect 1828 232 1841 242
rect 1812 228 1841 232
rect 1846 228 1876 254
rect 1894 240 1910 242
rect 1982 240 2035 254
rect 1983 238 2047 240
rect 2090 238 2105 254
rect 2154 251 2184 254
rect 2154 248 2190 251
rect 2120 240 2136 242
rect 1894 228 1909 232
rect 1812 226 1909 228
rect 1937 226 2105 238
rect 2121 228 2136 232
rect 2154 229 2193 248
rect 2212 242 2219 243
rect 2218 235 2219 242
rect 2202 232 2203 235
rect 2218 232 2231 235
rect 2154 228 2184 229
rect 2193 228 2199 229
rect 2202 228 2231 232
rect 2121 227 2231 228
rect 2121 226 2237 227
rect 1796 218 1847 226
rect 1796 206 1821 218
rect 1828 206 1847 218
rect 1878 218 1928 226
rect 1878 210 1894 218
rect 1901 216 1928 218
rect 1937 216 2158 226
rect 1901 206 2158 216
rect 2187 218 2237 226
rect 2187 209 2203 218
rect 1796 198 1847 206
rect 1894 198 2158 206
rect 2184 206 2203 209
rect 2210 206 2237 218
rect 2184 198 2237 206
rect 1812 190 1813 198
rect 1828 190 1841 198
rect 1812 182 1828 190
rect 1809 175 1828 178
rect 1809 166 1831 175
rect 1782 156 1831 166
rect 1782 150 1812 156
rect 1831 151 1836 156
rect 1754 134 1828 150
rect 1846 142 1876 198
rect 1911 188 2119 198
rect 2154 194 2199 198
rect 2202 197 2203 198
rect 2218 197 2231 198
rect 1937 158 2126 188
rect 1952 155 2126 158
rect 1945 152 2126 155
rect 1754 132 1767 134
rect 1782 132 1816 134
rect 1754 116 1828 132
rect 1855 128 1868 142
rect 1883 128 1899 144
rect 1945 139 1956 152
rect 1738 94 1739 110
rect 1754 94 1767 116
rect 1782 94 1812 116
rect 1855 112 1917 128
rect 1945 121 1956 137
rect 1961 132 1971 152
rect 1981 132 1995 152
rect 1998 139 2007 152
rect 2023 139 2032 152
rect 1961 121 1995 132
rect 1998 121 2006 137
rect 2023 121 2032 137
rect 2039 132 2049 152
rect 2059 132 2073 152
rect 2074 139 2085 152
rect 2039 121 2073 132
rect 2074 121 2085 137
rect 2131 128 2147 144
rect 2154 142 2184 194
rect 2218 190 2219 197
rect 2203 182 2219 190
rect 2190 150 2203 169
rect 2218 150 2248 166
rect 2190 134 2264 150
rect 2190 132 2203 134
rect 2218 132 2252 134
rect 1855 110 1868 112
rect 1883 110 1917 112
rect 1855 94 1917 110
rect 1961 105 1974 108
rect 2039 105 2069 116
rect 2117 112 2163 128
rect 2190 116 2264 132
rect 2117 110 2151 112
rect 2116 94 2163 110
rect 2190 94 2203 116
rect 2218 94 2248 116
rect 2275 94 2276 110
rect 2291 94 2304 254
rect 2334 150 2347 254
rect 2392 232 2393 242
rect 2408 232 2421 242
rect 2392 228 2421 232
rect 2426 228 2456 254
rect 2474 240 2490 242
rect 2562 240 2615 254
rect 2563 238 2627 240
rect 2670 238 2685 254
rect 2734 251 2764 254
rect 2734 248 2770 251
rect 2700 240 2716 242
rect 2474 228 2489 232
rect 2392 226 2489 228
rect 2517 226 2685 238
rect 2701 228 2716 232
rect 2734 229 2773 248
rect 2792 242 2799 243
rect 2798 235 2799 242
rect 2782 232 2783 235
rect 2798 232 2811 235
rect 2734 228 2764 229
rect 2773 228 2779 229
rect 2782 228 2811 232
rect 2701 227 2811 228
rect 2701 226 2817 227
rect 2376 218 2427 226
rect 2376 206 2401 218
rect 2408 206 2427 218
rect 2458 218 2508 226
rect 2458 210 2474 218
rect 2481 216 2508 218
rect 2517 216 2738 226
rect 2481 206 2738 216
rect 2767 218 2817 226
rect 2767 209 2783 218
rect 2376 198 2427 206
rect 2474 198 2738 206
rect 2764 206 2783 209
rect 2790 206 2817 218
rect 2764 198 2817 206
rect 2392 190 2393 198
rect 2408 190 2421 198
rect 2392 182 2408 190
rect 2389 175 2408 178
rect 2389 166 2411 175
rect 2362 156 2411 166
rect 2362 150 2392 156
rect 2411 151 2416 156
rect 2334 134 2408 150
rect 2426 142 2456 198
rect 2491 188 2699 198
rect 2734 194 2779 198
rect 2782 197 2783 198
rect 2798 197 2811 198
rect 2517 158 2706 188
rect 2532 155 2706 158
rect 2525 152 2706 155
rect 2334 132 2347 134
rect 2362 132 2396 134
rect 2334 116 2408 132
rect 2435 128 2448 142
rect 2463 128 2479 144
rect 2525 139 2536 152
rect 2318 94 2319 110
rect 2334 94 2347 116
rect 2362 94 2392 116
rect 2435 112 2497 128
rect 2525 121 2536 137
rect 2541 132 2551 152
rect 2561 132 2575 152
rect 2578 139 2587 152
rect 2603 139 2612 152
rect 2541 121 2575 132
rect 2578 121 2586 137
rect 2603 121 2612 137
rect 2619 132 2629 152
rect 2639 132 2653 152
rect 2654 139 2665 152
rect 2619 121 2653 132
rect 2654 121 2665 137
rect 2711 128 2727 144
rect 2734 142 2764 194
rect 2798 190 2799 197
rect 2783 182 2799 190
rect 2770 150 2783 169
rect 2798 150 2828 166
rect 2770 134 2844 150
rect 2770 132 2783 134
rect 2798 132 2832 134
rect 2435 110 2448 112
rect 2463 110 2497 112
rect 2435 94 2497 110
rect 2541 105 2554 108
rect 2619 105 2649 116
rect 2697 112 2743 128
rect 2770 116 2844 132
rect 2697 110 2731 112
rect 2696 94 2743 110
rect 2770 94 2783 116
rect 2798 94 2828 116
rect 2855 94 2856 110
rect 2871 94 2884 254
rect 2914 150 2927 254
rect 2972 232 2973 242
rect 2988 232 3001 242
rect 2972 228 3001 232
rect 3006 228 3036 254
rect 3054 240 3070 242
rect 3142 240 3195 254
rect 3143 238 3205 240
rect 3250 238 3265 254
rect 3314 251 3344 254
rect 3314 248 3350 251
rect 3280 240 3296 242
rect 3054 228 3069 232
rect 2972 226 3069 228
rect 3097 226 3265 238
rect 3281 228 3296 232
rect 3314 229 3353 248
rect 3372 242 3379 243
rect 3378 235 3379 242
rect 3362 232 3363 235
rect 3378 232 3391 235
rect 3314 228 3344 229
rect 3353 228 3359 229
rect 3362 228 3391 232
rect 3281 227 3391 228
rect 3281 226 3397 227
rect 2956 218 3007 226
rect 2956 206 2981 218
rect 2988 206 3007 218
rect 3038 218 3088 226
rect 3038 210 3054 218
rect 3061 216 3088 218
rect 3097 216 3318 226
rect 3061 206 3318 216
rect 3347 218 3397 226
rect 3347 209 3363 218
rect 2956 198 3007 206
rect 3054 198 3318 206
rect 3344 206 3363 209
rect 3370 206 3397 218
rect 3344 198 3397 206
rect 2972 190 2973 198
rect 2988 190 3001 198
rect 2972 182 2988 190
rect 2969 175 2988 178
rect 2969 166 2991 175
rect 2942 156 2991 166
rect 2942 150 2972 156
rect 2991 151 2996 156
rect 2914 134 2988 150
rect 3006 142 3036 198
rect 3071 188 3279 198
rect 3314 194 3359 198
rect 3362 197 3363 198
rect 3378 197 3391 198
rect 3097 158 3286 188
rect 3112 155 3286 158
rect 3105 152 3286 155
rect 2914 132 2927 134
rect 2942 132 2976 134
rect 2914 116 2988 132
rect 3015 128 3028 142
rect 3043 128 3059 144
rect 3105 139 3116 152
rect 2898 94 2899 110
rect 2914 94 2927 116
rect 2942 94 2972 116
rect 3015 112 3077 128
rect 3105 121 3116 137
rect 3121 132 3131 152
rect 3141 132 3155 152
rect 3158 139 3167 152
rect 3183 139 3192 152
rect 3121 121 3155 132
rect 3158 121 3166 137
rect 3183 121 3192 137
rect 3199 132 3209 152
rect 3219 132 3233 152
rect 3234 139 3245 152
rect 3199 121 3233 132
rect 3234 121 3245 137
rect 3291 128 3307 144
rect 3314 142 3344 194
rect 3378 190 3379 197
rect 3363 182 3379 190
rect 3350 150 3363 169
rect 3378 150 3408 166
rect 3350 134 3424 150
rect 3350 132 3363 134
rect 3378 132 3412 134
rect 3015 110 3028 112
rect 3043 110 3077 112
rect 3015 94 3077 110
rect 3121 105 3134 108
rect 3199 105 3229 116
rect 3277 112 3323 128
rect 3350 116 3424 132
rect 3277 110 3311 112
rect 3276 94 3323 110
rect 3350 94 3363 116
rect 3378 94 3408 116
rect 3435 94 3436 110
rect 3451 94 3464 254
rect 3494 150 3507 254
rect 3552 232 3553 242
rect 3568 232 3581 242
rect 3552 228 3581 232
rect 3586 228 3616 254
rect 3634 240 3650 242
rect 3722 240 3775 254
rect 3723 238 3787 240
rect 3830 238 3845 254
rect 3894 251 3924 254
rect 3894 248 3930 251
rect 3860 240 3876 242
rect 3634 228 3649 232
rect 3552 226 3649 228
rect 3677 226 3845 238
rect 3861 228 3876 232
rect 3894 229 3933 248
rect 3952 242 3959 243
rect 3958 235 3959 242
rect 3942 232 3943 235
rect 3958 232 3971 235
rect 3894 228 3924 229
rect 3933 228 3939 229
rect 3942 228 3971 232
rect 3861 227 3971 228
rect 3861 226 3977 227
rect 3536 218 3587 226
rect 3536 206 3561 218
rect 3568 206 3587 218
rect 3618 218 3668 226
rect 3618 210 3634 218
rect 3641 216 3668 218
rect 3677 216 3898 226
rect 3641 206 3898 216
rect 3927 218 3977 226
rect 3927 209 3943 218
rect 3536 198 3587 206
rect 3634 198 3898 206
rect 3924 206 3943 209
rect 3950 206 3977 218
rect 3924 198 3977 206
rect 3552 190 3553 198
rect 3568 190 3581 198
rect 3552 182 3568 190
rect 3549 175 3568 178
rect 3549 166 3571 175
rect 3522 156 3571 166
rect 3522 150 3552 156
rect 3571 151 3576 156
rect 3494 134 3568 150
rect 3586 142 3616 198
rect 3651 188 3859 198
rect 3894 194 3939 198
rect 3942 197 3943 198
rect 3958 197 3971 198
rect 3677 158 3866 188
rect 3692 155 3866 158
rect 3685 152 3866 155
rect 3494 132 3507 134
rect 3522 132 3556 134
rect 3494 116 3568 132
rect 3595 128 3608 142
rect 3623 128 3639 144
rect 3685 139 3696 152
rect 3478 94 3479 110
rect 3494 94 3507 116
rect 3522 94 3552 116
rect 3595 112 3657 128
rect 3685 121 3696 137
rect 3701 132 3711 152
rect 3721 132 3735 152
rect 3738 139 3747 152
rect 3763 139 3772 152
rect 3701 121 3735 132
rect 3738 121 3746 137
rect 3763 121 3772 137
rect 3779 132 3789 152
rect 3799 132 3813 152
rect 3814 139 3825 152
rect 3779 121 3813 132
rect 3814 121 3825 137
rect 3871 128 3887 144
rect 3894 142 3924 194
rect 3958 190 3959 197
rect 3943 182 3959 190
rect 3930 150 3943 169
rect 3958 150 3988 166
rect 3930 134 4004 150
rect 3930 132 3943 134
rect 3958 132 3992 134
rect 3595 110 3608 112
rect 3623 110 3657 112
rect 3595 94 3657 110
rect 3701 105 3714 108
rect 3779 105 3809 116
rect 3857 112 3903 128
rect 3930 116 4004 132
rect 3857 110 3891 112
rect 3856 94 3903 110
rect 3930 94 3943 116
rect 3958 94 3988 116
rect 4015 94 4016 110
rect 4031 94 4044 254
rect 4074 150 4087 254
rect 4132 232 4133 242
rect 4148 232 4161 242
rect 4132 228 4161 232
rect 4166 228 4196 254
rect 4214 240 4230 242
rect 4302 240 4355 254
rect 4303 238 4367 240
rect 4410 238 4425 254
rect 4474 251 4504 254
rect 4611 253 6944 254
rect 4474 248 4510 251
rect 4440 240 4456 242
rect 4214 228 4229 232
rect 4132 226 4229 228
rect 4257 226 4425 238
rect 4441 228 4456 232
rect 4474 229 4513 248
rect 4532 242 4539 243
rect 4538 235 4539 242
rect 4522 232 4523 235
rect 4538 232 4551 235
rect 4474 228 4504 229
rect 4513 228 4519 229
rect 4522 228 4551 232
rect 4441 227 4551 228
rect 4441 226 4557 227
rect 4116 218 4167 226
rect 4116 206 4141 218
rect 4148 206 4167 218
rect 4198 218 4248 226
rect 4198 210 4214 218
rect 4221 216 4248 218
rect 4257 216 4478 226
rect 4221 206 4478 216
rect 4507 218 4557 226
rect 4507 209 4523 218
rect 4116 198 4167 206
rect 4214 198 4478 206
rect 4504 206 4523 209
rect 4530 206 4557 218
rect 4504 198 4557 206
rect 4132 190 4133 198
rect 4148 190 4161 198
rect 4132 182 4148 190
rect 4129 175 4148 178
rect 4129 166 4151 175
rect 4102 156 4151 166
rect 4102 150 4132 156
rect 4151 151 4156 156
rect 4074 134 4148 150
rect 4166 142 4196 198
rect 4231 188 4439 198
rect 4474 194 4519 198
rect 4522 197 4523 198
rect 4538 197 4551 198
rect 4257 158 4446 188
rect 4272 155 4446 158
rect 4265 152 4446 155
rect 4074 132 4087 134
rect 4102 132 4136 134
rect 4074 116 4148 132
rect 4175 128 4188 142
rect 4203 128 4219 144
rect 4265 139 4276 152
rect 4058 94 4059 110
rect 4074 94 4087 116
rect 4102 94 4132 116
rect 4175 112 4237 128
rect 4265 121 4276 137
rect 4281 132 4291 152
rect 4301 132 4315 152
rect 4318 139 4327 152
rect 4343 139 4352 152
rect 4281 121 4315 132
rect 4318 121 4326 137
rect 4343 121 4352 137
rect 4359 132 4369 152
rect 4379 132 4393 152
rect 4394 139 4405 152
rect 4359 121 4393 132
rect 4394 121 4405 137
rect 4451 128 4467 144
rect 4474 142 4504 194
rect 4538 190 4539 197
rect 4523 182 4539 190
rect 4510 150 4523 169
rect 4538 150 4568 166
rect 4510 134 4584 150
rect 4510 132 4523 134
rect 4538 132 4572 134
rect 4175 110 4188 112
rect 4203 110 4237 112
rect 4175 94 4237 110
rect 4281 105 4294 108
rect 4359 105 4389 116
rect 4437 112 4483 128
rect 4510 116 4584 132
rect 4437 110 4471 112
rect 4436 94 4483 110
rect 4510 94 4523 116
rect 4538 94 4568 116
rect 4595 94 4596 110
rect 4611 94 4624 253
rect 4654 149 4667 253
rect 4712 231 4713 241
rect 4733 239 4741 241
rect 4731 237 4741 239
rect 4728 231 4741 237
rect 4712 227 4741 231
rect 4746 227 4776 253
rect 4794 239 4810 241
rect 4882 239 4933 253
rect 4883 237 4947 239
rect 4990 237 5005 253
rect 5054 250 5084 253
rect 5054 247 5090 250
rect 5020 239 5036 241
rect 4794 227 4809 231
rect 4712 225 4809 227
rect 4837 225 5005 237
rect 5021 227 5036 231
rect 5054 228 5093 247
rect 5112 241 5119 242
rect 5118 234 5119 241
rect 5102 231 5103 234
rect 5118 231 5131 234
rect 5054 227 5084 228
rect 5093 227 5099 228
rect 5102 227 5131 231
rect 5021 226 5131 227
rect 5021 225 5137 226
rect 4696 217 4747 225
rect 4696 205 4721 217
rect 4728 205 4747 217
rect 4778 217 4828 225
rect 4778 209 4794 217
rect 4801 215 4828 217
rect 4837 215 5058 225
rect 4801 205 5058 215
rect 5087 217 5137 225
rect 5087 208 5103 217
rect 4696 197 4747 205
rect 4794 197 5058 205
rect 5084 205 5103 208
rect 5110 205 5137 217
rect 5084 197 5137 205
rect 4712 189 4713 197
rect 4728 189 4741 197
rect 4712 181 4728 189
rect 4709 174 4728 177
rect 4709 165 4731 174
rect 4682 155 4731 165
rect 4682 149 4712 155
rect 4731 150 4736 155
rect 4654 133 4728 149
rect 4746 141 4776 197
rect 4811 187 5019 197
rect 5054 193 5099 197
rect 5102 196 5103 197
rect 5118 196 5131 197
rect 4837 157 5026 187
rect 4852 154 5026 157
rect 4845 151 5026 154
rect 4654 131 4667 133
rect 4682 131 4716 133
rect 4654 115 4728 131
rect 4755 127 4768 141
rect 4783 127 4799 143
rect 4845 138 4856 151
rect -8 86 33 94
rect -8 60 7 86
rect 14 60 33 86
rect 97 82 159 94
rect 171 82 246 94
rect 304 82 379 94
rect 391 82 422 94
rect 428 82 463 94
rect 97 80 259 82
rect -8 52 33 60
rect 115 56 128 80
rect 143 78 158 80
rect -2 42 -1 52
rect 14 42 27 52
rect 42 42 72 56
rect 115 42 158 56
rect 182 53 189 60
rect 192 56 259 80
rect 291 80 463 82
rect 261 58 289 62
rect 291 58 371 80
rect 392 78 407 80
rect 261 56 371 58
rect 192 52 371 56
rect 165 42 195 52
rect 197 42 350 52
rect 358 42 388 52
rect 392 42 422 56
rect 450 42 463 80
rect 535 86 570 94
rect 535 60 536 86
rect 543 60 570 86
rect 478 42 508 56
rect 535 52 570 60
rect 572 86 613 94
rect 572 60 587 86
rect 594 60 613 86
rect 677 82 739 94
rect 751 82 826 94
rect 884 82 959 94
rect 971 82 1002 94
rect 1008 82 1043 94
rect 677 80 839 82
rect 572 52 613 60
rect 695 56 708 80
rect 723 78 738 80
rect 535 42 536 52
rect 551 42 564 52
rect 578 42 579 52
rect 594 42 607 52
rect 622 42 652 56
rect 695 42 738 56
rect 762 53 769 60
rect 772 56 839 80
rect 871 80 1043 82
rect 841 58 869 62
rect 871 58 951 80
rect 972 78 987 80
rect 841 56 951 58
rect 772 52 951 56
rect 745 42 775 52
rect 777 42 930 52
rect 938 42 968 52
rect 972 42 1002 56
rect 1030 42 1043 80
rect 1115 86 1150 94
rect 1115 60 1116 86
rect 1123 60 1150 86
rect 1058 42 1088 56
rect 1115 52 1150 60
rect 1152 86 1193 94
rect 1152 60 1167 86
rect 1174 60 1193 86
rect 1257 82 1319 94
rect 1331 82 1406 94
rect 1464 82 1539 94
rect 1551 82 1582 94
rect 1588 82 1623 94
rect 1257 80 1419 82
rect 1152 52 1193 60
rect 1275 56 1288 80
rect 1303 78 1318 80
rect 1115 42 1116 52
rect 1131 42 1144 52
rect 1158 42 1159 52
rect 1174 42 1187 52
rect 1202 42 1232 56
rect 1275 42 1318 56
rect 1342 53 1349 60
rect 1352 56 1419 80
rect 1451 80 1623 82
rect 1421 58 1449 62
rect 1451 58 1531 80
rect 1552 78 1567 80
rect 1421 56 1531 58
rect 1352 52 1531 56
rect 1325 42 1355 52
rect 1357 42 1510 52
rect 1518 42 1548 52
rect 1552 42 1582 56
rect 1610 42 1623 80
rect 1695 86 1730 94
rect 1695 60 1696 86
rect 1703 60 1730 86
rect 1638 42 1668 56
rect 1695 52 1730 60
rect 1732 86 1773 94
rect 1732 60 1747 86
rect 1754 60 1773 86
rect 1837 82 1899 94
rect 1911 82 1986 94
rect 2044 82 2119 94
rect 2131 82 2162 94
rect 2168 82 2203 94
rect 1837 80 1999 82
rect 1732 52 1773 60
rect 1855 56 1868 80
rect 1883 78 1898 80
rect 1695 42 1696 52
rect 1711 42 1724 52
rect 1738 42 1739 52
rect 1754 42 1767 52
rect 1782 42 1812 56
rect 1855 42 1898 56
rect 1922 53 1929 60
rect 1932 56 1999 80
rect 2031 80 2203 82
rect 2001 58 2029 62
rect 2031 58 2111 80
rect 2132 78 2147 80
rect 2001 56 2111 58
rect 1932 52 2111 56
rect 1905 42 1935 52
rect 1937 42 2090 52
rect 2098 42 2128 52
rect 2132 42 2162 56
rect 2190 42 2203 80
rect 2275 86 2310 94
rect 2275 60 2276 86
rect 2283 60 2310 86
rect 2218 42 2248 56
rect 2275 52 2310 60
rect 2312 86 2353 94
rect 2312 60 2327 86
rect 2334 60 2353 86
rect 2417 82 2479 94
rect 2491 82 2566 94
rect 2624 82 2699 94
rect 2711 82 2742 94
rect 2748 82 2783 94
rect 2417 80 2579 82
rect 2312 52 2353 60
rect 2435 56 2448 80
rect 2463 78 2478 80
rect 2275 42 2276 52
rect 2291 42 2304 52
rect 2318 42 2319 52
rect 2334 42 2347 52
rect 2362 42 2392 56
rect 2435 42 2478 56
rect 2502 53 2509 60
rect 2512 56 2579 80
rect 2611 80 2783 82
rect 2581 58 2609 62
rect 2611 58 2691 80
rect 2712 78 2727 80
rect 2581 56 2691 58
rect 2512 52 2691 56
rect 2485 42 2515 52
rect 2517 42 2670 52
rect 2678 42 2708 52
rect 2712 42 2742 56
rect 2770 42 2783 80
rect 2855 86 2890 94
rect 2855 60 2856 86
rect 2863 60 2890 86
rect 2798 42 2828 56
rect 2855 52 2890 60
rect 2892 86 2933 94
rect 2892 60 2907 86
rect 2914 60 2933 86
rect 2997 82 3059 94
rect 3071 82 3146 94
rect 3204 82 3279 94
rect 3291 82 3322 94
rect 3328 82 3363 94
rect 2997 80 3159 82
rect 2892 52 2933 60
rect 3015 56 3028 80
rect 3043 78 3058 80
rect 2855 42 2856 52
rect 2871 42 2884 52
rect 2898 42 2899 52
rect 2914 42 2927 52
rect 2942 42 2972 56
rect 3015 42 3058 56
rect 3082 53 3089 60
rect 3092 56 3159 80
rect 3191 80 3363 82
rect 3161 58 3189 62
rect 3191 58 3271 80
rect 3292 78 3307 80
rect 3161 56 3271 58
rect 3092 52 3271 56
rect 3065 42 3095 52
rect 3097 42 3250 52
rect 3258 42 3288 52
rect 3292 42 3322 56
rect 3350 42 3363 80
rect 3435 86 3470 94
rect 3435 60 3436 86
rect 3443 60 3470 86
rect 3378 42 3408 56
rect 3435 52 3470 60
rect 3472 86 3513 94
rect 3472 60 3487 86
rect 3494 60 3513 86
rect 3577 82 3639 94
rect 3651 82 3726 94
rect 3784 82 3859 94
rect 3871 82 3902 94
rect 3908 82 3943 94
rect 3577 80 3739 82
rect 3472 52 3513 60
rect 3595 56 3608 80
rect 3623 78 3638 80
rect 3435 42 3436 52
rect 3451 42 3464 52
rect 3478 42 3479 52
rect 3494 42 3507 52
rect 3522 42 3552 56
rect 3595 42 3638 56
rect 3662 53 3669 60
rect 3672 56 3739 80
rect 3771 80 3943 82
rect 3741 58 3769 62
rect 3771 58 3851 80
rect 3872 78 3887 80
rect 3741 56 3851 58
rect 3672 52 3851 56
rect 3645 42 3675 52
rect 3677 42 3830 52
rect 3838 42 3868 52
rect 3872 42 3902 56
rect 3930 42 3943 80
rect 4015 86 4050 94
rect 4015 60 4016 86
rect 4023 60 4050 86
rect 3958 42 3988 56
rect 4015 52 4050 60
rect 4052 86 4093 94
rect 4052 60 4067 86
rect 4074 60 4093 86
rect 4157 82 4219 94
rect 4231 82 4306 94
rect 4364 82 4439 94
rect 4451 82 4482 94
rect 4488 82 4523 94
rect 4157 80 4319 82
rect 4052 52 4093 60
rect 4175 56 4188 80
rect 4203 78 4218 80
rect 4015 42 4016 52
rect 4031 42 4044 52
rect 4058 42 4059 52
rect 4074 42 4087 52
rect 4102 42 4132 56
rect 4175 42 4218 56
rect 4242 53 4249 60
rect 4252 56 4319 80
rect 4351 80 4523 82
rect 4321 58 4349 62
rect 4351 58 4431 80
rect 4452 78 4467 80
rect 4321 56 4431 58
rect 4252 52 4431 56
rect 4225 42 4255 52
rect 4257 42 4410 52
rect 4418 42 4448 52
rect 4452 42 4482 56
rect 4510 42 4523 80
rect 4595 86 4630 94
rect 4638 93 4639 109
rect 4654 93 4667 115
rect 4682 93 4712 115
rect 4755 111 4817 127
rect 4845 120 4856 136
rect 4861 131 4871 151
rect 4881 131 4895 151
rect 4898 138 4907 151
rect 4923 138 4932 151
rect 4861 120 4895 131
rect 4898 120 4907 136
rect 4923 120 4932 136
rect 4939 131 4949 151
rect 4959 131 4973 151
rect 4974 138 4985 151
rect 4939 120 4973 131
rect 4974 120 4985 136
rect 5031 127 5047 143
rect 5054 141 5084 193
rect 5118 189 5119 196
rect 5103 181 5119 189
rect 5090 149 5103 168
rect 5118 149 5148 165
rect 5090 133 5164 149
rect 5090 131 5103 133
rect 5118 131 5152 133
rect 4755 109 4768 111
rect 4783 109 4817 111
rect 4755 93 4817 109
rect 4861 104 4877 107
rect 4939 104 4969 115
rect 5017 111 5063 127
rect 5090 115 5164 131
rect 5017 109 5051 111
rect 5016 93 5063 109
rect 5090 93 5103 115
rect 5118 93 5148 115
rect 5175 93 5176 109
rect 5191 93 5204 253
rect 5234 149 5247 253
rect 5292 231 5293 241
rect 5313 239 5321 241
rect 5311 237 5321 239
rect 5308 231 5321 237
rect 5292 227 5321 231
rect 5326 227 5356 253
rect 5374 239 5390 241
rect 5462 239 5513 253
rect 5463 237 5527 239
rect 5570 237 5585 253
rect 5634 250 5664 253
rect 5634 247 5670 250
rect 5600 239 5616 241
rect 5374 227 5389 231
rect 5292 225 5389 227
rect 5417 225 5585 237
rect 5601 227 5616 231
rect 5634 228 5673 247
rect 5692 241 5699 242
rect 5698 234 5699 241
rect 5682 231 5683 234
rect 5698 231 5711 234
rect 5634 227 5664 228
rect 5673 227 5679 228
rect 5682 227 5711 231
rect 5601 226 5711 227
rect 5601 225 5717 226
rect 5276 217 5327 225
rect 5276 205 5301 217
rect 5308 205 5327 217
rect 5358 217 5408 225
rect 5358 209 5374 217
rect 5381 215 5408 217
rect 5417 215 5638 225
rect 5381 205 5638 215
rect 5667 217 5717 225
rect 5667 208 5683 217
rect 5276 197 5327 205
rect 5374 197 5638 205
rect 5664 205 5683 208
rect 5690 205 5717 217
rect 5664 197 5717 205
rect 5292 189 5293 197
rect 5308 189 5321 197
rect 5292 181 5308 189
rect 5289 174 5308 177
rect 5289 165 5311 174
rect 5262 155 5311 165
rect 5262 149 5292 155
rect 5311 150 5316 155
rect 5234 133 5308 149
rect 5326 141 5356 197
rect 5391 187 5599 197
rect 5634 193 5679 197
rect 5682 196 5683 197
rect 5698 196 5711 197
rect 5417 157 5606 187
rect 5432 154 5606 157
rect 5425 151 5606 154
rect 5234 131 5247 133
rect 5262 131 5296 133
rect 5234 115 5308 131
rect 5335 127 5348 141
rect 5363 127 5379 143
rect 5425 138 5436 151
rect 5218 93 5219 109
rect 5234 93 5247 115
rect 5262 93 5292 115
rect 5335 111 5397 127
rect 5425 120 5436 136
rect 5441 131 5451 151
rect 5461 131 5475 151
rect 5478 138 5487 151
rect 5503 138 5512 151
rect 5441 120 5475 131
rect 5478 120 5487 136
rect 5503 120 5512 136
rect 5519 131 5529 151
rect 5539 131 5553 151
rect 5554 138 5565 151
rect 5519 120 5553 131
rect 5554 120 5565 136
rect 5611 127 5627 143
rect 5634 141 5664 193
rect 5698 189 5699 196
rect 5683 181 5699 189
rect 5670 149 5683 168
rect 5698 149 5728 165
rect 5670 133 5744 149
rect 5670 131 5683 133
rect 5698 131 5732 133
rect 5335 109 5348 111
rect 5363 109 5397 111
rect 5335 93 5397 109
rect 5441 104 5457 107
rect 5519 104 5549 115
rect 5597 111 5643 127
rect 5670 115 5744 131
rect 5597 109 5631 111
rect 5596 93 5643 109
rect 5670 93 5683 115
rect 5698 93 5728 115
rect 5755 93 5756 109
rect 5771 93 5784 253
rect 5814 149 5827 253
rect 5872 231 5873 241
rect 5893 239 5901 241
rect 5891 237 5901 239
rect 5888 231 5901 237
rect 5872 227 5901 231
rect 5906 227 5936 253
rect 5954 239 5970 241
rect 6042 239 6093 253
rect 6043 237 6107 239
rect 6150 237 6165 253
rect 6214 250 6244 253
rect 6214 247 6250 250
rect 6180 239 6196 241
rect 5954 227 5969 231
rect 5872 225 5969 227
rect 5997 225 6165 237
rect 6181 227 6196 231
rect 6214 228 6253 247
rect 6272 241 6279 242
rect 6278 234 6279 241
rect 6262 231 6263 234
rect 6278 231 6291 234
rect 6214 227 6244 228
rect 6253 227 6259 228
rect 6262 227 6291 231
rect 6181 226 6291 227
rect 6181 225 6297 226
rect 5856 217 5907 225
rect 5856 205 5881 217
rect 5888 205 5907 217
rect 5938 217 5988 225
rect 5938 209 5954 217
rect 5961 215 5988 217
rect 5997 215 6218 225
rect 5961 205 6218 215
rect 6247 217 6297 225
rect 6247 208 6263 217
rect 5856 197 5907 205
rect 5954 197 6218 205
rect 6244 205 6263 208
rect 6270 205 6297 217
rect 6244 197 6297 205
rect 5872 189 5873 197
rect 5888 189 5901 197
rect 5872 181 5888 189
rect 5869 174 5888 177
rect 5869 165 5891 174
rect 5842 155 5891 165
rect 5842 149 5872 155
rect 5891 150 5896 155
rect 5814 133 5888 149
rect 5906 141 5936 197
rect 5971 187 6179 197
rect 6214 193 6259 197
rect 6262 196 6263 197
rect 6278 196 6291 197
rect 5997 157 6186 187
rect 6012 154 6186 157
rect 6005 151 6186 154
rect 5814 131 5827 133
rect 5842 131 5876 133
rect 5814 115 5888 131
rect 5915 127 5928 141
rect 5943 127 5959 143
rect 6005 138 6016 151
rect 5798 93 5799 109
rect 5814 93 5827 115
rect 5842 93 5872 115
rect 5915 111 5977 127
rect 6005 120 6016 136
rect 6021 131 6031 151
rect 6041 131 6055 151
rect 6058 138 6067 151
rect 6083 138 6092 151
rect 6021 120 6055 131
rect 6058 120 6067 136
rect 6083 120 6092 136
rect 6099 131 6109 151
rect 6119 131 6133 151
rect 6134 138 6145 151
rect 6099 120 6133 131
rect 6134 120 6145 136
rect 6191 127 6207 143
rect 6214 141 6244 193
rect 6278 189 6279 196
rect 6263 181 6279 189
rect 6250 149 6263 168
rect 6278 149 6308 165
rect 6250 133 6324 149
rect 6250 131 6263 133
rect 6278 131 6312 133
rect 5915 109 5928 111
rect 5943 109 5977 111
rect 5915 93 5977 109
rect 6021 104 6037 107
rect 6099 104 6129 115
rect 6177 111 6223 127
rect 6250 115 6324 131
rect 6177 109 6211 111
rect 6176 93 6223 109
rect 6250 93 6263 115
rect 6278 93 6308 115
rect 6335 93 6336 109
rect 6351 93 6364 253
rect 6394 149 6407 253
rect 6452 231 6453 241
rect 6473 239 6481 241
rect 6471 237 6481 239
rect 6468 231 6481 237
rect 6452 227 6481 231
rect 6486 227 6516 253
rect 6534 239 6550 241
rect 6622 239 6673 253
rect 6623 237 6687 239
rect 6730 237 6745 253
rect 6794 250 6824 253
rect 6794 247 6830 250
rect 6760 239 6776 241
rect 6534 227 6549 231
rect 6452 225 6549 227
rect 6577 225 6745 237
rect 6761 227 6776 231
rect 6794 228 6833 247
rect 6852 241 6859 242
rect 6858 234 6859 241
rect 6842 231 6843 234
rect 6858 231 6871 234
rect 6794 227 6824 228
rect 6833 227 6839 228
rect 6842 227 6871 231
rect 6761 226 6871 227
rect 6761 225 6877 226
rect 6436 217 6487 225
rect 6436 205 6461 217
rect 6468 205 6487 217
rect 6518 217 6568 225
rect 6518 209 6534 217
rect 6541 215 6568 217
rect 6577 215 6798 225
rect 6541 205 6798 215
rect 6827 217 6877 225
rect 6827 208 6843 217
rect 6436 197 6487 205
rect 6534 197 6798 205
rect 6824 205 6843 208
rect 6850 205 6877 217
rect 6824 197 6877 205
rect 6452 189 6453 197
rect 6468 189 6481 197
rect 6452 181 6468 189
rect 6449 174 6468 177
rect 6449 165 6471 174
rect 6422 155 6471 165
rect 6422 149 6452 155
rect 6471 150 6476 155
rect 6394 133 6468 149
rect 6486 141 6516 197
rect 6551 187 6759 197
rect 6794 193 6839 197
rect 6842 196 6843 197
rect 6858 196 6871 197
rect 6577 157 6766 187
rect 6592 154 6766 157
rect 6585 151 6766 154
rect 6394 131 6407 133
rect 6422 131 6456 133
rect 6394 115 6468 131
rect 6495 127 6508 141
rect 6523 127 6539 143
rect 6585 138 6596 151
rect 6378 93 6379 109
rect 6394 93 6407 115
rect 6422 93 6452 115
rect 6495 111 6557 127
rect 6585 120 6596 136
rect 6601 131 6611 151
rect 6621 131 6635 151
rect 6638 138 6647 151
rect 6663 138 6672 151
rect 6601 120 6635 131
rect 6638 120 6647 136
rect 6663 120 6672 136
rect 6679 131 6689 151
rect 6699 131 6713 151
rect 6714 138 6725 151
rect 6679 120 6713 131
rect 6714 120 6725 136
rect 6771 127 6787 143
rect 6794 141 6824 193
rect 6858 189 6859 196
rect 6843 181 6859 189
rect 6830 149 6843 168
rect 6858 149 6888 165
rect 6830 133 6904 149
rect 6830 131 6843 133
rect 6858 131 6892 133
rect 6495 109 6508 111
rect 6523 109 6557 111
rect 6495 93 6557 109
rect 6601 104 6617 107
rect 6679 104 6709 115
rect 6757 111 6803 127
rect 6830 115 6904 131
rect 6757 109 6791 111
rect 6756 93 6803 109
rect 6830 93 6843 115
rect 6858 93 6888 115
rect 6915 93 6916 109
rect 6931 93 6944 253
rect 4595 60 4596 86
rect 4603 60 4630 86
rect 4538 42 4568 56
rect 4595 52 4630 60
rect 4632 85 4673 93
rect 4632 59 4647 85
rect 4654 59 4673 85
rect 4737 81 4799 93
rect 4811 81 4886 93
rect 4944 81 5019 93
rect 5031 81 5062 93
rect 5068 81 5103 93
rect 4737 79 4899 81
rect 4755 61 4768 79
rect 4783 77 4798 79
rect 4595 42 4596 52
rect 4611 42 4624 52
rect 4632 51 4673 59
rect 4756 55 4768 61
rect 4832 61 4899 79
rect 4931 79 5103 81
rect 4931 61 5011 79
rect 5032 77 5047 79
rect -2 41 4624 42
rect 4638 41 4639 51
rect 4654 41 4667 51
rect 4682 41 4712 55
rect 4756 41 4798 55
rect 4822 52 4829 59
rect 4832 51 5011 61
rect 4805 41 4835 51
rect 4837 41 4990 51
rect 4998 41 5028 51
rect 5032 41 5062 55
rect 5090 41 5103 79
rect 5175 85 5210 93
rect 5175 59 5176 85
rect 5183 59 5210 85
rect 5118 41 5148 55
rect 5175 51 5210 59
rect 5212 85 5253 93
rect 5212 59 5227 85
rect 5234 59 5253 85
rect 5317 81 5379 93
rect 5391 81 5466 93
rect 5524 81 5599 93
rect 5611 81 5642 93
rect 5648 81 5683 93
rect 5317 79 5479 81
rect 5335 61 5348 79
rect 5363 77 5378 79
rect 5212 51 5253 59
rect 5336 55 5348 61
rect 5412 61 5479 79
rect 5511 79 5683 81
rect 5511 61 5591 79
rect 5612 77 5627 79
rect 5175 41 5176 51
rect 5191 41 5204 51
rect 5218 41 5219 51
rect 5234 41 5247 51
rect 5262 41 5292 55
rect 5336 41 5378 55
rect 5402 52 5409 59
rect 5412 51 5591 61
rect 5385 41 5415 51
rect 5417 41 5570 51
rect 5578 41 5608 51
rect 5612 41 5642 55
rect 5670 41 5683 79
rect 5755 85 5790 93
rect 5755 59 5756 85
rect 5763 59 5790 85
rect 5698 41 5728 55
rect 5755 51 5790 59
rect 5792 85 5833 93
rect 5792 59 5807 85
rect 5814 59 5833 85
rect 5897 81 5959 93
rect 5971 81 6046 93
rect 6104 81 6179 93
rect 6191 81 6222 93
rect 6228 81 6263 93
rect 5897 79 6059 81
rect 5915 61 5928 79
rect 5943 77 5958 79
rect 5792 51 5833 59
rect 5916 55 5928 61
rect 5992 61 6059 79
rect 6091 79 6263 81
rect 6091 61 6171 79
rect 6192 77 6207 79
rect 5755 41 5756 51
rect 5771 41 5784 51
rect 5798 41 5799 51
rect 5814 41 5827 51
rect 5842 41 5872 55
rect 5916 41 5958 55
rect 5982 52 5989 59
rect 5992 51 6171 61
rect 5965 41 5995 51
rect 5997 41 6150 51
rect 6158 41 6188 51
rect 6192 41 6222 55
rect 6250 41 6263 79
rect 6335 85 6370 93
rect 6335 59 6336 85
rect 6343 59 6370 85
rect 6278 41 6308 55
rect 6335 51 6370 59
rect 6372 85 6413 93
rect 6372 59 6387 85
rect 6394 59 6413 85
rect 6477 81 6539 93
rect 6551 81 6626 93
rect 6684 81 6759 93
rect 6771 81 6802 93
rect 6808 81 6843 93
rect 6477 79 6639 81
rect 6495 61 6508 79
rect 6523 77 6538 79
rect 6372 51 6413 59
rect 6496 55 6508 61
rect 6572 61 6639 79
rect 6671 79 6843 81
rect 6671 61 6751 79
rect 6772 77 6787 79
rect 6335 41 6336 51
rect 6351 41 6364 51
rect 6378 41 6379 51
rect 6394 41 6407 51
rect 6422 41 6452 55
rect 6496 41 6538 55
rect 6562 52 6569 59
rect 6572 51 6751 61
rect 6545 41 6575 51
rect 6577 41 6730 51
rect 6738 41 6768 51
rect 6772 41 6802 55
rect 6830 41 6843 79
rect 6915 85 6950 93
rect 6915 59 6916 85
rect 6923 59 6950 85
rect 6858 41 6888 55
rect 6915 51 6950 59
rect 6915 41 6916 51
rect 6931 41 6944 51
rect -2 36 6944 41
rect -1 28 6944 36
rect 14 -2 27 28
rect 42 10 72 28
rect 115 14 129 28
rect 165 14 385 28
rect 116 12 129 14
rect 82 0 97 12
rect 79 -2 101 0
rect 106 -2 136 12
rect 197 10 350 14
rect 179 -2 371 10
rect 414 -2 444 12
rect 450 -2 463 28
rect 478 10 508 28
rect 551 -2 564 28
rect 594 -2 607 28
rect 622 10 652 28
rect 695 14 709 28
rect 745 14 965 28
rect 696 12 709 14
rect 662 0 677 12
rect 659 -2 681 0
rect 686 -2 716 12
rect 777 10 930 14
rect 759 -2 951 10
rect 994 -2 1024 12
rect 1030 -2 1043 28
rect 1058 10 1088 28
rect 1131 -2 1144 28
rect 1174 -2 1187 28
rect 1202 10 1232 28
rect 1275 14 1289 28
rect 1325 14 1545 28
rect 1276 12 1289 14
rect 1242 0 1257 12
rect 1239 -2 1261 0
rect 1266 -2 1296 12
rect 1357 10 1510 14
rect 1339 -2 1531 10
rect 1574 -2 1604 12
rect 1610 -2 1623 28
rect 1638 10 1668 28
rect 1711 -2 1724 28
rect 1754 -2 1767 28
rect 1782 10 1812 28
rect 1855 14 1869 28
rect 1905 14 2125 28
rect 1856 12 1869 14
rect 1822 0 1837 12
rect 1819 -2 1841 0
rect 1846 -2 1876 12
rect 1937 10 2090 14
rect 1919 -2 2111 10
rect 2154 -2 2184 12
rect 2190 -2 2203 28
rect 2218 10 2248 28
rect 2291 -2 2304 28
rect 2334 -2 2347 28
rect 2362 10 2392 28
rect 2435 14 2449 28
rect 2485 14 2705 28
rect 2436 12 2449 14
rect 2402 0 2417 12
rect 2399 -2 2421 0
rect 2426 -2 2456 12
rect 2517 10 2670 14
rect 2499 -2 2691 10
rect 2734 -2 2764 12
rect 2770 -2 2783 28
rect 2798 10 2828 28
rect 2871 -2 2884 28
rect 2914 -2 2927 28
rect 2942 10 2972 28
rect 3015 14 3029 28
rect 3065 14 3285 28
rect 3016 12 3029 14
rect 2982 0 2997 12
rect 2979 -2 3001 0
rect 3006 -2 3036 12
rect 3097 10 3250 14
rect 3079 -2 3271 10
rect 3314 -2 3344 12
rect 3350 -2 3363 28
rect 3378 10 3408 28
rect 3451 -2 3464 28
rect 3494 -2 3507 28
rect 3522 10 3552 28
rect 3595 14 3609 28
rect 3645 14 3865 28
rect 3596 12 3609 14
rect 3562 0 3577 12
rect 3559 -2 3581 0
rect 3586 -2 3616 12
rect 3677 10 3830 14
rect 3659 -2 3851 10
rect 3894 -2 3924 12
rect 3930 -2 3943 28
rect 3958 10 3988 28
rect 4031 -2 4044 28
rect 4074 -2 4087 28
rect 4102 10 4132 28
rect 4175 14 4189 28
rect 4225 14 4445 28
rect 4176 12 4189 14
rect 4142 0 4157 12
rect 4139 -2 4161 0
rect 4166 -2 4196 12
rect 4257 10 4410 14
rect 4239 -2 4431 10
rect 4474 -2 4504 12
rect 4510 -2 4523 28
rect 4538 10 4568 28
rect 4611 27 6944 28
rect 4611 -2 4624 27
rect -1 -3 4624 -2
rect 4654 -3 4667 27
rect 4682 9 4712 27
rect 4756 11 4769 27
rect 4805 13 5025 27
rect 4722 -1 4737 11
rect 4719 -3 4741 -1
rect 4746 -3 4776 11
rect 4837 9 4990 13
rect 4819 -3 5011 9
rect 5054 -3 5084 11
rect 5090 -3 5103 27
rect 5118 9 5148 27
rect 5191 -3 5204 27
rect 5234 -3 5247 27
rect 5262 9 5292 27
rect 5336 11 5349 27
rect 5385 13 5605 27
rect 5302 -1 5317 11
rect 5299 -3 5321 -1
rect 5326 -3 5356 11
rect 5417 9 5570 13
rect 5399 -3 5591 9
rect 5634 -3 5664 11
rect 5670 -3 5683 27
rect 5698 9 5728 27
rect 5771 -3 5784 27
rect 5814 -3 5827 27
rect 5842 9 5872 27
rect 5916 11 5929 27
rect 5965 13 6185 27
rect 5882 -1 5897 11
rect 5879 -3 5901 -1
rect 5906 -3 5936 11
rect 5997 9 6150 13
rect 5979 -3 6171 9
rect 6214 -3 6244 11
rect 6250 -3 6263 27
rect 6278 9 6308 27
rect 6351 -3 6364 27
rect 6394 -3 6407 27
rect 6422 9 6452 27
rect 6496 11 6509 27
rect 6545 13 6765 27
rect 6462 -1 6477 11
rect 6459 -3 6481 -1
rect 6486 -3 6516 11
rect 6577 9 6730 13
rect 6559 -3 6751 9
rect 6794 -3 6824 11
rect 6830 -3 6843 27
rect 6858 9 6888 27
rect 6931 -3 6944 27
rect -1 -16 6944 -3
rect 14 -120 27 -16
rect 72 -38 73 -28
rect 88 -38 101 -28
rect 72 -42 101 -38
rect 106 -42 136 -16
rect 154 -30 170 -28
rect 242 -30 295 -16
rect 243 -32 307 -30
rect 350 -32 365 -16
rect 414 -19 444 -16
rect 414 -22 450 -19
rect 380 -30 396 -28
rect 154 -42 169 -38
rect 72 -44 169 -42
rect 197 -44 365 -32
rect 381 -42 396 -38
rect 414 -41 453 -22
rect 472 -28 479 -27
rect 478 -35 479 -28
rect 462 -38 463 -35
rect 478 -38 491 -35
rect 414 -42 444 -41
rect 453 -42 459 -41
rect 462 -42 491 -38
rect 381 -43 491 -42
rect 381 -44 497 -43
rect 56 -52 107 -44
rect 56 -64 81 -52
rect 88 -64 107 -52
rect 138 -52 188 -44
rect 138 -60 154 -52
rect 161 -54 188 -52
rect 197 -54 418 -44
rect 161 -64 418 -54
rect 447 -52 497 -44
rect 447 -61 463 -52
rect 56 -72 107 -64
rect 154 -72 418 -64
rect 444 -64 463 -61
rect 470 -64 497 -52
rect 444 -72 497 -64
rect 72 -80 73 -72
rect 88 -80 101 -72
rect 72 -88 88 -80
rect 69 -95 88 -92
rect 69 -104 91 -95
rect 42 -114 91 -104
rect 42 -120 72 -114
rect 91 -119 96 -114
rect 14 -136 88 -120
rect 106 -128 136 -72
rect 171 -82 379 -72
rect 414 -76 459 -72
rect 462 -73 463 -72
rect 478 -73 491 -72
rect 197 -112 386 -82
rect 212 -115 386 -112
rect 205 -118 386 -115
rect 14 -138 27 -136
rect 42 -138 76 -136
rect 14 -154 88 -138
rect 115 -142 128 -128
rect 143 -142 159 -126
rect 205 -131 216 -118
rect -2 -176 -1 -160
rect 14 -176 27 -154
rect 42 -176 72 -154
rect 115 -158 177 -142
rect 205 -149 216 -133
rect 221 -138 231 -118
rect 241 -138 255 -118
rect 258 -131 267 -118
rect 283 -131 292 -118
rect 221 -149 255 -138
rect 258 -149 267 -133
rect 283 -149 292 -133
rect 299 -138 309 -118
rect 319 -138 333 -118
rect 334 -131 345 -118
rect 299 -149 333 -138
rect 334 -149 345 -133
rect 391 -142 407 -126
rect 414 -128 444 -76
rect 478 -80 479 -73
rect 463 -88 479 -80
rect 450 -120 463 -101
rect 478 -120 508 -104
rect 450 -136 524 -120
rect 450 -138 463 -136
rect 478 -138 512 -136
rect 115 -160 128 -158
rect 143 -160 177 -158
rect 115 -176 177 -160
rect 221 -165 237 -162
rect 299 -165 329 -154
rect 377 -158 423 -142
rect 450 -154 524 -138
rect 377 -160 411 -158
rect 376 -176 423 -160
rect 450 -176 463 -154
rect 478 -176 508 -154
rect 535 -176 536 -160
rect 551 -176 564 -16
rect 594 -120 607 -16
rect 652 -38 653 -28
rect 668 -38 681 -28
rect 652 -42 681 -38
rect 686 -42 716 -16
rect 734 -30 750 -28
rect 822 -30 875 -16
rect 823 -32 887 -30
rect 930 -32 945 -16
rect 994 -19 1024 -16
rect 994 -22 1030 -19
rect 960 -30 976 -28
rect 734 -42 749 -38
rect 652 -44 749 -42
rect 777 -44 945 -32
rect 961 -42 976 -38
rect 994 -41 1033 -22
rect 1052 -28 1059 -27
rect 1058 -35 1059 -28
rect 1042 -38 1043 -35
rect 1058 -38 1071 -35
rect 994 -42 1024 -41
rect 1033 -42 1039 -41
rect 1042 -42 1071 -38
rect 961 -43 1071 -42
rect 961 -44 1077 -43
rect 636 -52 687 -44
rect 636 -64 661 -52
rect 668 -64 687 -52
rect 718 -52 768 -44
rect 718 -60 734 -52
rect 741 -54 768 -52
rect 777 -54 998 -44
rect 741 -64 998 -54
rect 1027 -52 1077 -44
rect 1027 -61 1043 -52
rect 636 -72 687 -64
rect 734 -72 998 -64
rect 1024 -64 1043 -61
rect 1050 -64 1077 -52
rect 1024 -72 1077 -64
rect 652 -80 653 -72
rect 668 -80 681 -72
rect 652 -88 668 -80
rect 649 -95 668 -92
rect 649 -104 671 -95
rect 622 -114 671 -104
rect 622 -120 652 -114
rect 671 -119 676 -114
rect 594 -136 668 -120
rect 686 -128 716 -72
rect 751 -82 959 -72
rect 994 -76 1039 -72
rect 1042 -73 1043 -72
rect 1058 -73 1071 -72
rect 777 -112 966 -82
rect 792 -115 966 -112
rect 785 -118 966 -115
rect 594 -138 607 -136
rect 622 -138 656 -136
rect 594 -154 668 -138
rect 695 -142 708 -128
rect 723 -142 739 -126
rect 785 -131 796 -118
rect 578 -176 579 -160
rect 594 -176 607 -154
rect 622 -176 652 -154
rect 695 -158 757 -142
rect 785 -149 796 -133
rect 801 -138 811 -118
rect 821 -138 835 -118
rect 838 -131 847 -118
rect 863 -131 872 -118
rect 801 -149 835 -138
rect 838 -149 847 -133
rect 863 -149 872 -133
rect 879 -138 889 -118
rect 899 -138 913 -118
rect 914 -131 925 -118
rect 879 -149 913 -138
rect 914 -149 925 -133
rect 971 -142 987 -126
rect 994 -128 1024 -76
rect 1058 -80 1059 -73
rect 1043 -88 1059 -80
rect 1030 -120 1043 -101
rect 1058 -120 1088 -104
rect 1030 -136 1104 -120
rect 1030 -138 1043 -136
rect 1058 -138 1092 -136
rect 695 -160 708 -158
rect 723 -160 757 -158
rect 695 -176 757 -160
rect 801 -165 817 -162
rect 879 -165 909 -154
rect 957 -158 1003 -142
rect 1030 -154 1104 -138
rect 957 -160 991 -158
rect 956 -176 1003 -160
rect 1030 -176 1043 -154
rect 1058 -176 1088 -154
rect 1115 -176 1116 -160
rect 1131 -176 1144 -16
rect 1174 -120 1187 -16
rect 1232 -38 1233 -28
rect 1248 -38 1261 -28
rect 1232 -42 1261 -38
rect 1266 -42 1296 -16
rect 1314 -30 1330 -28
rect 1402 -30 1455 -16
rect 1403 -32 1467 -30
rect 1510 -32 1525 -16
rect 1574 -19 1604 -16
rect 1574 -22 1610 -19
rect 1540 -30 1556 -28
rect 1314 -42 1329 -38
rect 1232 -44 1329 -42
rect 1357 -44 1525 -32
rect 1541 -42 1556 -38
rect 1574 -41 1613 -22
rect 1632 -28 1639 -27
rect 1638 -35 1639 -28
rect 1622 -38 1623 -35
rect 1638 -38 1651 -35
rect 1574 -42 1604 -41
rect 1613 -42 1619 -41
rect 1622 -42 1651 -38
rect 1541 -43 1651 -42
rect 1541 -44 1657 -43
rect 1216 -52 1267 -44
rect 1216 -64 1241 -52
rect 1248 -64 1267 -52
rect 1298 -52 1348 -44
rect 1298 -60 1314 -52
rect 1321 -54 1348 -52
rect 1357 -54 1578 -44
rect 1321 -64 1578 -54
rect 1607 -52 1657 -44
rect 1607 -61 1623 -52
rect 1216 -72 1267 -64
rect 1314 -72 1578 -64
rect 1604 -64 1623 -61
rect 1630 -64 1657 -52
rect 1604 -72 1657 -64
rect 1232 -80 1233 -72
rect 1248 -80 1261 -72
rect 1232 -88 1248 -80
rect 1229 -95 1248 -92
rect 1229 -104 1251 -95
rect 1202 -114 1251 -104
rect 1202 -120 1232 -114
rect 1251 -119 1256 -114
rect 1174 -136 1248 -120
rect 1266 -128 1296 -72
rect 1331 -82 1539 -72
rect 1574 -76 1619 -72
rect 1622 -73 1623 -72
rect 1638 -73 1651 -72
rect 1357 -112 1546 -82
rect 1372 -115 1546 -112
rect 1365 -118 1546 -115
rect 1174 -138 1187 -136
rect 1202 -138 1236 -136
rect 1174 -154 1248 -138
rect 1275 -142 1288 -128
rect 1303 -142 1319 -126
rect 1365 -131 1376 -118
rect 1158 -176 1159 -160
rect 1174 -176 1187 -154
rect 1202 -176 1232 -154
rect 1275 -158 1337 -142
rect 1365 -149 1376 -133
rect 1381 -138 1391 -118
rect 1401 -138 1415 -118
rect 1418 -131 1427 -118
rect 1443 -131 1452 -118
rect 1381 -149 1415 -138
rect 1418 -149 1427 -133
rect 1443 -149 1452 -133
rect 1459 -138 1469 -118
rect 1479 -138 1493 -118
rect 1494 -131 1505 -118
rect 1459 -149 1493 -138
rect 1494 -149 1505 -133
rect 1551 -142 1567 -126
rect 1574 -128 1604 -76
rect 1638 -80 1639 -73
rect 1623 -88 1639 -80
rect 1610 -120 1623 -101
rect 1638 -120 1668 -104
rect 1610 -136 1684 -120
rect 1610 -138 1623 -136
rect 1638 -138 1672 -136
rect 1275 -160 1288 -158
rect 1303 -160 1337 -158
rect 1275 -176 1337 -160
rect 1381 -165 1397 -162
rect 1459 -165 1489 -154
rect 1537 -158 1583 -142
rect 1610 -154 1684 -138
rect 1537 -160 1571 -158
rect 1536 -176 1583 -160
rect 1610 -176 1623 -154
rect 1638 -176 1668 -154
rect 1695 -176 1696 -160
rect 1711 -176 1724 -16
rect 1754 -120 1767 -16
rect 1812 -38 1813 -28
rect 1828 -38 1841 -28
rect 1812 -42 1841 -38
rect 1846 -42 1876 -16
rect 1894 -30 1910 -28
rect 1982 -30 2035 -16
rect 1983 -32 2047 -30
rect 2090 -32 2105 -16
rect 2154 -19 2184 -16
rect 2154 -22 2190 -19
rect 2120 -30 2136 -28
rect 1894 -42 1909 -38
rect 1812 -44 1909 -42
rect 1937 -44 2105 -32
rect 2121 -42 2136 -38
rect 2154 -41 2193 -22
rect 2212 -28 2219 -27
rect 2218 -35 2219 -28
rect 2202 -38 2203 -35
rect 2218 -38 2231 -35
rect 2154 -42 2184 -41
rect 2193 -42 2199 -41
rect 2202 -42 2231 -38
rect 2121 -43 2231 -42
rect 2121 -44 2237 -43
rect 1796 -52 1847 -44
rect 1796 -64 1821 -52
rect 1828 -64 1847 -52
rect 1878 -52 1928 -44
rect 1878 -60 1894 -52
rect 1901 -54 1928 -52
rect 1937 -54 2158 -44
rect 1901 -64 2158 -54
rect 2187 -52 2237 -44
rect 2187 -61 2203 -52
rect 1796 -72 1847 -64
rect 1894 -72 2158 -64
rect 2184 -64 2203 -61
rect 2210 -64 2237 -52
rect 2184 -72 2237 -64
rect 1812 -80 1813 -72
rect 1828 -80 1841 -72
rect 1812 -88 1828 -80
rect 1809 -95 1828 -92
rect 1809 -104 1831 -95
rect 1782 -114 1831 -104
rect 1782 -120 1812 -114
rect 1831 -119 1836 -114
rect 1754 -136 1828 -120
rect 1846 -128 1876 -72
rect 1911 -82 2119 -72
rect 2154 -76 2199 -72
rect 2202 -73 2203 -72
rect 2218 -73 2231 -72
rect 1937 -112 2126 -82
rect 1952 -115 2126 -112
rect 1945 -118 2126 -115
rect 1754 -138 1767 -136
rect 1782 -138 1816 -136
rect 1754 -154 1828 -138
rect 1855 -142 1868 -128
rect 1883 -142 1899 -126
rect 1945 -131 1956 -118
rect 1738 -176 1739 -160
rect 1754 -176 1767 -154
rect 1782 -176 1812 -154
rect 1855 -158 1917 -142
rect 1945 -149 1956 -133
rect 1961 -138 1971 -118
rect 1981 -138 1995 -118
rect 1998 -131 2007 -118
rect 2023 -131 2032 -118
rect 1961 -149 1995 -138
rect 1998 -149 2007 -133
rect 2023 -149 2032 -133
rect 2039 -138 2049 -118
rect 2059 -138 2073 -118
rect 2074 -131 2085 -118
rect 2039 -149 2073 -138
rect 2074 -149 2085 -133
rect 2131 -142 2147 -126
rect 2154 -128 2184 -76
rect 2218 -80 2219 -73
rect 2203 -88 2219 -80
rect 2190 -120 2203 -101
rect 2218 -120 2248 -104
rect 2190 -136 2264 -120
rect 2190 -138 2203 -136
rect 2218 -138 2252 -136
rect 1855 -160 1868 -158
rect 1883 -160 1917 -158
rect 1855 -176 1917 -160
rect 1961 -165 1977 -162
rect 2039 -165 2069 -154
rect 2117 -158 2163 -142
rect 2190 -154 2264 -138
rect 2117 -160 2151 -158
rect 2116 -176 2163 -160
rect 2190 -176 2203 -154
rect 2218 -176 2248 -154
rect 2275 -176 2276 -160
rect 2291 -176 2304 -16
rect 2334 -120 2347 -16
rect 2392 -38 2393 -28
rect 2408 -38 2421 -28
rect 2392 -42 2421 -38
rect 2426 -42 2456 -16
rect 2474 -30 2490 -28
rect 2562 -30 2615 -16
rect 2563 -32 2627 -30
rect 2670 -32 2685 -16
rect 2734 -19 2764 -16
rect 2734 -22 2770 -19
rect 2700 -30 2716 -28
rect 2474 -42 2489 -38
rect 2392 -44 2489 -42
rect 2517 -44 2685 -32
rect 2701 -42 2716 -38
rect 2734 -41 2773 -22
rect 2792 -28 2799 -27
rect 2798 -35 2799 -28
rect 2782 -38 2783 -35
rect 2798 -38 2811 -35
rect 2734 -42 2764 -41
rect 2773 -42 2779 -41
rect 2782 -42 2811 -38
rect 2701 -43 2811 -42
rect 2701 -44 2817 -43
rect 2376 -52 2427 -44
rect 2376 -64 2401 -52
rect 2408 -64 2427 -52
rect 2458 -52 2508 -44
rect 2458 -60 2474 -52
rect 2481 -54 2508 -52
rect 2517 -54 2738 -44
rect 2481 -64 2738 -54
rect 2767 -52 2817 -44
rect 2767 -61 2783 -52
rect 2376 -72 2427 -64
rect 2474 -72 2738 -64
rect 2764 -64 2783 -61
rect 2790 -64 2817 -52
rect 2764 -72 2817 -64
rect 2392 -80 2393 -72
rect 2408 -80 2421 -72
rect 2392 -88 2408 -80
rect 2389 -95 2408 -92
rect 2389 -104 2411 -95
rect 2362 -114 2411 -104
rect 2362 -120 2392 -114
rect 2411 -119 2416 -114
rect 2334 -136 2408 -120
rect 2426 -128 2456 -72
rect 2491 -82 2699 -72
rect 2734 -76 2779 -72
rect 2782 -73 2783 -72
rect 2798 -73 2811 -72
rect 2517 -112 2706 -82
rect 2532 -115 2706 -112
rect 2525 -118 2706 -115
rect 2334 -138 2347 -136
rect 2362 -138 2396 -136
rect 2334 -154 2408 -138
rect 2435 -142 2448 -128
rect 2463 -142 2479 -126
rect 2525 -131 2536 -118
rect 2318 -176 2319 -160
rect 2334 -176 2347 -154
rect 2362 -176 2392 -154
rect 2435 -158 2497 -142
rect 2525 -149 2536 -133
rect 2541 -138 2551 -118
rect 2561 -138 2575 -118
rect 2578 -131 2587 -118
rect 2603 -131 2612 -118
rect 2541 -149 2575 -138
rect 2578 -149 2587 -133
rect 2603 -149 2612 -133
rect 2619 -138 2629 -118
rect 2639 -138 2653 -118
rect 2654 -131 2665 -118
rect 2619 -149 2653 -138
rect 2654 -149 2665 -133
rect 2711 -142 2727 -126
rect 2734 -128 2764 -76
rect 2798 -80 2799 -73
rect 2783 -88 2799 -80
rect 2770 -120 2783 -101
rect 2798 -120 2828 -104
rect 2770 -136 2844 -120
rect 2770 -138 2783 -136
rect 2798 -138 2832 -136
rect 2435 -160 2448 -158
rect 2463 -160 2497 -158
rect 2435 -176 2497 -160
rect 2541 -165 2557 -162
rect 2619 -165 2649 -154
rect 2697 -158 2743 -142
rect 2770 -154 2844 -138
rect 2697 -160 2731 -158
rect 2696 -176 2743 -160
rect 2770 -176 2783 -154
rect 2798 -176 2828 -154
rect 2855 -176 2856 -160
rect 2871 -176 2884 -16
rect 2914 -120 2927 -16
rect 2972 -38 2973 -28
rect 2988 -38 3001 -28
rect 2972 -42 3001 -38
rect 3006 -42 3036 -16
rect 3054 -30 3070 -28
rect 3142 -30 3195 -16
rect 3143 -32 3205 -30
rect 3250 -32 3265 -16
rect 3314 -19 3344 -16
rect 3314 -22 3350 -19
rect 3280 -30 3296 -28
rect 3054 -42 3069 -38
rect 2972 -44 3069 -42
rect 3097 -44 3265 -32
rect 3281 -42 3296 -38
rect 3314 -41 3353 -22
rect 3372 -28 3379 -27
rect 3378 -35 3379 -28
rect 3362 -38 3363 -35
rect 3378 -38 3391 -35
rect 3314 -42 3344 -41
rect 3353 -42 3359 -41
rect 3362 -42 3391 -38
rect 3281 -43 3391 -42
rect 3281 -44 3397 -43
rect 2956 -52 3007 -44
rect 2956 -64 2981 -52
rect 2988 -64 3007 -52
rect 3038 -52 3088 -44
rect 3038 -60 3054 -52
rect 3061 -54 3088 -52
rect 3097 -54 3318 -44
rect 3061 -64 3318 -54
rect 3347 -52 3397 -44
rect 3347 -61 3363 -52
rect 2956 -72 3007 -64
rect 3054 -72 3318 -64
rect 3344 -64 3363 -61
rect 3370 -64 3397 -52
rect 3344 -72 3397 -64
rect 2972 -80 2973 -72
rect 2988 -80 3001 -72
rect 2972 -88 2988 -80
rect 2969 -95 2988 -92
rect 2969 -104 2991 -95
rect 2942 -114 2991 -104
rect 2942 -120 2972 -114
rect 2991 -119 2996 -114
rect 2914 -136 2988 -120
rect 3006 -128 3036 -72
rect 3071 -82 3279 -72
rect 3314 -76 3359 -72
rect 3362 -73 3363 -72
rect 3378 -73 3391 -72
rect 3097 -112 3286 -82
rect 3112 -115 3286 -112
rect 3105 -118 3286 -115
rect 2914 -138 2927 -136
rect 2942 -138 2976 -136
rect 2914 -154 2988 -138
rect 3015 -142 3028 -128
rect 3043 -142 3059 -126
rect 3105 -131 3116 -118
rect 2898 -176 2899 -160
rect 2914 -176 2927 -154
rect 2942 -176 2972 -154
rect 3015 -158 3077 -142
rect 3105 -149 3116 -133
rect 3121 -138 3131 -118
rect 3141 -138 3155 -118
rect 3158 -131 3167 -118
rect 3183 -131 3192 -118
rect 3121 -149 3155 -138
rect 3158 -149 3167 -133
rect 3183 -149 3192 -133
rect 3199 -138 3209 -118
rect 3219 -138 3233 -118
rect 3234 -131 3245 -118
rect 3199 -149 3233 -138
rect 3234 -149 3245 -133
rect 3291 -142 3307 -126
rect 3314 -128 3344 -76
rect 3378 -80 3379 -73
rect 3363 -88 3379 -80
rect 3350 -120 3363 -101
rect 3378 -120 3408 -104
rect 3350 -136 3424 -120
rect 3350 -138 3363 -136
rect 3378 -138 3412 -136
rect 3015 -160 3028 -158
rect 3043 -160 3077 -158
rect 3015 -176 3077 -160
rect 3121 -165 3137 -162
rect 3199 -165 3229 -154
rect 3277 -158 3323 -142
rect 3350 -154 3424 -138
rect 3277 -160 3311 -158
rect 3276 -176 3323 -160
rect 3350 -176 3363 -154
rect 3378 -176 3408 -154
rect 3435 -176 3436 -160
rect 3451 -176 3464 -16
rect 3494 -120 3507 -16
rect 3552 -38 3553 -28
rect 3568 -38 3581 -28
rect 3552 -42 3581 -38
rect 3586 -42 3616 -16
rect 3634 -30 3650 -28
rect 3722 -30 3775 -16
rect 3723 -32 3787 -30
rect 3830 -32 3845 -16
rect 3894 -19 3924 -16
rect 3894 -22 3930 -19
rect 3860 -30 3876 -28
rect 3634 -42 3649 -38
rect 3552 -44 3649 -42
rect 3677 -44 3845 -32
rect 3861 -42 3876 -38
rect 3894 -41 3933 -22
rect 3952 -28 3959 -27
rect 3958 -35 3959 -28
rect 3942 -38 3943 -35
rect 3958 -38 3971 -35
rect 3894 -42 3924 -41
rect 3933 -42 3939 -41
rect 3942 -42 3971 -38
rect 3861 -43 3971 -42
rect 3861 -44 3977 -43
rect 3536 -52 3587 -44
rect 3536 -64 3561 -52
rect 3568 -64 3587 -52
rect 3618 -52 3668 -44
rect 3618 -60 3634 -52
rect 3641 -54 3668 -52
rect 3677 -54 3898 -44
rect 3641 -64 3898 -54
rect 3927 -52 3977 -44
rect 3927 -61 3943 -52
rect 3536 -72 3587 -64
rect 3634 -72 3898 -64
rect 3924 -64 3943 -61
rect 3950 -64 3977 -52
rect 3924 -72 3977 -64
rect 3552 -80 3553 -72
rect 3568 -80 3581 -72
rect 3552 -88 3568 -80
rect 3549 -95 3568 -92
rect 3549 -104 3571 -95
rect 3522 -114 3571 -104
rect 3522 -120 3552 -114
rect 3571 -119 3576 -114
rect 3494 -136 3568 -120
rect 3586 -128 3616 -72
rect 3651 -82 3859 -72
rect 3894 -76 3939 -72
rect 3942 -73 3943 -72
rect 3958 -73 3971 -72
rect 3677 -112 3866 -82
rect 3692 -115 3866 -112
rect 3685 -118 3866 -115
rect 3494 -138 3507 -136
rect 3522 -138 3556 -136
rect 3494 -154 3568 -138
rect 3595 -142 3608 -128
rect 3623 -142 3639 -126
rect 3685 -131 3696 -118
rect 3478 -176 3479 -160
rect 3494 -176 3507 -154
rect 3522 -176 3552 -154
rect 3595 -158 3657 -142
rect 3685 -149 3696 -133
rect 3701 -138 3711 -118
rect 3721 -138 3735 -118
rect 3738 -131 3747 -118
rect 3763 -131 3772 -118
rect 3701 -149 3735 -138
rect 3738 -149 3747 -133
rect 3763 -149 3772 -133
rect 3779 -138 3789 -118
rect 3799 -138 3813 -118
rect 3814 -131 3825 -118
rect 3779 -149 3813 -138
rect 3814 -149 3825 -133
rect 3871 -142 3887 -126
rect 3894 -128 3924 -76
rect 3958 -80 3959 -73
rect 3943 -88 3959 -80
rect 3930 -120 3943 -101
rect 3958 -120 3988 -104
rect 3930 -136 4004 -120
rect 3930 -138 3943 -136
rect 3958 -138 3992 -136
rect 3595 -160 3608 -158
rect 3623 -160 3657 -158
rect 3595 -176 3657 -160
rect 3701 -165 3717 -162
rect 3779 -165 3809 -154
rect 3857 -158 3903 -142
rect 3930 -154 4004 -138
rect 3857 -160 3891 -158
rect 3856 -176 3903 -160
rect 3930 -176 3943 -154
rect 3958 -176 3988 -154
rect 4015 -176 4016 -160
rect 4031 -176 4044 -16
rect 4074 -120 4087 -16
rect 4132 -38 4133 -28
rect 4148 -38 4161 -28
rect 4132 -42 4161 -38
rect 4166 -42 4196 -16
rect 4214 -30 4230 -28
rect 4302 -30 4355 -16
rect 4303 -32 4367 -30
rect 4410 -32 4425 -16
rect 4474 -19 4504 -16
rect 4611 -17 6944 -16
rect 4474 -22 4510 -19
rect 4440 -30 4456 -28
rect 4214 -42 4229 -38
rect 4132 -44 4229 -42
rect 4257 -44 4425 -32
rect 4441 -42 4456 -38
rect 4474 -41 4513 -22
rect 4532 -28 4539 -27
rect 4538 -35 4539 -28
rect 4522 -38 4523 -35
rect 4538 -38 4551 -35
rect 4474 -42 4504 -41
rect 4513 -42 4519 -41
rect 4522 -42 4551 -38
rect 4441 -43 4551 -42
rect 4441 -44 4557 -43
rect 4116 -52 4167 -44
rect 4116 -64 4141 -52
rect 4148 -64 4167 -52
rect 4198 -52 4248 -44
rect 4198 -60 4214 -52
rect 4221 -54 4248 -52
rect 4257 -54 4478 -44
rect 4221 -64 4478 -54
rect 4507 -52 4557 -44
rect 4507 -61 4523 -52
rect 4116 -72 4167 -64
rect 4214 -72 4478 -64
rect 4504 -64 4523 -61
rect 4530 -64 4557 -52
rect 4504 -72 4557 -64
rect 4132 -80 4133 -72
rect 4148 -80 4161 -72
rect 4132 -88 4148 -80
rect 4129 -95 4148 -92
rect 4129 -104 4151 -95
rect 4102 -114 4151 -104
rect 4102 -120 4132 -114
rect 4151 -119 4156 -114
rect 4074 -136 4148 -120
rect 4166 -128 4196 -72
rect 4231 -82 4439 -72
rect 4474 -76 4519 -72
rect 4522 -73 4523 -72
rect 4538 -73 4551 -72
rect 4257 -112 4446 -82
rect 4272 -115 4446 -112
rect 4265 -118 4446 -115
rect 4074 -138 4087 -136
rect 4102 -138 4136 -136
rect 4074 -154 4148 -138
rect 4175 -142 4188 -128
rect 4203 -142 4219 -126
rect 4265 -131 4276 -118
rect 4058 -176 4059 -160
rect 4074 -176 4087 -154
rect 4102 -176 4132 -154
rect 4175 -158 4237 -142
rect 4265 -149 4276 -133
rect 4281 -138 4291 -118
rect 4301 -138 4315 -118
rect 4318 -131 4327 -118
rect 4343 -131 4352 -118
rect 4281 -149 4315 -138
rect 4318 -149 4327 -133
rect 4343 -149 4352 -133
rect 4359 -138 4369 -118
rect 4379 -138 4393 -118
rect 4394 -131 4405 -118
rect 4359 -149 4393 -138
rect 4394 -149 4405 -133
rect 4451 -142 4467 -126
rect 4474 -128 4504 -76
rect 4538 -80 4539 -73
rect 4523 -88 4539 -80
rect 4510 -120 4523 -101
rect 4538 -120 4568 -104
rect 4510 -136 4584 -120
rect 4510 -138 4523 -136
rect 4538 -138 4572 -136
rect 4175 -160 4188 -158
rect 4203 -160 4237 -158
rect 4175 -176 4237 -160
rect 4281 -165 4297 -162
rect 4359 -165 4389 -154
rect 4437 -158 4483 -142
rect 4510 -154 4584 -138
rect 4437 -160 4471 -158
rect 4436 -176 4483 -160
rect 4510 -176 4523 -154
rect 4538 -176 4568 -154
rect 4595 -176 4596 -160
rect 4611 -176 4624 -17
rect 4654 -121 4667 -17
rect 4712 -39 4713 -29
rect 4733 -31 4741 -29
rect 4731 -33 4741 -31
rect 4729 -35 4741 -33
rect 4728 -39 4741 -35
rect 4712 -43 4741 -39
rect 4746 -43 4776 -17
rect 4794 -31 4810 -29
rect 4882 -31 4933 -17
rect 4883 -33 4947 -31
rect 4990 -33 5005 -17
rect 5054 -20 5084 -17
rect 5054 -23 5090 -20
rect 5020 -31 5036 -29
rect 4794 -43 4809 -39
rect 4712 -45 4809 -43
rect 4837 -45 5005 -33
rect 5021 -43 5036 -39
rect 5054 -42 5093 -23
rect 5112 -29 5119 -28
rect 5118 -36 5119 -29
rect 5102 -39 5103 -36
rect 5118 -39 5131 -36
rect 5054 -43 5084 -42
rect 5093 -43 5099 -42
rect 5102 -43 5131 -39
rect 5021 -44 5131 -43
rect 5021 -45 5137 -44
rect 4696 -53 4747 -45
rect 4696 -65 4721 -53
rect 4728 -65 4747 -53
rect 4778 -53 4828 -45
rect 4778 -61 4794 -53
rect 4801 -55 4828 -53
rect 4837 -55 5058 -45
rect 4801 -65 5058 -55
rect 5087 -53 5137 -45
rect 5087 -62 5103 -53
rect 4696 -73 4747 -65
rect 4794 -73 5058 -65
rect 5084 -65 5103 -62
rect 5110 -65 5137 -53
rect 5084 -73 5137 -65
rect 4712 -81 4713 -73
rect 4728 -81 4741 -73
rect 4712 -89 4728 -81
rect 4709 -96 4728 -93
rect 4709 -105 4731 -96
rect 4682 -115 4731 -105
rect 4682 -121 4712 -115
rect 4731 -120 4736 -115
rect 4654 -137 4728 -121
rect 4746 -129 4776 -73
rect 4811 -83 5019 -73
rect 5054 -77 5099 -73
rect 5102 -74 5103 -73
rect 5118 -74 5131 -73
rect 4837 -113 5026 -83
rect 4852 -116 5026 -113
rect 4845 -119 5026 -116
rect 4654 -139 4667 -137
rect 4682 -139 4716 -137
rect 4654 -155 4728 -139
rect 4755 -143 4768 -129
rect 4783 -143 4799 -127
rect 4845 -132 4856 -119
rect -8 -184 33 -176
rect -8 -210 7 -184
rect 14 -210 33 -184
rect 97 -188 159 -176
rect 171 -188 246 -176
rect 304 -188 379 -176
rect 391 -188 422 -176
rect 428 -188 463 -176
rect 97 -190 259 -188
rect -8 -218 33 -210
rect 115 -214 128 -190
rect 143 -192 158 -190
rect -2 -228 -1 -218
rect 14 -228 27 -218
rect 42 -228 72 -214
rect 115 -228 158 -214
rect 182 -217 189 -210
rect 192 -214 259 -190
rect 291 -190 463 -188
rect 261 -212 289 -208
rect 291 -212 371 -190
rect 392 -192 407 -190
rect 261 -214 371 -212
rect 192 -218 371 -214
rect 165 -228 195 -218
rect 197 -228 350 -218
rect 358 -228 388 -218
rect 392 -228 422 -214
rect 450 -228 463 -190
rect 535 -184 570 -176
rect 535 -210 536 -184
rect 543 -210 570 -184
rect 478 -228 508 -214
rect 535 -218 570 -210
rect 572 -184 613 -176
rect 572 -210 587 -184
rect 594 -210 613 -184
rect 677 -188 739 -176
rect 751 -188 826 -176
rect 884 -188 959 -176
rect 971 -188 1002 -176
rect 1008 -188 1043 -176
rect 677 -190 839 -188
rect 572 -218 613 -210
rect 695 -214 708 -190
rect 723 -192 738 -190
rect 535 -228 536 -218
rect 551 -228 564 -218
rect 578 -228 579 -218
rect 594 -228 607 -218
rect 622 -228 652 -214
rect 695 -228 738 -214
rect 762 -217 769 -210
rect 772 -214 839 -190
rect 871 -190 1043 -188
rect 841 -212 869 -208
rect 871 -212 951 -190
rect 972 -192 987 -190
rect 841 -214 951 -212
rect 772 -218 951 -214
rect 745 -228 775 -218
rect 777 -228 930 -218
rect 938 -228 968 -218
rect 972 -228 1002 -214
rect 1030 -228 1043 -190
rect 1115 -184 1150 -176
rect 1115 -210 1116 -184
rect 1123 -210 1150 -184
rect 1058 -228 1088 -214
rect 1115 -218 1150 -210
rect 1152 -184 1193 -176
rect 1152 -210 1167 -184
rect 1174 -210 1193 -184
rect 1257 -188 1319 -176
rect 1331 -188 1406 -176
rect 1464 -188 1539 -176
rect 1551 -188 1582 -176
rect 1588 -188 1623 -176
rect 1257 -190 1419 -188
rect 1152 -218 1193 -210
rect 1275 -214 1288 -190
rect 1303 -192 1318 -190
rect 1115 -228 1116 -218
rect 1131 -228 1144 -218
rect 1158 -228 1159 -218
rect 1174 -228 1187 -218
rect 1202 -228 1232 -214
rect 1275 -228 1318 -214
rect 1342 -217 1349 -210
rect 1352 -214 1419 -190
rect 1451 -190 1623 -188
rect 1421 -212 1449 -208
rect 1451 -212 1531 -190
rect 1552 -192 1567 -190
rect 1421 -214 1531 -212
rect 1352 -218 1531 -214
rect 1325 -228 1355 -218
rect 1357 -228 1510 -218
rect 1518 -228 1548 -218
rect 1552 -228 1582 -214
rect 1610 -228 1623 -190
rect 1695 -184 1730 -176
rect 1695 -210 1696 -184
rect 1703 -210 1730 -184
rect 1638 -228 1668 -214
rect 1695 -218 1730 -210
rect 1732 -184 1773 -176
rect 1732 -210 1747 -184
rect 1754 -210 1773 -184
rect 1837 -188 1899 -176
rect 1911 -188 1986 -176
rect 2044 -188 2119 -176
rect 2131 -188 2162 -176
rect 2168 -188 2203 -176
rect 1837 -190 1999 -188
rect 1732 -218 1773 -210
rect 1855 -214 1868 -190
rect 1883 -192 1898 -190
rect 1695 -228 1696 -218
rect 1711 -228 1724 -218
rect 1738 -228 1739 -218
rect 1754 -228 1767 -218
rect 1782 -228 1812 -214
rect 1855 -228 1898 -214
rect 1922 -217 1929 -210
rect 1932 -214 1999 -190
rect 2031 -190 2203 -188
rect 2001 -212 2029 -208
rect 2031 -212 2111 -190
rect 2132 -192 2147 -190
rect 2001 -214 2111 -212
rect 1932 -218 2111 -214
rect 1905 -228 1935 -218
rect 1937 -228 2090 -218
rect 2098 -228 2128 -218
rect 2132 -228 2162 -214
rect 2190 -228 2203 -190
rect 2275 -184 2310 -176
rect 2275 -210 2276 -184
rect 2283 -210 2310 -184
rect 2218 -228 2248 -214
rect 2275 -218 2310 -210
rect 2312 -184 2353 -176
rect 2312 -210 2327 -184
rect 2334 -210 2353 -184
rect 2417 -188 2479 -176
rect 2491 -188 2566 -176
rect 2624 -188 2699 -176
rect 2711 -188 2742 -176
rect 2748 -188 2783 -176
rect 2417 -190 2579 -188
rect 2312 -218 2353 -210
rect 2435 -214 2448 -190
rect 2463 -192 2478 -190
rect 2275 -228 2276 -218
rect 2291 -228 2304 -218
rect 2318 -228 2319 -218
rect 2334 -228 2347 -218
rect 2362 -228 2392 -214
rect 2435 -228 2478 -214
rect 2502 -217 2509 -210
rect 2512 -214 2579 -190
rect 2611 -190 2783 -188
rect 2581 -212 2609 -208
rect 2611 -212 2691 -190
rect 2712 -192 2727 -190
rect 2581 -214 2691 -212
rect 2512 -218 2691 -214
rect 2485 -228 2515 -218
rect 2517 -228 2670 -218
rect 2678 -228 2708 -218
rect 2712 -228 2742 -214
rect 2770 -228 2783 -190
rect 2855 -184 2890 -176
rect 2855 -210 2856 -184
rect 2863 -210 2890 -184
rect 2798 -228 2828 -214
rect 2855 -218 2890 -210
rect 2892 -184 2933 -176
rect 2892 -210 2907 -184
rect 2914 -210 2933 -184
rect 2997 -188 3059 -176
rect 3071 -188 3146 -176
rect 3204 -188 3279 -176
rect 3291 -188 3322 -176
rect 3328 -188 3363 -176
rect 2997 -190 3159 -188
rect 2892 -218 2933 -210
rect 3015 -214 3028 -190
rect 3043 -192 3058 -190
rect 2855 -228 2856 -218
rect 2871 -228 2884 -218
rect 2898 -228 2899 -218
rect 2914 -228 2927 -218
rect 2942 -228 2972 -214
rect 3015 -228 3058 -214
rect 3082 -217 3089 -210
rect 3092 -214 3159 -190
rect 3191 -190 3363 -188
rect 3161 -212 3189 -208
rect 3191 -212 3271 -190
rect 3292 -192 3307 -190
rect 3161 -214 3271 -212
rect 3092 -218 3271 -214
rect 3065 -228 3095 -218
rect 3097 -228 3250 -218
rect 3258 -228 3288 -218
rect 3292 -228 3322 -214
rect 3350 -228 3363 -190
rect 3435 -184 3470 -176
rect 3435 -210 3436 -184
rect 3443 -210 3470 -184
rect 3378 -228 3408 -214
rect 3435 -218 3470 -210
rect 3472 -184 3513 -176
rect 3472 -210 3487 -184
rect 3494 -210 3513 -184
rect 3577 -188 3639 -176
rect 3651 -188 3726 -176
rect 3784 -188 3859 -176
rect 3871 -188 3902 -176
rect 3908 -188 3943 -176
rect 3577 -190 3739 -188
rect 3472 -218 3513 -210
rect 3595 -214 3608 -190
rect 3623 -192 3638 -190
rect 3435 -228 3436 -218
rect 3451 -228 3464 -218
rect 3478 -228 3479 -218
rect 3494 -228 3507 -218
rect 3522 -228 3552 -214
rect 3595 -228 3638 -214
rect 3662 -217 3669 -210
rect 3672 -214 3739 -190
rect 3771 -190 3943 -188
rect 3741 -212 3769 -208
rect 3771 -212 3851 -190
rect 3872 -192 3887 -190
rect 3741 -214 3851 -212
rect 3672 -218 3851 -214
rect 3645 -228 3675 -218
rect 3677 -228 3830 -218
rect 3838 -228 3868 -218
rect 3872 -228 3902 -214
rect 3930 -228 3943 -190
rect 4015 -184 4050 -176
rect 4015 -210 4016 -184
rect 4023 -210 4050 -184
rect 3958 -228 3988 -214
rect 4015 -218 4050 -210
rect 4052 -184 4093 -176
rect 4052 -210 4067 -184
rect 4074 -210 4093 -184
rect 4157 -188 4219 -176
rect 4231 -188 4306 -176
rect 4364 -188 4439 -176
rect 4451 -188 4482 -176
rect 4488 -188 4523 -176
rect 4157 -190 4319 -188
rect 4052 -218 4093 -210
rect 4175 -214 4188 -190
rect 4203 -192 4218 -190
rect 4015 -228 4016 -218
rect 4031 -228 4044 -218
rect 4058 -228 4059 -218
rect 4074 -228 4087 -218
rect 4102 -228 4132 -214
rect 4175 -228 4218 -214
rect 4242 -217 4249 -210
rect 4252 -214 4319 -190
rect 4351 -190 4523 -188
rect 4321 -212 4349 -208
rect 4351 -212 4431 -190
rect 4452 -192 4467 -190
rect 4321 -214 4431 -212
rect 4252 -218 4431 -214
rect 4225 -228 4255 -218
rect 4257 -228 4410 -218
rect 4418 -228 4448 -218
rect 4452 -228 4482 -214
rect 4510 -228 4523 -190
rect 4595 -184 4630 -176
rect 4638 -177 4639 -161
rect 4654 -177 4667 -155
rect 4682 -177 4712 -155
rect 4755 -159 4817 -143
rect 4845 -150 4856 -134
rect 4861 -139 4871 -119
rect 4881 -139 4895 -119
rect 4898 -132 4907 -119
rect 4923 -132 4932 -119
rect 4861 -150 4895 -139
rect 4898 -150 4907 -134
rect 4923 -150 4932 -134
rect 4939 -139 4949 -119
rect 4959 -139 4973 -119
rect 4974 -132 4985 -119
rect 4939 -150 4973 -139
rect 4974 -150 4985 -134
rect 5031 -143 5047 -127
rect 5054 -129 5084 -77
rect 5118 -81 5119 -74
rect 5103 -89 5119 -81
rect 5090 -121 5103 -102
rect 5118 -121 5148 -105
rect 5090 -137 5164 -121
rect 5090 -139 5103 -137
rect 5118 -139 5152 -137
rect 4755 -161 4768 -159
rect 4783 -161 4817 -159
rect 4755 -177 4817 -161
rect 4861 -166 4877 -163
rect 4939 -166 4969 -155
rect 5017 -159 5063 -143
rect 5090 -155 5164 -139
rect 5017 -161 5051 -159
rect 5016 -177 5063 -161
rect 5090 -177 5103 -155
rect 5118 -177 5148 -155
rect 5175 -177 5176 -161
rect 5191 -177 5204 -17
rect 5234 -121 5247 -17
rect 5292 -39 5293 -29
rect 5313 -31 5321 -29
rect 5311 -33 5321 -31
rect 5309 -35 5321 -33
rect 5308 -39 5321 -35
rect 5292 -43 5321 -39
rect 5326 -43 5356 -17
rect 5374 -31 5390 -29
rect 5462 -31 5513 -17
rect 5463 -33 5527 -31
rect 5570 -33 5585 -17
rect 5634 -20 5664 -17
rect 5634 -23 5670 -20
rect 5600 -31 5616 -29
rect 5374 -43 5389 -39
rect 5292 -45 5389 -43
rect 5417 -45 5585 -33
rect 5601 -43 5616 -39
rect 5634 -42 5673 -23
rect 5692 -29 5699 -28
rect 5698 -36 5699 -29
rect 5682 -39 5683 -36
rect 5698 -39 5711 -36
rect 5634 -43 5664 -42
rect 5673 -43 5679 -42
rect 5682 -43 5711 -39
rect 5601 -44 5711 -43
rect 5601 -45 5717 -44
rect 5276 -53 5327 -45
rect 5276 -65 5301 -53
rect 5308 -65 5327 -53
rect 5358 -53 5408 -45
rect 5358 -61 5374 -53
rect 5381 -55 5408 -53
rect 5417 -55 5638 -45
rect 5381 -65 5638 -55
rect 5667 -53 5717 -45
rect 5667 -62 5683 -53
rect 5276 -73 5327 -65
rect 5374 -73 5638 -65
rect 5664 -65 5683 -62
rect 5690 -65 5717 -53
rect 5664 -73 5717 -65
rect 5292 -81 5293 -73
rect 5308 -81 5321 -73
rect 5292 -89 5308 -81
rect 5289 -96 5308 -93
rect 5289 -105 5311 -96
rect 5262 -115 5311 -105
rect 5262 -121 5292 -115
rect 5311 -120 5316 -115
rect 5234 -137 5308 -121
rect 5326 -129 5356 -73
rect 5391 -83 5599 -73
rect 5634 -77 5679 -73
rect 5682 -74 5683 -73
rect 5698 -74 5711 -73
rect 5417 -113 5606 -83
rect 5432 -116 5606 -113
rect 5425 -119 5606 -116
rect 5234 -139 5247 -137
rect 5262 -139 5296 -137
rect 5234 -155 5308 -139
rect 5335 -143 5348 -129
rect 5363 -143 5379 -127
rect 5425 -132 5436 -119
rect 5218 -177 5219 -161
rect 5234 -177 5247 -155
rect 5262 -177 5292 -155
rect 5335 -159 5397 -143
rect 5425 -150 5436 -134
rect 5441 -139 5451 -119
rect 5461 -139 5475 -119
rect 5478 -132 5487 -119
rect 5503 -132 5512 -119
rect 5441 -150 5475 -139
rect 5478 -150 5487 -134
rect 5503 -150 5512 -134
rect 5519 -139 5529 -119
rect 5539 -139 5553 -119
rect 5554 -132 5565 -119
rect 5519 -150 5553 -139
rect 5554 -150 5565 -134
rect 5611 -143 5627 -127
rect 5634 -129 5664 -77
rect 5698 -81 5699 -74
rect 5683 -89 5699 -81
rect 5670 -121 5683 -102
rect 5698 -121 5728 -105
rect 5670 -137 5744 -121
rect 5670 -139 5683 -137
rect 5698 -139 5732 -137
rect 5335 -161 5348 -159
rect 5363 -161 5397 -159
rect 5335 -177 5397 -161
rect 5441 -166 5457 -163
rect 5519 -166 5549 -155
rect 5597 -159 5643 -143
rect 5670 -155 5744 -139
rect 5597 -161 5631 -159
rect 5596 -177 5643 -161
rect 5670 -177 5683 -155
rect 5698 -177 5728 -155
rect 5755 -177 5756 -161
rect 5771 -177 5784 -17
rect 5814 -121 5827 -17
rect 5872 -39 5873 -29
rect 5893 -31 5901 -29
rect 5891 -33 5901 -31
rect 5889 -35 5901 -33
rect 5888 -39 5901 -35
rect 5872 -43 5901 -39
rect 5906 -43 5936 -17
rect 5954 -31 5970 -29
rect 6042 -31 6093 -17
rect 6043 -33 6107 -31
rect 6150 -33 6165 -17
rect 6214 -20 6244 -17
rect 6214 -23 6250 -20
rect 6180 -31 6196 -29
rect 5954 -43 5969 -39
rect 5872 -45 5969 -43
rect 5997 -45 6165 -33
rect 6181 -43 6196 -39
rect 6214 -42 6253 -23
rect 6272 -29 6279 -28
rect 6278 -36 6279 -29
rect 6262 -39 6263 -36
rect 6278 -39 6291 -36
rect 6214 -43 6244 -42
rect 6253 -43 6259 -42
rect 6262 -43 6291 -39
rect 6181 -44 6291 -43
rect 6181 -45 6297 -44
rect 5856 -53 5907 -45
rect 5856 -65 5881 -53
rect 5888 -65 5907 -53
rect 5938 -53 5988 -45
rect 5938 -61 5954 -53
rect 5961 -55 5988 -53
rect 5997 -55 6218 -45
rect 5961 -65 6218 -55
rect 6247 -53 6297 -45
rect 6247 -62 6263 -53
rect 5856 -73 5907 -65
rect 5954 -73 6218 -65
rect 6244 -65 6263 -62
rect 6270 -65 6297 -53
rect 6244 -73 6297 -65
rect 5872 -81 5873 -73
rect 5888 -81 5901 -73
rect 5872 -89 5888 -81
rect 5869 -96 5888 -93
rect 5869 -105 5891 -96
rect 5842 -115 5891 -105
rect 5842 -121 5872 -115
rect 5891 -120 5896 -115
rect 5814 -137 5888 -121
rect 5906 -129 5936 -73
rect 5971 -83 6179 -73
rect 6214 -77 6259 -73
rect 6262 -74 6263 -73
rect 6278 -74 6291 -73
rect 5997 -113 6186 -83
rect 6012 -116 6186 -113
rect 6005 -119 6186 -116
rect 5814 -139 5827 -137
rect 5842 -139 5876 -137
rect 5814 -155 5888 -139
rect 5915 -143 5928 -129
rect 5943 -143 5959 -127
rect 6005 -132 6016 -119
rect 5798 -177 5799 -161
rect 5814 -177 5827 -155
rect 5842 -177 5872 -155
rect 5915 -159 5977 -143
rect 6005 -150 6016 -134
rect 6021 -139 6031 -119
rect 6041 -139 6055 -119
rect 6058 -132 6067 -119
rect 6083 -132 6092 -119
rect 6021 -150 6055 -139
rect 6058 -150 6067 -134
rect 6083 -150 6092 -134
rect 6099 -139 6109 -119
rect 6119 -139 6133 -119
rect 6134 -132 6145 -119
rect 6099 -150 6133 -139
rect 6134 -150 6145 -134
rect 6191 -143 6207 -127
rect 6214 -129 6244 -77
rect 6278 -81 6279 -74
rect 6263 -89 6279 -81
rect 6250 -121 6263 -102
rect 6278 -121 6308 -105
rect 6250 -137 6324 -121
rect 6250 -139 6263 -137
rect 6278 -139 6312 -137
rect 5915 -161 5928 -159
rect 5943 -161 5977 -159
rect 5915 -177 5977 -161
rect 6021 -166 6037 -163
rect 6099 -166 6129 -155
rect 6177 -159 6223 -143
rect 6250 -155 6324 -139
rect 6177 -161 6211 -159
rect 6176 -177 6223 -161
rect 6250 -177 6263 -155
rect 6278 -177 6308 -155
rect 6335 -177 6336 -161
rect 6351 -177 6364 -17
rect 6394 -121 6407 -17
rect 6452 -39 6453 -29
rect 6473 -31 6481 -29
rect 6471 -33 6481 -31
rect 6469 -35 6481 -33
rect 6468 -39 6481 -35
rect 6452 -43 6481 -39
rect 6486 -43 6516 -17
rect 6534 -31 6550 -29
rect 6622 -31 6673 -17
rect 6623 -33 6687 -31
rect 6730 -33 6745 -17
rect 6794 -20 6824 -17
rect 6794 -23 6830 -20
rect 6760 -31 6776 -29
rect 6534 -43 6549 -39
rect 6452 -45 6549 -43
rect 6577 -45 6745 -33
rect 6761 -43 6776 -39
rect 6794 -42 6833 -23
rect 6852 -29 6859 -28
rect 6858 -36 6859 -29
rect 6842 -39 6843 -36
rect 6858 -39 6871 -36
rect 6794 -43 6824 -42
rect 6833 -43 6839 -42
rect 6842 -43 6871 -39
rect 6761 -44 6871 -43
rect 6761 -45 6877 -44
rect 6436 -53 6487 -45
rect 6436 -65 6461 -53
rect 6468 -65 6487 -53
rect 6518 -53 6568 -45
rect 6518 -61 6534 -53
rect 6541 -55 6568 -53
rect 6577 -55 6798 -45
rect 6541 -65 6798 -55
rect 6827 -53 6877 -45
rect 6827 -62 6843 -53
rect 6436 -73 6487 -65
rect 6534 -73 6798 -65
rect 6824 -65 6843 -62
rect 6850 -65 6877 -53
rect 6824 -73 6877 -65
rect 6452 -81 6453 -73
rect 6468 -81 6481 -73
rect 6452 -89 6468 -81
rect 6449 -96 6468 -93
rect 6449 -105 6471 -96
rect 6422 -115 6471 -105
rect 6422 -121 6452 -115
rect 6471 -120 6476 -115
rect 6394 -137 6468 -121
rect 6486 -129 6516 -73
rect 6551 -83 6759 -73
rect 6794 -77 6839 -73
rect 6842 -74 6843 -73
rect 6858 -74 6871 -73
rect 6577 -113 6766 -83
rect 6592 -116 6766 -113
rect 6585 -119 6766 -116
rect 6394 -139 6407 -137
rect 6422 -139 6456 -137
rect 6394 -155 6468 -139
rect 6495 -143 6508 -129
rect 6523 -143 6539 -127
rect 6585 -132 6596 -119
rect 6378 -177 6379 -161
rect 6394 -177 6407 -155
rect 6422 -177 6452 -155
rect 6495 -159 6557 -143
rect 6585 -150 6596 -134
rect 6601 -139 6611 -119
rect 6621 -139 6635 -119
rect 6638 -132 6647 -119
rect 6663 -132 6672 -119
rect 6601 -150 6635 -139
rect 6638 -150 6647 -134
rect 6663 -150 6672 -134
rect 6679 -139 6689 -119
rect 6699 -139 6713 -119
rect 6714 -132 6725 -119
rect 6679 -150 6713 -139
rect 6714 -150 6725 -134
rect 6771 -143 6787 -127
rect 6794 -129 6824 -77
rect 6858 -81 6859 -74
rect 6843 -89 6859 -81
rect 6830 -121 6843 -102
rect 6858 -121 6888 -105
rect 6830 -137 6904 -121
rect 6830 -139 6843 -137
rect 6858 -139 6892 -137
rect 6495 -161 6508 -159
rect 6523 -161 6557 -159
rect 6495 -177 6557 -161
rect 6601 -166 6617 -163
rect 6679 -166 6709 -155
rect 6757 -159 6803 -143
rect 6830 -155 6904 -139
rect 6757 -161 6791 -159
rect 6756 -177 6803 -161
rect 6830 -177 6843 -155
rect 6858 -177 6888 -155
rect 6915 -177 6916 -161
rect 6931 -177 6944 -17
rect 4595 -210 4596 -184
rect 4603 -210 4630 -184
rect 4538 -228 4568 -214
rect 4595 -218 4630 -210
rect 4632 -185 4673 -177
rect 4632 -211 4647 -185
rect 4654 -211 4673 -185
rect 4737 -189 4799 -177
rect 4811 -189 4886 -177
rect 4944 -189 5019 -177
rect 5031 -189 5062 -177
rect 5068 -189 5103 -177
rect 4737 -191 4899 -189
rect 4595 -228 4596 -218
rect 4611 -228 4624 -218
rect 4632 -219 4673 -211
rect 4755 -215 4768 -191
rect 4783 -193 4798 -191
rect 4832 -209 4899 -191
rect 4931 -191 5103 -189
rect 4931 -209 5011 -191
rect 5032 -193 5047 -191
rect -2 -229 4624 -228
rect 4638 -229 4639 -219
rect 4654 -229 4667 -219
rect 4682 -229 4712 -215
rect 4755 -229 4798 -215
rect 4822 -218 4829 -211
rect 4832 -219 5011 -209
rect 4805 -229 4835 -219
rect 4837 -229 4990 -219
rect 4998 -229 5028 -219
rect 5032 -229 5062 -215
rect 5090 -229 5103 -191
rect 5175 -185 5210 -177
rect 5175 -211 5176 -185
rect 5183 -211 5210 -185
rect 5118 -229 5148 -215
rect 5175 -219 5210 -211
rect 5212 -185 5253 -177
rect 5212 -211 5227 -185
rect 5234 -211 5253 -185
rect 5317 -189 5379 -177
rect 5391 -189 5466 -177
rect 5524 -189 5599 -177
rect 5611 -189 5642 -177
rect 5648 -189 5683 -177
rect 5317 -191 5479 -189
rect 5212 -219 5253 -211
rect 5335 -215 5348 -191
rect 5363 -193 5378 -191
rect 5412 -209 5479 -191
rect 5511 -191 5683 -189
rect 5511 -209 5591 -191
rect 5612 -193 5627 -191
rect 5175 -229 5176 -219
rect 5191 -229 5204 -219
rect 5218 -229 5219 -219
rect 5234 -229 5247 -219
rect 5262 -229 5292 -215
rect 5335 -229 5378 -215
rect 5402 -218 5409 -211
rect 5412 -219 5591 -209
rect 5385 -229 5415 -219
rect 5417 -229 5570 -219
rect 5578 -229 5608 -219
rect 5612 -229 5642 -215
rect 5670 -229 5683 -191
rect 5755 -185 5790 -177
rect 5755 -211 5756 -185
rect 5763 -211 5790 -185
rect 5698 -229 5728 -215
rect 5755 -219 5790 -211
rect 5792 -185 5833 -177
rect 5792 -211 5807 -185
rect 5814 -211 5833 -185
rect 5897 -189 5959 -177
rect 5971 -189 6046 -177
rect 6104 -189 6179 -177
rect 6191 -189 6222 -177
rect 6228 -189 6263 -177
rect 5897 -191 6059 -189
rect 5792 -219 5833 -211
rect 5915 -215 5928 -191
rect 5943 -193 5958 -191
rect 5992 -209 6059 -191
rect 6091 -191 6263 -189
rect 6091 -209 6171 -191
rect 6192 -193 6207 -191
rect 5755 -229 5756 -219
rect 5771 -229 5784 -219
rect 5798 -229 5799 -219
rect 5814 -229 5827 -219
rect 5842 -229 5872 -215
rect 5915 -229 5958 -215
rect 5982 -218 5989 -211
rect 5992 -219 6171 -209
rect 5965 -229 5995 -219
rect 5997 -229 6150 -219
rect 6158 -229 6188 -219
rect 6192 -229 6222 -215
rect 6250 -229 6263 -191
rect 6335 -185 6370 -177
rect 6335 -211 6336 -185
rect 6343 -211 6370 -185
rect 6278 -229 6308 -215
rect 6335 -219 6370 -211
rect 6372 -185 6413 -177
rect 6372 -211 6387 -185
rect 6394 -211 6413 -185
rect 6477 -189 6539 -177
rect 6551 -189 6626 -177
rect 6684 -189 6759 -177
rect 6771 -189 6802 -177
rect 6808 -189 6843 -177
rect 6477 -191 6639 -189
rect 6372 -219 6413 -211
rect 6495 -215 6508 -191
rect 6523 -193 6538 -191
rect 6572 -209 6639 -191
rect 6671 -191 6843 -189
rect 6671 -209 6751 -191
rect 6772 -193 6787 -191
rect 6335 -229 6336 -219
rect 6351 -229 6364 -219
rect 6378 -229 6379 -219
rect 6394 -229 6407 -219
rect 6422 -229 6452 -215
rect 6495 -229 6538 -215
rect 6562 -218 6569 -211
rect 6572 -219 6751 -209
rect 6545 -229 6575 -219
rect 6577 -229 6730 -219
rect 6738 -229 6768 -219
rect 6772 -229 6802 -215
rect 6830 -229 6843 -191
rect 6915 -185 6950 -177
rect 6915 -211 6916 -185
rect 6923 -211 6950 -185
rect 6858 -229 6888 -215
rect 6915 -219 6950 -211
rect 6915 -229 6916 -219
rect 6931 -229 6944 -219
rect -2 -234 6944 -229
rect -1 -242 6944 -234
rect 14 -272 27 -242
rect 42 -260 72 -242
rect 115 -256 129 -242
rect 165 -256 385 -242
rect 116 -258 129 -256
rect 82 -270 97 -258
rect 79 -272 101 -270
rect 106 -272 136 -258
rect 197 -260 350 -256
rect 179 -272 371 -260
rect 414 -272 444 -258
rect 450 -272 463 -242
rect 478 -260 508 -242
rect 551 -272 564 -242
rect 594 -272 607 -242
rect 622 -260 652 -242
rect 695 -256 709 -242
rect 745 -256 965 -242
rect 696 -258 709 -256
rect 662 -270 677 -258
rect 659 -272 681 -270
rect 686 -272 716 -258
rect 777 -260 930 -256
rect 759 -272 951 -260
rect 994 -272 1024 -258
rect 1030 -272 1043 -242
rect 1058 -260 1088 -242
rect 1131 -272 1144 -242
rect 1174 -272 1187 -242
rect 1202 -260 1232 -242
rect 1275 -256 1289 -242
rect 1325 -256 1545 -242
rect 1276 -258 1289 -256
rect 1242 -270 1257 -258
rect 1239 -272 1261 -270
rect 1266 -272 1296 -258
rect 1357 -260 1510 -256
rect 1339 -272 1531 -260
rect 1574 -272 1604 -258
rect 1610 -272 1623 -242
rect 1638 -260 1668 -242
rect 1711 -272 1724 -242
rect 1754 -272 1767 -242
rect 1782 -260 1812 -242
rect 1855 -256 1869 -242
rect 1905 -256 2125 -242
rect 1856 -258 1869 -256
rect 1822 -270 1837 -258
rect 1819 -272 1841 -270
rect 1846 -272 1876 -258
rect 1937 -260 2090 -256
rect 1919 -272 2111 -260
rect 2154 -272 2184 -258
rect 2190 -272 2203 -242
rect 2218 -260 2248 -242
rect 2291 -272 2304 -242
rect 2334 -272 2347 -242
rect 2362 -260 2392 -242
rect 2435 -256 2449 -242
rect 2485 -256 2705 -242
rect 2436 -258 2449 -256
rect 2402 -270 2417 -258
rect 2399 -272 2421 -270
rect 2426 -272 2456 -258
rect 2517 -260 2670 -256
rect 2499 -272 2691 -260
rect 2734 -272 2764 -258
rect 2770 -272 2783 -242
rect 2798 -260 2828 -242
rect 2871 -272 2884 -242
rect 2914 -272 2927 -242
rect 2942 -260 2972 -242
rect 3015 -256 3029 -242
rect 3065 -256 3285 -242
rect 3016 -258 3029 -256
rect 2982 -270 2997 -258
rect 2979 -272 3001 -270
rect 3006 -272 3036 -258
rect 3097 -260 3250 -256
rect 3079 -272 3271 -260
rect 3314 -272 3344 -258
rect 3350 -272 3363 -242
rect 3378 -260 3408 -242
rect 3451 -272 3464 -242
rect 3494 -272 3507 -242
rect 3522 -260 3552 -242
rect 3595 -256 3609 -242
rect 3645 -256 3865 -242
rect 3596 -258 3609 -256
rect 3562 -270 3577 -258
rect 3559 -272 3581 -270
rect 3586 -272 3616 -258
rect 3677 -260 3830 -256
rect 3659 -272 3851 -260
rect 3894 -272 3924 -258
rect 3930 -272 3943 -242
rect 3958 -260 3988 -242
rect 4031 -272 4044 -242
rect 4074 -272 4087 -242
rect 4102 -260 4132 -242
rect 4175 -256 4189 -242
rect 4225 -256 4445 -242
rect 4176 -258 4189 -256
rect 4142 -270 4157 -258
rect 4139 -272 4161 -270
rect 4166 -272 4196 -258
rect 4257 -260 4410 -256
rect 4239 -272 4431 -260
rect 4474 -272 4504 -258
rect 4510 -272 4523 -242
rect 4538 -260 4568 -242
rect 4611 -243 6944 -242
rect 4611 -272 4624 -243
rect -1 -273 4624 -272
rect 4654 -273 4667 -243
rect 4682 -261 4712 -243
rect 4755 -257 4769 -243
rect 4805 -257 5025 -243
rect 4756 -259 4769 -257
rect 4722 -271 4737 -259
rect 4719 -273 4741 -271
rect 4746 -273 4776 -259
rect 4837 -261 4990 -257
rect 4819 -273 5011 -261
rect 5054 -273 5084 -259
rect 5090 -273 5103 -243
rect 5118 -261 5148 -243
rect 5191 -273 5204 -243
rect 5234 -273 5247 -243
rect 5262 -261 5292 -243
rect 5335 -257 5349 -243
rect 5385 -257 5605 -243
rect 5336 -259 5349 -257
rect 5302 -271 5317 -259
rect 5299 -273 5321 -271
rect 5326 -273 5356 -259
rect 5417 -261 5570 -257
rect 5399 -273 5591 -261
rect 5634 -273 5664 -259
rect 5670 -273 5683 -243
rect 5698 -261 5728 -243
rect 5771 -273 5784 -243
rect 5814 -273 5827 -243
rect 5842 -261 5872 -243
rect 5915 -257 5929 -243
rect 5965 -257 6185 -243
rect 5916 -259 5929 -257
rect 5882 -271 5897 -259
rect 5879 -273 5901 -271
rect 5906 -273 5936 -259
rect 5997 -261 6150 -257
rect 5979 -273 6171 -261
rect 6214 -273 6244 -259
rect 6250 -273 6263 -243
rect 6278 -261 6308 -243
rect 6351 -273 6364 -243
rect 6394 -273 6407 -243
rect 6422 -261 6452 -243
rect 6495 -257 6509 -243
rect 6545 -257 6765 -243
rect 6496 -259 6509 -257
rect 6462 -271 6477 -259
rect 6459 -273 6481 -271
rect 6486 -273 6516 -259
rect 6577 -261 6730 -257
rect 6559 -273 6751 -261
rect 6794 -273 6824 -259
rect 6830 -273 6843 -243
rect 6858 -261 6888 -243
rect 6931 -273 6944 -243
rect -1 -286 6944 -273
rect 14 -390 27 -286
rect 72 -308 73 -298
rect 88 -308 101 -298
rect 72 -312 101 -308
rect 106 -312 136 -286
rect 154 -300 170 -298
rect 242 -300 295 -286
rect 243 -302 307 -300
rect 350 -302 365 -286
rect 414 -289 444 -286
rect 414 -292 450 -289
rect 380 -300 396 -298
rect 154 -312 169 -308
rect 72 -314 169 -312
rect 197 -314 365 -302
rect 381 -312 396 -308
rect 414 -311 453 -292
rect 472 -298 479 -297
rect 478 -305 479 -298
rect 462 -308 463 -305
rect 478 -308 491 -305
rect 414 -312 444 -311
rect 453 -312 459 -311
rect 462 -312 491 -308
rect 381 -313 491 -312
rect 381 -314 497 -313
rect 56 -322 107 -314
rect 56 -334 81 -322
rect 88 -334 107 -322
rect 138 -322 188 -314
rect 138 -330 154 -322
rect 161 -324 188 -322
rect 197 -324 418 -314
rect 161 -334 418 -324
rect 447 -322 497 -314
rect 447 -331 463 -322
rect 56 -342 107 -334
rect 154 -342 418 -334
rect 444 -334 463 -331
rect 470 -334 497 -322
rect 444 -342 497 -334
rect 72 -350 73 -342
rect 88 -350 101 -342
rect 72 -358 88 -350
rect 69 -365 88 -362
rect 69 -374 91 -365
rect 42 -384 91 -374
rect 42 -390 72 -384
rect 91 -389 96 -384
rect 14 -406 88 -390
rect 106 -398 136 -342
rect 171 -352 379 -342
rect 414 -346 459 -342
rect 462 -343 463 -342
rect 478 -343 491 -342
rect 197 -382 386 -352
rect 212 -385 386 -382
rect 205 -388 386 -385
rect 14 -408 27 -406
rect 42 -408 76 -406
rect 14 -424 88 -408
rect 115 -412 128 -398
rect 143 -412 159 -396
rect 205 -401 216 -388
rect -2 -446 -1 -430
rect 14 -446 27 -424
rect 42 -446 72 -424
rect 115 -428 177 -412
rect 205 -419 216 -403
rect 221 -408 231 -388
rect 241 -408 255 -388
rect 258 -401 267 -388
rect 283 -401 292 -388
rect 221 -419 255 -408
rect 258 -419 267 -403
rect 283 -419 292 -403
rect 299 -408 309 -388
rect 319 -408 333 -388
rect 334 -401 345 -388
rect 299 -419 333 -408
rect 334 -419 345 -403
rect 391 -412 407 -396
rect 414 -398 444 -346
rect 478 -350 479 -343
rect 463 -358 479 -350
rect 450 -390 463 -371
rect 478 -390 508 -374
rect 450 -406 524 -390
rect 450 -408 463 -406
rect 478 -408 512 -406
rect 115 -430 128 -428
rect 143 -430 177 -428
rect 115 -446 177 -430
rect 221 -435 237 -432
rect 299 -435 329 -424
rect 377 -428 423 -412
rect 450 -424 524 -408
rect 377 -430 411 -428
rect 376 -446 423 -430
rect 450 -446 463 -424
rect 478 -446 508 -424
rect 535 -446 536 -430
rect 551 -446 564 -286
rect 594 -390 607 -286
rect 652 -308 653 -298
rect 668 -308 681 -298
rect 652 -312 681 -308
rect 686 -312 716 -286
rect 734 -300 750 -298
rect 822 -300 875 -286
rect 823 -302 887 -300
rect 930 -302 945 -286
rect 994 -289 1024 -286
rect 994 -292 1030 -289
rect 960 -300 976 -298
rect 734 -312 749 -308
rect 652 -314 749 -312
rect 777 -314 945 -302
rect 961 -312 976 -308
rect 994 -311 1033 -292
rect 1052 -298 1059 -297
rect 1058 -305 1059 -298
rect 1042 -308 1043 -305
rect 1058 -308 1071 -305
rect 994 -312 1024 -311
rect 1033 -312 1039 -311
rect 1042 -312 1071 -308
rect 961 -313 1071 -312
rect 961 -314 1077 -313
rect 636 -322 687 -314
rect 636 -334 661 -322
rect 668 -334 687 -322
rect 718 -322 768 -314
rect 718 -330 734 -322
rect 741 -324 768 -322
rect 777 -324 998 -314
rect 741 -334 998 -324
rect 1027 -322 1077 -314
rect 1027 -331 1043 -322
rect 636 -342 687 -334
rect 734 -342 998 -334
rect 1024 -334 1043 -331
rect 1050 -334 1077 -322
rect 1024 -342 1077 -334
rect 652 -350 653 -342
rect 668 -350 681 -342
rect 652 -358 668 -350
rect 649 -365 668 -362
rect 649 -374 671 -365
rect 622 -384 671 -374
rect 622 -390 652 -384
rect 671 -389 676 -384
rect 594 -406 668 -390
rect 686 -398 716 -342
rect 751 -352 959 -342
rect 994 -346 1039 -342
rect 1042 -343 1043 -342
rect 1058 -343 1071 -342
rect 777 -382 966 -352
rect 792 -385 966 -382
rect 785 -388 966 -385
rect 594 -408 607 -406
rect 622 -408 656 -406
rect 594 -424 668 -408
rect 695 -412 708 -398
rect 723 -412 739 -396
rect 785 -401 796 -388
rect 578 -446 579 -430
rect 594 -446 607 -424
rect 622 -446 652 -424
rect 695 -428 757 -412
rect 785 -419 796 -403
rect 801 -408 811 -388
rect 821 -408 835 -388
rect 838 -401 847 -388
rect 863 -401 872 -388
rect 801 -419 835 -408
rect 838 -419 847 -403
rect 863 -419 872 -403
rect 879 -408 889 -388
rect 899 -408 913 -388
rect 914 -401 925 -388
rect 879 -419 913 -408
rect 914 -419 925 -403
rect 971 -412 987 -396
rect 994 -398 1024 -346
rect 1058 -350 1059 -343
rect 1043 -358 1059 -350
rect 1030 -390 1043 -371
rect 1058 -390 1088 -374
rect 1030 -406 1104 -390
rect 1030 -408 1043 -406
rect 1058 -408 1092 -406
rect 695 -430 708 -428
rect 723 -430 757 -428
rect 695 -446 757 -430
rect 801 -435 817 -432
rect 879 -435 909 -424
rect 957 -428 1003 -412
rect 1030 -424 1104 -408
rect 957 -430 991 -428
rect 956 -446 1003 -430
rect 1030 -446 1043 -424
rect 1058 -446 1088 -424
rect 1115 -446 1116 -430
rect 1131 -446 1144 -286
rect 1174 -390 1187 -286
rect 1232 -308 1233 -298
rect 1248 -308 1261 -298
rect 1232 -312 1261 -308
rect 1266 -312 1296 -286
rect 1314 -300 1330 -298
rect 1402 -300 1455 -286
rect 1403 -302 1467 -300
rect 1510 -302 1525 -286
rect 1574 -289 1604 -286
rect 1574 -292 1610 -289
rect 1540 -300 1556 -298
rect 1314 -312 1329 -308
rect 1232 -314 1329 -312
rect 1357 -314 1525 -302
rect 1541 -312 1556 -308
rect 1574 -311 1613 -292
rect 1632 -298 1639 -297
rect 1638 -305 1639 -298
rect 1622 -308 1623 -305
rect 1638 -308 1651 -305
rect 1574 -312 1604 -311
rect 1613 -312 1619 -311
rect 1622 -312 1651 -308
rect 1541 -313 1651 -312
rect 1541 -314 1657 -313
rect 1216 -322 1267 -314
rect 1216 -334 1241 -322
rect 1248 -334 1267 -322
rect 1298 -322 1348 -314
rect 1298 -330 1314 -322
rect 1321 -324 1348 -322
rect 1357 -324 1578 -314
rect 1321 -334 1578 -324
rect 1607 -322 1657 -314
rect 1607 -331 1623 -322
rect 1216 -342 1267 -334
rect 1314 -342 1578 -334
rect 1604 -334 1623 -331
rect 1630 -334 1657 -322
rect 1604 -342 1657 -334
rect 1232 -350 1233 -342
rect 1248 -350 1261 -342
rect 1232 -358 1248 -350
rect 1229 -365 1248 -362
rect 1229 -374 1251 -365
rect 1202 -384 1251 -374
rect 1202 -390 1232 -384
rect 1251 -389 1256 -384
rect 1174 -406 1248 -390
rect 1266 -398 1296 -342
rect 1331 -352 1539 -342
rect 1574 -346 1619 -342
rect 1622 -343 1623 -342
rect 1638 -343 1651 -342
rect 1357 -382 1546 -352
rect 1372 -385 1546 -382
rect 1365 -388 1546 -385
rect 1174 -408 1187 -406
rect 1202 -408 1236 -406
rect 1174 -424 1248 -408
rect 1275 -412 1288 -398
rect 1303 -412 1319 -396
rect 1365 -401 1376 -388
rect 1158 -446 1159 -430
rect 1174 -446 1187 -424
rect 1202 -446 1232 -424
rect 1275 -428 1337 -412
rect 1365 -419 1376 -403
rect 1381 -408 1391 -388
rect 1401 -408 1415 -388
rect 1418 -401 1427 -388
rect 1443 -401 1452 -388
rect 1381 -419 1415 -408
rect 1418 -419 1427 -403
rect 1443 -419 1452 -403
rect 1459 -408 1469 -388
rect 1479 -408 1493 -388
rect 1494 -401 1505 -388
rect 1459 -419 1493 -408
rect 1494 -419 1505 -403
rect 1551 -412 1567 -396
rect 1574 -398 1604 -346
rect 1638 -350 1639 -343
rect 1623 -358 1639 -350
rect 1610 -390 1623 -371
rect 1638 -390 1668 -374
rect 1610 -406 1684 -390
rect 1610 -408 1623 -406
rect 1638 -408 1672 -406
rect 1275 -430 1288 -428
rect 1303 -430 1337 -428
rect 1275 -446 1337 -430
rect 1381 -435 1397 -432
rect 1459 -435 1489 -424
rect 1537 -428 1583 -412
rect 1610 -424 1684 -408
rect 1537 -430 1571 -428
rect 1536 -446 1583 -430
rect 1610 -446 1623 -424
rect 1638 -446 1668 -424
rect 1695 -446 1696 -430
rect 1711 -446 1724 -286
rect 1754 -390 1767 -286
rect 1812 -308 1813 -298
rect 1828 -308 1841 -298
rect 1812 -312 1841 -308
rect 1846 -312 1876 -286
rect 1894 -300 1910 -298
rect 1982 -300 2035 -286
rect 1983 -302 2047 -300
rect 2090 -302 2105 -286
rect 2154 -289 2184 -286
rect 2154 -292 2190 -289
rect 2120 -300 2136 -298
rect 1894 -312 1909 -308
rect 1812 -314 1909 -312
rect 1937 -314 2105 -302
rect 2121 -312 2136 -308
rect 2154 -311 2193 -292
rect 2212 -298 2219 -297
rect 2218 -305 2219 -298
rect 2202 -308 2203 -305
rect 2218 -308 2231 -305
rect 2154 -312 2184 -311
rect 2193 -312 2199 -311
rect 2202 -312 2231 -308
rect 2121 -313 2231 -312
rect 2121 -314 2237 -313
rect 1796 -322 1847 -314
rect 1796 -334 1821 -322
rect 1828 -334 1847 -322
rect 1878 -322 1928 -314
rect 1878 -330 1894 -322
rect 1901 -324 1928 -322
rect 1937 -324 2158 -314
rect 1901 -334 2158 -324
rect 2187 -322 2237 -314
rect 2187 -331 2203 -322
rect 1796 -342 1847 -334
rect 1894 -342 2158 -334
rect 2184 -334 2203 -331
rect 2210 -334 2237 -322
rect 2184 -342 2237 -334
rect 1812 -350 1813 -342
rect 1828 -350 1841 -342
rect 1812 -358 1828 -350
rect 1809 -365 1828 -362
rect 1809 -374 1831 -365
rect 1782 -384 1831 -374
rect 1782 -390 1812 -384
rect 1831 -389 1836 -384
rect 1754 -406 1828 -390
rect 1846 -398 1876 -342
rect 1911 -352 2119 -342
rect 2154 -346 2199 -342
rect 2202 -343 2203 -342
rect 2218 -343 2231 -342
rect 1937 -382 2126 -352
rect 1952 -385 2126 -382
rect 1945 -388 2126 -385
rect 1754 -408 1767 -406
rect 1782 -408 1816 -406
rect 1754 -424 1828 -408
rect 1855 -412 1868 -398
rect 1883 -412 1899 -396
rect 1945 -401 1956 -388
rect 1738 -446 1739 -430
rect 1754 -446 1767 -424
rect 1782 -446 1812 -424
rect 1855 -428 1917 -412
rect 1945 -419 1956 -403
rect 1961 -408 1971 -388
rect 1981 -408 1995 -388
rect 1998 -401 2007 -388
rect 2023 -401 2032 -388
rect 1961 -419 1995 -408
rect 1998 -419 2007 -403
rect 2023 -419 2032 -403
rect 2039 -408 2049 -388
rect 2059 -408 2073 -388
rect 2074 -401 2085 -388
rect 2039 -419 2073 -408
rect 2074 -419 2085 -403
rect 2131 -412 2147 -396
rect 2154 -398 2184 -346
rect 2218 -350 2219 -343
rect 2203 -358 2219 -350
rect 2190 -390 2203 -371
rect 2218 -390 2248 -374
rect 2190 -406 2264 -390
rect 2190 -408 2203 -406
rect 2218 -408 2252 -406
rect 1855 -430 1868 -428
rect 1883 -430 1917 -428
rect 1855 -446 1917 -430
rect 1961 -435 1977 -432
rect 2039 -435 2069 -424
rect 2117 -428 2163 -412
rect 2190 -424 2264 -408
rect 2117 -430 2151 -428
rect 2116 -446 2163 -430
rect 2190 -446 2203 -424
rect 2218 -446 2248 -424
rect 2275 -446 2276 -430
rect 2291 -446 2304 -286
rect 2334 -390 2347 -286
rect 2392 -308 2393 -298
rect 2408 -308 2421 -298
rect 2392 -312 2421 -308
rect 2426 -312 2456 -286
rect 2474 -300 2490 -298
rect 2562 -300 2615 -286
rect 2563 -302 2627 -300
rect 2670 -302 2685 -286
rect 2734 -289 2764 -286
rect 2734 -292 2770 -289
rect 2700 -300 2716 -298
rect 2474 -312 2489 -308
rect 2392 -314 2489 -312
rect 2517 -314 2685 -302
rect 2701 -312 2716 -308
rect 2734 -311 2773 -292
rect 2792 -298 2799 -297
rect 2798 -305 2799 -298
rect 2782 -308 2783 -305
rect 2798 -308 2811 -305
rect 2734 -312 2764 -311
rect 2773 -312 2779 -311
rect 2782 -312 2811 -308
rect 2701 -313 2811 -312
rect 2701 -314 2817 -313
rect 2376 -322 2427 -314
rect 2376 -334 2401 -322
rect 2408 -334 2427 -322
rect 2458 -322 2508 -314
rect 2458 -330 2474 -322
rect 2481 -324 2508 -322
rect 2517 -324 2738 -314
rect 2481 -334 2738 -324
rect 2767 -322 2817 -314
rect 2767 -331 2783 -322
rect 2376 -342 2427 -334
rect 2474 -342 2738 -334
rect 2764 -334 2783 -331
rect 2790 -334 2817 -322
rect 2764 -342 2817 -334
rect 2392 -350 2393 -342
rect 2408 -350 2421 -342
rect 2392 -358 2408 -350
rect 2389 -365 2408 -362
rect 2389 -374 2411 -365
rect 2362 -384 2411 -374
rect 2362 -390 2392 -384
rect 2411 -389 2416 -384
rect 2334 -406 2408 -390
rect 2426 -398 2456 -342
rect 2491 -352 2699 -342
rect 2734 -346 2779 -342
rect 2782 -343 2783 -342
rect 2798 -343 2811 -342
rect 2517 -382 2706 -352
rect 2532 -385 2706 -382
rect 2525 -388 2706 -385
rect 2334 -408 2347 -406
rect 2362 -408 2396 -406
rect 2334 -424 2408 -408
rect 2435 -412 2448 -398
rect 2463 -412 2479 -396
rect 2525 -401 2536 -388
rect 2318 -446 2319 -430
rect 2334 -446 2347 -424
rect 2362 -446 2392 -424
rect 2435 -428 2497 -412
rect 2525 -419 2536 -403
rect 2541 -408 2551 -388
rect 2561 -408 2575 -388
rect 2578 -401 2587 -388
rect 2603 -401 2612 -388
rect 2541 -419 2575 -408
rect 2578 -419 2587 -403
rect 2603 -419 2612 -403
rect 2619 -408 2629 -388
rect 2639 -408 2653 -388
rect 2654 -401 2665 -388
rect 2619 -419 2653 -408
rect 2654 -419 2665 -403
rect 2711 -412 2727 -396
rect 2734 -398 2764 -346
rect 2798 -350 2799 -343
rect 2783 -358 2799 -350
rect 2770 -390 2783 -371
rect 2798 -390 2828 -374
rect 2770 -406 2844 -390
rect 2770 -408 2783 -406
rect 2798 -408 2832 -406
rect 2435 -430 2448 -428
rect 2463 -430 2497 -428
rect 2435 -446 2497 -430
rect 2541 -435 2557 -432
rect 2619 -435 2649 -424
rect 2697 -428 2743 -412
rect 2770 -424 2844 -408
rect 2697 -430 2731 -428
rect 2696 -446 2743 -430
rect 2770 -446 2783 -424
rect 2798 -446 2828 -424
rect 2855 -446 2856 -430
rect 2871 -446 2884 -286
rect 2914 -390 2927 -286
rect 2972 -308 2973 -298
rect 2988 -308 3001 -298
rect 2972 -312 3001 -308
rect 3006 -312 3036 -286
rect 3054 -300 3070 -298
rect 3142 -300 3195 -286
rect 3143 -302 3205 -300
rect 3250 -302 3265 -286
rect 3314 -289 3344 -286
rect 3314 -292 3350 -289
rect 3280 -300 3296 -298
rect 3054 -312 3069 -308
rect 2972 -314 3069 -312
rect 3097 -314 3265 -302
rect 3281 -312 3296 -308
rect 3314 -311 3353 -292
rect 3372 -298 3379 -297
rect 3378 -305 3379 -298
rect 3362 -308 3363 -305
rect 3378 -308 3391 -305
rect 3314 -312 3344 -311
rect 3353 -312 3359 -311
rect 3362 -312 3391 -308
rect 3281 -313 3391 -312
rect 3281 -314 3397 -313
rect 2956 -322 3007 -314
rect 2956 -334 2981 -322
rect 2988 -334 3007 -322
rect 3038 -322 3088 -314
rect 3038 -330 3054 -322
rect 3061 -324 3088 -322
rect 3097 -324 3318 -314
rect 3061 -334 3318 -324
rect 3347 -322 3397 -314
rect 3347 -331 3363 -322
rect 2956 -342 3007 -334
rect 3054 -342 3318 -334
rect 3344 -334 3363 -331
rect 3370 -334 3397 -322
rect 3344 -342 3397 -334
rect 2972 -350 2973 -342
rect 2988 -350 3001 -342
rect 2972 -358 2988 -350
rect 2969 -365 2988 -362
rect 2969 -374 2991 -365
rect 2942 -384 2991 -374
rect 2942 -390 2972 -384
rect 2991 -389 2996 -384
rect 2914 -406 2988 -390
rect 3006 -398 3036 -342
rect 3071 -352 3279 -342
rect 3314 -346 3359 -342
rect 3362 -343 3363 -342
rect 3378 -343 3391 -342
rect 3097 -382 3286 -352
rect 3112 -385 3286 -382
rect 3105 -388 3286 -385
rect 2914 -408 2927 -406
rect 2942 -408 2976 -406
rect 2914 -424 2988 -408
rect 3015 -412 3028 -398
rect 3043 -412 3059 -396
rect 3105 -401 3116 -388
rect 2898 -446 2899 -430
rect 2914 -446 2927 -424
rect 2942 -446 2972 -424
rect 3015 -428 3077 -412
rect 3105 -419 3116 -403
rect 3121 -408 3131 -388
rect 3141 -408 3155 -388
rect 3158 -401 3167 -388
rect 3183 -401 3192 -388
rect 3121 -419 3155 -408
rect 3158 -419 3167 -403
rect 3183 -419 3192 -403
rect 3199 -408 3209 -388
rect 3219 -408 3233 -388
rect 3234 -401 3245 -388
rect 3199 -419 3233 -408
rect 3234 -419 3245 -403
rect 3291 -412 3307 -396
rect 3314 -398 3344 -346
rect 3378 -350 3379 -343
rect 3363 -358 3379 -350
rect 3350 -390 3363 -371
rect 3378 -390 3408 -374
rect 3350 -406 3424 -390
rect 3350 -408 3363 -406
rect 3378 -408 3412 -406
rect 3015 -430 3028 -428
rect 3043 -430 3077 -428
rect 3015 -446 3077 -430
rect 3121 -435 3137 -432
rect 3199 -435 3229 -424
rect 3277 -428 3323 -412
rect 3350 -424 3424 -408
rect 3277 -430 3311 -428
rect 3276 -446 3323 -430
rect 3350 -446 3363 -424
rect 3378 -446 3408 -424
rect 3435 -446 3436 -430
rect 3451 -446 3464 -286
rect 3494 -390 3507 -286
rect 3552 -308 3553 -298
rect 3568 -308 3581 -298
rect 3552 -312 3581 -308
rect 3586 -312 3616 -286
rect 3634 -300 3650 -298
rect 3722 -300 3775 -286
rect 3723 -302 3787 -300
rect 3830 -302 3845 -286
rect 3894 -289 3924 -286
rect 3894 -292 3930 -289
rect 3860 -300 3876 -298
rect 3634 -312 3649 -308
rect 3552 -314 3649 -312
rect 3677 -314 3845 -302
rect 3861 -312 3876 -308
rect 3894 -311 3933 -292
rect 3952 -298 3959 -297
rect 3958 -305 3959 -298
rect 3942 -308 3943 -305
rect 3958 -308 3971 -305
rect 3894 -312 3924 -311
rect 3933 -312 3939 -311
rect 3942 -312 3971 -308
rect 3861 -313 3971 -312
rect 3861 -314 3977 -313
rect 3536 -322 3587 -314
rect 3536 -334 3561 -322
rect 3568 -334 3587 -322
rect 3618 -322 3668 -314
rect 3618 -330 3634 -322
rect 3641 -324 3668 -322
rect 3677 -324 3898 -314
rect 3641 -334 3898 -324
rect 3927 -322 3977 -314
rect 3927 -331 3943 -322
rect 3536 -342 3587 -334
rect 3634 -342 3898 -334
rect 3924 -334 3943 -331
rect 3950 -334 3977 -322
rect 3924 -342 3977 -334
rect 3552 -350 3553 -342
rect 3568 -350 3581 -342
rect 3552 -358 3568 -350
rect 3549 -365 3568 -362
rect 3549 -374 3571 -365
rect 3522 -384 3571 -374
rect 3522 -390 3552 -384
rect 3571 -389 3576 -384
rect 3494 -406 3568 -390
rect 3586 -398 3616 -342
rect 3651 -352 3859 -342
rect 3894 -346 3939 -342
rect 3942 -343 3943 -342
rect 3958 -343 3971 -342
rect 3677 -382 3866 -352
rect 3692 -385 3866 -382
rect 3685 -388 3866 -385
rect 3494 -408 3507 -406
rect 3522 -408 3556 -406
rect 3494 -424 3568 -408
rect 3595 -412 3608 -398
rect 3623 -412 3639 -396
rect 3685 -401 3696 -388
rect 3478 -446 3479 -430
rect 3494 -446 3507 -424
rect 3522 -446 3552 -424
rect 3595 -428 3657 -412
rect 3685 -419 3696 -403
rect 3701 -408 3711 -388
rect 3721 -408 3735 -388
rect 3738 -401 3747 -388
rect 3763 -401 3772 -388
rect 3701 -419 3735 -408
rect 3738 -419 3747 -403
rect 3763 -419 3772 -403
rect 3779 -408 3789 -388
rect 3799 -408 3813 -388
rect 3814 -401 3825 -388
rect 3779 -419 3813 -408
rect 3814 -419 3825 -403
rect 3871 -412 3887 -396
rect 3894 -398 3924 -346
rect 3958 -350 3959 -343
rect 3943 -358 3959 -350
rect 3930 -390 3943 -371
rect 3958 -390 3988 -374
rect 3930 -406 4004 -390
rect 3930 -408 3943 -406
rect 3958 -408 3992 -406
rect 3595 -430 3608 -428
rect 3623 -430 3657 -428
rect 3595 -446 3657 -430
rect 3701 -435 3717 -432
rect 3779 -435 3809 -424
rect 3857 -428 3903 -412
rect 3930 -424 4004 -408
rect 3857 -430 3891 -428
rect 3856 -446 3903 -430
rect 3930 -446 3943 -424
rect 3958 -446 3988 -424
rect 4015 -446 4016 -430
rect 4031 -446 4044 -286
rect 4074 -390 4087 -286
rect 4132 -308 4133 -298
rect 4148 -308 4161 -298
rect 4132 -312 4161 -308
rect 4166 -312 4196 -286
rect 4214 -300 4230 -298
rect 4302 -300 4355 -286
rect 4303 -302 4367 -300
rect 4410 -302 4425 -286
rect 4474 -289 4504 -286
rect 4611 -287 6944 -286
rect 4474 -292 4510 -289
rect 4440 -300 4456 -298
rect 4214 -312 4229 -308
rect 4132 -314 4229 -312
rect 4257 -314 4425 -302
rect 4441 -312 4456 -308
rect 4474 -311 4513 -292
rect 4532 -298 4539 -297
rect 4538 -305 4539 -298
rect 4522 -308 4523 -305
rect 4538 -308 4551 -305
rect 4474 -312 4504 -311
rect 4513 -312 4519 -311
rect 4522 -312 4551 -308
rect 4441 -313 4551 -312
rect 4441 -314 4557 -313
rect 4116 -322 4167 -314
rect 4116 -334 4141 -322
rect 4148 -334 4167 -322
rect 4198 -322 4248 -314
rect 4198 -330 4214 -322
rect 4221 -324 4248 -322
rect 4257 -324 4478 -314
rect 4221 -334 4478 -324
rect 4507 -322 4557 -314
rect 4507 -331 4523 -322
rect 4116 -342 4167 -334
rect 4214 -342 4478 -334
rect 4504 -334 4523 -331
rect 4530 -334 4557 -322
rect 4504 -342 4557 -334
rect 4132 -350 4133 -342
rect 4148 -350 4161 -342
rect 4132 -358 4148 -350
rect 4129 -365 4148 -362
rect 4129 -374 4151 -365
rect 4102 -384 4151 -374
rect 4102 -390 4132 -384
rect 4151 -389 4156 -384
rect 4074 -406 4148 -390
rect 4166 -398 4196 -342
rect 4231 -352 4439 -342
rect 4474 -346 4519 -342
rect 4522 -343 4523 -342
rect 4538 -343 4551 -342
rect 4257 -382 4446 -352
rect 4272 -385 4446 -382
rect 4265 -388 4446 -385
rect 4074 -408 4087 -406
rect 4102 -408 4136 -406
rect 4074 -424 4148 -408
rect 4175 -412 4188 -398
rect 4203 -412 4219 -396
rect 4265 -401 4276 -388
rect 4058 -446 4059 -430
rect 4074 -446 4087 -424
rect 4102 -446 4132 -424
rect 4175 -428 4237 -412
rect 4265 -419 4276 -403
rect 4281 -408 4291 -388
rect 4301 -408 4315 -388
rect 4318 -401 4327 -388
rect 4343 -401 4352 -388
rect 4281 -419 4315 -408
rect 4318 -419 4327 -403
rect 4343 -419 4352 -403
rect 4359 -408 4369 -388
rect 4379 -408 4393 -388
rect 4394 -401 4405 -388
rect 4359 -419 4393 -408
rect 4394 -419 4405 -403
rect 4451 -412 4467 -396
rect 4474 -398 4504 -346
rect 4538 -350 4539 -343
rect 4523 -358 4539 -350
rect 4510 -390 4523 -371
rect 4538 -390 4568 -374
rect 4510 -406 4584 -390
rect 4510 -408 4523 -406
rect 4538 -408 4572 -406
rect 4175 -430 4188 -428
rect 4203 -430 4237 -428
rect 4175 -446 4237 -430
rect 4281 -435 4297 -432
rect 4359 -435 4389 -424
rect 4437 -428 4483 -412
rect 4510 -424 4584 -408
rect 4437 -430 4471 -428
rect 4436 -446 4483 -430
rect 4510 -446 4523 -424
rect 4538 -446 4568 -424
rect 4595 -446 4596 -430
rect 4611 -446 4624 -287
rect 4654 -391 4667 -287
rect 4712 -309 4713 -299
rect 4733 -301 4741 -299
rect 4731 -303 4741 -301
rect 4728 -309 4741 -303
rect 4712 -313 4741 -309
rect 4746 -313 4776 -287
rect 4794 -301 4810 -299
rect 4882 -301 4933 -287
rect 4883 -303 4947 -301
rect 4990 -303 5005 -287
rect 5054 -290 5084 -287
rect 5054 -293 5090 -290
rect 5020 -301 5036 -299
rect 4794 -313 4809 -309
rect 4712 -315 4809 -313
rect 4837 -315 5005 -303
rect 5021 -313 5036 -309
rect 5054 -312 5093 -293
rect 5112 -299 5119 -298
rect 5118 -306 5119 -299
rect 5102 -309 5103 -306
rect 5118 -309 5131 -306
rect 5054 -313 5084 -312
rect 5093 -313 5099 -312
rect 5102 -313 5131 -309
rect 5021 -314 5131 -313
rect 5021 -315 5137 -314
rect 4696 -323 4747 -315
rect 4696 -335 4721 -323
rect 4728 -335 4747 -323
rect 4778 -323 4828 -315
rect 4778 -331 4794 -323
rect 4801 -325 4828 -323
rect 4837 -325 5058 -315
rect 4801 -335 5058 -325
rect 5087 -323 5137 -315
rect 5087 -332 5103 -323
rect 4696 -343 4747 -335
rect 4794 -343 5058 -335
rect 5084 -335 5103 -332
rect 5110 -335 5137 -323
rect 5084 -343 5137 -335
rect 4712 -351 4713 -343
rect 4728 -351 4741 -343
rect 4712 -359 4728 -351
rect 4709 -366 4728 -363
rect 4709 -375 4731 -366
rect 4682 -385 4731 -375
rect 4682 -391 4712 -385
rect 4731 -390 4736 -385
rect 4654 -407 4728 -391
rect 4746 -399 4776 -343
rect 4811 -353 5019 -343
rect 5054 -347 5099 -343
rect 5102 -344 5103 -343
rect 5118 -344 5131 -343
rect 4837 -383 5026 -353
rect 4852 -386 5026 -383
rect 4845 -389 5026 -386
rect 4654 -409 4667 -407
rect 4682 -409 4716 -407
rect 4654 -425 4728 -409
rect 4755 -413 4768 -399
rect 4783 -413 4799 -397
rect 4845 -402 4856 -389
rect -8 -454 33 -446
rect -8 -480 7 -454
rect 14 -480 33 -454
rect 97 -458 159 -446
rect 171 -458 246 -446
rect 304 -458 379 -446
rect 391 -458 422 -446
rect 428 -458 463 -446
rect 97 -460 259 -458
rect -8 -488 33 -480
rect 115 -484 128 -460
rect 143 -462 158 -460
rect -2 -498 -1 -488
rect 14 -498 27 -488
rect 42 -498 72 -484
rect 115 -498 158 -484
rect 182 -487 189 -480
rect 192 -484 259 -460
rect 291 -460 463 -458
rect 261 -482 289 -478
rect 291 -482 371 -460
rect 392 -462 407 -460
rect 261 -484 371 -482
rect 192 -488 371 -484
rect 165 -498 195 -488
rect 197 -498 350 -488
rect 358 -498 388 -488
rect 392 -498 422 -484
rect 450 -498 463 -460
rect 535 -454 570 -446
rect 535 -480 536 -454
rect 543 -480 570 -454
rect 478 -498 508 -484
rect 535 -488 570 -480
rect 572 -454 613 -446
rect 572 -480 587 -454
rect 594 -480 613 -454
rect 677 -458 739 -446
rect 751 -458 826 -446
rect 884 -458 959 -446
rect 971 -458 1002 -446
rect 1008 -458 1043 -446
rect 677 -460 839 -458
rect 572 -488 613 -480
rect 695 -484 708 -460
rect 723 -462 738 -460
rect 535 -498 536 -488
rect 551 -498 564 -488
rect 578 -498 579 -488
rect 594 -498 607 -488
rect 622 -498 652 -484
rect 695 -498 738 -484
rect 762 -487 769 -480
rect 772 -484 839 -460
rect 871 -460 1043 -458
rect 841 -482 869 -478
rect 871 -482 951 -460
rect 972 -462 987 -460
rect 841 -484 951 -482
rect 772 -488 951 -484
rect 745 -498 775 -488
rect 777 -498 930 -488
rect 938 -498 968 -488
rect 972 -498 1002 -484
rect 1030 -498 1043 -460
rect 1115 -454 1150 -446
rect 1115 -480 1116 -454
rect 1123 -480 1150 -454
rect 1058 -498 1088 -484
rect 1115 -488 1150 -480
rect 1152 -454 1193 -446
rect 1152 -480 1167 -454
rect 1174 -480 1193 -454
rect 1257 -458 1319 -446
rect 1331 -458 1406 -446
rect 1464 -458 1539 -446
rect 1551 -458 1582 -446
rect 1588 -458 1623 -446
rect 1257 -460 1419 -458
rect 1152 -488 1193 -480
rect 1275 -484 1288 -460
rect 1303 -462 1318 -460
rect 1115 -498 1116 -488
rect 1131 -498 1144 -488
rect 1158 -498 1159 -488
rect 1174 -498 1187 -488
rect 1202 -498 1232 -484
rect 1275 -498 1318 -484
rect 1342 -487 1349 -480
rect 1352 -484 1419 -460
rect 1451 -460 1623 -458
rect 1421 -482 1449 -478
rect 1451 -482 1531 -460
rect 1552 -462 1567 -460
rect 1421 -484 1531 -482
rect 1352 -488 1531 -484
rect 1325 -498 1355 -488
rect 1357 -498 1510 -488
rect 1518 -498 1548 -488
rect 1552 -498 1582 -484
rect 1610 -498 1623 -460
rect 1695 -454 1730 -446
rect 1695 -480 1696 -454
rect 1703 -480 1730 -454
rect 1638 -498 1668 -484
rect 1695 -488 1730 -480
rect 1732 -454 1773 -446
rect 1732 -480 1747 -454
rect 1754 -480 1773 -454
rect 1837 -458 1899 -446
rect 1911 -458 1986 -446
rect 2044 -458 2119 -446
rect 2131 -458 2162 -446
rect 2168 -458 2203 -446
rect 1837 -460 1999 -458
rect 1732 -488 1773 -480
rect 1855 -484 1868 -460
rect 1883 -462 1898 -460
rect 1695 -498 1696 -488
rect 1711 -498 1724 -488
rect 1738 -498 1739 -488
rect 1754 -498 1767 -488
rect 1782 -498 1812 -484
rect 1855 -498 1898 -484
rect 1922 -487 1929 -480
rect 1932 -484 1999 -460
rect 2031 -460 2203 -458
rect 2001 -482 2029 -478
rect 2031 -482 2111 -460
rect 2132 -462 2147 -460
rect 2001 -484 2111 -482
rect 1932 -488 2111 -484
rect 1905 -498 1935 -488
rect 1937 -498 2090 -488
rect 2098 -498 2128 -488
rect 2132 -498 2162 -484
rect 2190 -498 2203 -460
rect 2275 -454 2310 -446
rect 2275 -480 2276 -454
rect 2283 -480 2310 -454
rect 2218 -498 2248 -484
rect 2275 -488 2310 -480
rect 2312 -454 2353 -446
rect 2312 -480 2327 -454
rect 2334 -480 2353 -454
rect 2417 -458 2479 -446
rect 2491 -458 2566 -446
rect 2624 -458 2699 -446
rect 2711 -458 2742 -446
rect 2748 -458 2783 -446
rect 2417 -460 2579 -458
rect 2312 -488 2353 -480
rect 2435 -484 2448 -460
rect 2463 -462 2478 -460
rect 2275 -498 2276 -488
rect 2291 -498 2304 -488
rect 2318 -498 2319 -488
rect 2334 -498 2347 -488
rect 2362 -498 2392 -484
rect 2435 -498 2478 -484
rect 2502 -487 2509 -480
rect 2512 -484 2579 -460
rect 2611 -460 2783 -458
rect 2581 -482 2609 -478
rect 2611 -482 2691 -460
rect 2712 -462 2727 -460
rect 2581 -484 2691 -482
rect 2512 -488 2691 -484
rect 2485 -498 2515 -488
rect 2517 -498 2670 -488
rect 2678 -498 2708 -488
rect 2712 -498 2742 -484
rect 2770 -498 2783 -460
rect 2855 -454 2890 -446
rect 2855 -480 2856 -454
rect 2863 -480 2890 -454
rect 2798 -498 2828 -484
rect 2855 -488 2890 -480
rect 2892 -454 2933 -446
rect 2892 -480 2907 -454
rect 2914 -480 2933 -454
rect 2997 -458 3059 -446
rect 3071 -458 3146 -446
rect 3204 -458 3279 -446
rect 3291 -458 3322 -446
rect 3328 -458 3363 -446
rect 2997 -460 3159 -458
rect 2892 -488 2933 -480
rect 3015 -484 3028 -460
rect 3043 -462 3058 -460
rect 2855 -498 2856 -488
rect 2871 -498 2884 -488
rect 2898 -498 2899 -488
rect 2914 -498 2927 -488
rect 2942 -498 2972 -484
rect 3015 -498 3058 -484
rect 3082 -487 3089 -480
rect 3092 -484 3159 -460
rect 3191 -460 3363 -458
rect 3161 -482 3189 -478
rect 3191 -482 3271 -460
rect 3292 -462 3307 -460
rect 3161 -484 3271 -482
rect 3092 -488 3271 -484
rect 3065 -498 3095 -488
rect 3097 -498 3250 -488
rect 3258 -498 3288 -488
rect 3292 -498 3322 -484
rect 3350 -498 3363 -460
rect 3435 -454 3470 -446
rect 3435 -480 3436 -454
rect 3443 -480 3470 -454
rect 3378 -498 3408 -484
rect 3435 -488 3470 -480
rect 3472 -454 3513 -446
rect 3472 -480 3487 -454
rect 3494 -480 3513 -454
rect 3577 -458 3639 -446
rect 3651 -458 3726 -446
rect 3784 -458 3859 -446
rect 3871 -458 3902 -446
rect 3908 -458 3943 -446
rect 3577 -460 3739 -458
rect 3472 -488 3513 -480
rect 3595 -484 3608 -460
rect 3623 -462 3638 -460
rect 3435 -498 3436 -488
rect 3451 -498 3464 -488
rect 3478 -498 3479 -488
rect 3494 -498 3507 -488
rect 3522 -498 3552 -484
rect 3595 -498 3638 -484
rect 3662 -487 3669 -480
rect 3672 -484 3739 -460
rect 3771 -460 3943 -458
rect 3741 -482 3769 -478
rect 3771 -482 3851 -460
rect 3872 -462 3887 -460
rect 3741 -484 3851 -482
rect 3672 -488 3851 -484
rect 3645 -498 3675 -488
rect 3677 -498 3830 -488
rect 3838 -498 3868 -488
rect 3872 -498 3902 -484
rect 3930 -498 3943 -460
rect 4015 -454 4050 -446
rect 4015 -480 4016 -454
rect 4023 -480 4050 -454
rect 3958 -498 3988 -484
rect 4015 -488 4050 -480
rect 4052 -454 4093 -446
rect 4052 -480 4067 -454
rect 4074 -480 4093 -454
rect 4157 -458 4219 -446
rect 4231 -458 4306 -446
rect 4364 -458 4439 -446
rect 4451 -458 4482 -446
rect 4488 -458 4523 -446
rect 4157 -460 4319 -458
rect 4052 -488 4093 -480
rect 4175 -484 4188 -460
rect 4203 -462 4218 -460
rect 4015 -498 4016 -488
rect 4031 -498 4044 -488
rect 4058 -498 4059 -488
rect 4074 -498 4087 -488
rect 4102 -498 4132 -484
rect 4175 -498 4218 -484
rect 4242 -487 4249 -480
rect 4252 -484 4319 -460
rect 4351 -460 4523 -458
rect 4321 -482 4349 -478
rect 4351 -482 4431 -460
rect 4452 -462 4467 -460
rect 4321 -484 4431 -482
rect 4252 -488 4431 -484
rect 4225 -498 4255 -488
rect 4257 -498 4410 -488
rect 4418 -498 4448 -488
rect 4452 -498 4482 -484
rect 4510 -498 4523 -460
rect 4595 -454 4630 -446
rect 4638 -447 4639 -431
rect 4654 -447 4667 -425
rect 4682 -447 4712 -425
rect 4755 -429 4817 -413
rect 4845 -420 4856 -404
rect 4861 -409 4871 -389
rect 4881 -409 4895 -389
rect 4898 -402 4907 -389
rect 4923 -402 4932 -389
rect 4861 -420 4895 -409
rect 4898 -420 4907 -404
rect 4923 -420 4932 -404
rect 4939 -409 4949 -389
rect 4959 -409 4973 -389
rect 4974 -402 4985 -389
rect 4939 -420 4973 -409
rect 4974 -420 4985 -404
rect 5031 -413 5047 -397
rect 5054 -399 5084 -347
rect 5118 -351 5119 -344
rect 5103 -359 5119 -351
rect 5090 -391 5103 -372
rect 5118 -391 5148 -375
rect 5090 -407 5164 -391
rect 5090 -409 5103 -407
rect 5118 -409 5152 -407
rect 4755 -431 4768 -429
rect 4783 -431 4817 -429
rect 4755 -447 4817 -431
rect 4861 -436 4877 -433
rect 4939 -436 4969 -425
rect 5017 -429 5063 -413
rect 5090 -425 5164 -409
rect 5017 -431 5051 -429
rect 5016 -447 5063 -431
rect 5090 -447 5103 -425
rect 5118 -447 5148 -425
rect 5175 -447 5176 -431
rect 5191 -447 5204 -287
rect 5234 -391 5247 -287
rect 5292 -309 5293 -299
rect 5313 -301 5321 -299
rect 5311 -303 5321 -301
rect 5308 -309 5321 -303
rect 5292 -313 5321 -309
rect 5326 -313 5356 -287
rect 5374 -301 5390 -299
rect 5462 -301 5513 -287
rect 5463 -303 5527 -301
rect 5570 -303 5585 -287
rect 5634 -290 5664 -287
rect 5634 -293 5670 -290
rect 5600 -301 5616 -299
rect 5374 -313 5389 -309
rect 5292 -315 5389 -313
rect 5417 -315 5585 -303
rect 5601 -313 5616 -309
rect 5634 -312 5673 -293
rect 5692 -299 5699 -298
rect 5698 -306 5699 -299
rect 5682 -309 5683 -306
rect 5698 -309 5711 -306
rect 5634 -313 5664 -312
rect 5673 -313 5679 -312
rect 5682 -313 5711 -309
rect 5601 -314 5711 -313
rect 5601 -315 5717 -314
rect 5276 -323 5327 -315
rect 5276 -335 5301 -323
rect 5308 -335 5327 -323
rect 5358 -323 5408 -315
rect 5358 -331 5374 -323
rect 5381 -325 5408 -323
rect 5417 -325 5638 -315
rect 5381 -335 5638 -325
rect 5667 -323 5717 -315
rect 5667 -332 5683 -323
rect 5276 -343 5327 -335
rect 5374 -343 5638 -335
rect 5664 -335 5683 -332
rect 5690 -335 5717 -323
rect 5664 -343 5717 -335
rect 5292 -351 5293 -343
rect 5308 -351 5321 -343
rect 5292 -359 5308 -351
rect 5289 -366 5308 -363
rect 5289 -375 5311 -366
rect 5262 -385 5311 -375
rect 5262 -391 5292 -385
rect 5311 -390 5316 -385
rect 5234 -407 5308 -391
rect 5326 -399 5356 -343
rect 5391 -353 5599 -343
rect 5634 -347 5679 -343
rect 5682 -344 5683 -343
rect 5698 -344 5711 -343
rect 5417 -383 5606 -353
rect 5432 -386 5606 -383
rect 5425 -389 5606 -386
rect 5234 -409 5247 -407
rect 5262 -409 5296 -407
rect 5234 -425 5308 -409
rect 5335 -413 5348 -399
rect 5363 -413 5379 -397
rect 5425 -402 5436 -389
rect 5218 -447 5219 -431
rect 5234 -447 5247 -425
rect 5262 -447 5292 -425
rect 5335 -429 5397 -413
rect 5425 -420 5436 -404
rect 5441 -409 5451 -389
rect 5461 -409 5475 -389
rect 5478 -402 5487 -389
rect 5503 -402 5512 -389
rect 5441 -420 5475 -409
rect 5478 -420 5487 -404
rect 5503 -420 5512 -404
rect 5519 -409 5529 -389
rect 5539 -409 5553 -389
rect 5554 -402 5565 -389
rect 5519 -420 5553 -409
rect 5554 -420 5565 -404
rect 5611 -413 5627 -397
rect 5634 -399 5664 -347
rect 5698 -351 5699 -344
rect 5683 -359 5699 -351
rect 5670 -391 5683 -372
rect 5698 -391 5728 -375
rect 5670 -407 5744 -391
rect 5670 -409 5683 -407
rect 5698 -409 5732 -407
rect 5335 -431 5348 -429
rect 5363 -431 5397 -429
rect 5335 -447 5397 -431
rect 5441 -436 5457 -433
rect 5519 -436 5549 -425
rect 5597 -429 5643 -413
rect 5670 -425 5744 -409
rect 5597 -431 5631 -429
rect 5596 -447 5643 -431
rect 5670 -447 5683 -425
rect 5698 -447 5728 -425
rect 5755 -447 5756 -431
rect 5771 -447 5784 -287
rect 5814 -391 5827 -287
rect 5872 -309 5873 -299
rect 5893 -301 5901 -299
rect 5891 -303 5901 -301
rect 5888 -309 5901 -303
rect 5872 -313 5901 -309
rect 5906 -313 5936 -287
rect 5954 -301 5970 -299
rect 6042 -301 6093 -287
rect 6043 -303 6107 -301
rect 6150 -303 6165 -287
rect 6214 -290 6244 -287
rect 6214 -293 6250 -290
rect 6180 -301 6196 -299
rect 5954 -313 5969 -309
rect 5872 -315 5969 -313
rect 5997 -315 6165 -303
rect 6181 -313 6196 -309
rect 6214 -312 6253 -293
rect 6272 -299 6279 -298
rect 6278 -306 6279 -299
rect 6262 -309 6263 -306
rect 6278 -309 6291 -306
rect 6214 -313 6244 -312
rect 6253 -313 6259 -312
rect 6262 -313 6291 -309
rect 6181 -314 6291 -313
rect 6181 -315 6297 -314
rect 5856 -323 5907 -315
rect 5856 -335 5881 -323
rect 5888 -335 5907 -323
rect 5938 -323 5988 -315
rect 5938 -331 5954 -323
rect 5961 -325 5988 -323
rect 5997 -325 6218 -315
rect 5961 -335 6218 -325
rect 6247 -323 6297 -315
rect 6247 -332 6263 -323
rect 5856 -343 5907 -335
rect 5954 -343 6218 -335
rect 6244 -335 6263 -332
rect 6270 -335 6297 -323
rect 6244 -343 6297 -335
rect 5872 -351 5873 -343
rect 5888 -351 5901 -343
rect 5872 -359 5888 -351
rect 5869 -366 5888 -363
rect 5869 -375 5891 -366
rect 5842 -385 5891 -375
rect 5842 -391 5872 -385
rect 5891 -390 5896 -385
rect 5814 -407 5888 -391
rect 5906 -399 5936 -343
rect 5971 -353 6179 -343
rect 6214 -347 6259 -343
rect 6262 -344 6263 -343
rect 6278 -344 6291 -343
rect 5997 -383 6186 -353
rect 6012 -386 6186 -383
rect 6005 -389 6186 -386
rect 5814 -409 5827 -407
rect 5842 -409 5876 -407
rect 5814 -425 5888 -409
rect 5915 -413 5928 -399
rect 5943 -413 5959 -397
rect 6005 -402 6016 -389
rect 5798 -447 5799 -431
rect 5814 -447 5827 -425
rect 5842 -447 5872 -425
rect 5915 -429 5977 -413
rect 6005 -420 6016 -404
rect 6021 -409 6031 -389
rect 6041 -409 6055 -389
rect 6058 -402 6067 -389
rect 6083 -402 6092 -389
rect 6021 -420 6055 -409
rect 6058 -420 6067 -404
rect 6083 -420 6092 -404
rect 6099 -409 6109 -389
rect 6119 -409 6133 -389
rect 6134 -402 6145 -389
rect 6099 -420 6133 -409
rect 6134 -420 6145 -404
rect 6191 -413 6207 -397
rect 6214 -399 6244 -347
rect 6278 -351 6279 -344
rect 6263 -359 6279 -351
rect 6250 -391 6263 -372
rect 6278 -391 6308 -375
rect 6250 -407 6324 -391
rect 6250 -409 6263 -407
rect 6278 -409 6312 -407
rect 5915 -431 5928 -429
rect 5943 -431 5977 -429
rect 5915 -447 5977 -431
rect 6021 -436 6037 -433
rect 6099 -436 6129 -425
rect 6177 -429 6223 -413
rect 6250 -425 6324 -409
rect 6177 -431 6211 -429
rect 6176 -447 6223 -431
rect 6250 -447 6263 -425
rect 6278 -447 6308 -425
rect 6335 -447 6336 -431
rect 6351 -447 6364 -287
rect 6394 -391 6407 -287
rect 6452 -309 6453 -299
rect 6473 -301 6481 -299
rect 6471 -303 6481 -301
rect 6468 -309 6481 -303
rect 6452 -313 6481 -309
rect 6486 -313 6516 -287
rect 6534 -301 6550 -299
rect 6622 -301 6673 -287
rect 6623 -303 6687 -301
rect 6730 -303 6745 -287
rect 6794 -290 6824 -287
rect 6794 -293 6830 -290
rect 6760 -301 6776 -299
rect 6534 -313 6549 -309
rect 6452 -315 6549 -313
rect 6577 -315 6745 -303
rect 6761 -313 6776 -309
rect 6794 -312 6833 -293
rect 6852 -299 6859 -298
rect 6858 -306 6859 -299
rect 6842 -309 6843 -306
rect 6858 -309 6871 -306
rect 6794 -313 6824 -312
rect 6833 -313 6839 -312
rect 6842 -313 6871 -309
rect 6761 -314 6871 -313
rect 6761 -315 6877 -314
rect 6436 -323 6487 -315
rect 6436 -335 6461 -323
rect 6468 -335 6487 -323
rect 6518 -323 6568 -315
rect 6518 -331 6534 -323
rect 6541 -325 6568 -323
rect 6577 -325 6798 -315
rect 6541 -335 6798 -325
rect 6827 -323 6877 -315
rect 6827 -332 6843 -323
rect 6436 -343 6487 -335
rect 6534 -343 6798 -335
rect 6824 -335 6843 -332
rect 6850 -335 6877 -323
rect 6824 -343 6877 -335
rect 6452 -351 6453 -343
rect 6468 -351 6481 -343
rect 6452 -359 6468 -351
rect 6449 -366 6468 -363
rect 6449 -375 6471 -366
rect 6422 -385 6471 -375
rect 6422 -391 6452 -385
rect 6471 -390 6476 -385
rect 6394 -407 6468 -391
rect 6486 -399 6516 -343
rect 6551 -353 6759 -343
rect 6794 -347 6839 -343
rect 6842 -344 6843 -343
rect 6858 -344 6871 -343
rect 6577 -383 6766 -353
rect 6592 -386 6766 -383
rect 6585 -389 6766 -386
rect 6394 -409 6407 -407
rect 6422 -409 6456 -407
rect 6394 -425 6468 -409
rect 6495 -413 6508 -399
rect 6523 -413 6539 -397
rect 6585 -402 6596 -389
rect 6378 -447 6379 -431
rect 6394 -447 6407 -425
rect 6422 -447 6452 -425
rect 6495 -429 6557 -413
rect 6585 -420 6596 -404
rect 6601 -409 6611 -389
rect 6621 -409 6635 -389
rect 6638 -402 6647 -389
rect 6663 -402 6672 -389
rect 6601 -420 6635 -409
rect 6638 -420 6647 -404
rect 6663 -420 6672 -404
rect 6679 -409 6689 -389
rect 6699 -409 6713 -389
rect 6714 -402 6725 -389
rect 6679 -420 6713 -409
rect 6714 -420 6725 -404
rect 6771 -413 6787 -397
rect 6794 -399 6824 -347
rect 6858 -351 6859 -344
rect 6843 -359 6859 -351
rect 6830 -391 6843 -372
rect 6858 -391 6888 -375
rect 6830 -407 6904 -391
rect 6830 -409 6843 -407
rect 6858 -409 6892 -407
rect 6495 -431 6508 -429
rect 6523 -431 6557 -429
rect 6495 -447 6557 -431
rect 6601 -436 6617 -433
rect 6679 -436 6709 -425
rect 6757 -429 6803 -413
rect 6830 -425 6904 -409
rect 6757 -431 6791 -429
rect 6756 -447 6803 -431
rect 6830 -447 6843 -425
rect 6858 -447 6888 -425
rect 6915 -447 6916 -431
rect 6931 -447 6944 -287
rect 4595 -480 4596 -454
rect 4603 -480 4630 -454
rect 4538 -498 4568 -484
rect 4595 -488 4630 -480
rect 4632 -455 4673 -447
rect 4632 -481 4647 -455
rect 4654 -481 4673 -455
rect 4737 -459 4799 -447
rect 4811 -459 4886 -447
rect 4944 -459 5019 -447
rect 5031 -459 5062 -447
rect 5068 -459 5103 -447
rect 4737 -461 4899 -459
rect 4755 -479 4768 -461
rect 4783 -463 4798 -461
rect 4595 -498 4596 -488
rect 4611 -498 4624 -488
rect 4632 -489 4673 -481
rect 4756 -485 4768 -479
rect 4832 -479 4899 -461
rect 4931 -461 5103 -459
rect 4931 -479 5011 -461
rect 5032 -463 5047 -461
rect -2 -499 4624 -498
rect 4638 -499 4639 -489
rect 4654 -499 4667 -489
rect 4682 -499 4712 -485
rect 4756 -499 4798 -485
rect 4822 -488 4829 -481
rect 4832 -489 5011 -479
rect 4805 -499 4835 -489
rect 4837 -499 4990 -489
rect 4998 -499 5028 -489
rect 5032 -499 5062 -485
rect 5090 -499 5103 -461
rect 5175 -455 5210 -447
rect 5175 -481 5176 -455
rect 5183 -481 5210 -455
rect 5118 -499 5148 -485
rect 5175 -489 5210 -481
rect 5212 -455 5253 -447
rect 5212 -481 5227 -455
rect 5234 -481 5253 -455
rect 5317 -459 5379 -447
rect 5391 -459 5466 -447
rect 5524 -459 5599 -447
rect 5611 -459 5642 -447
rect 5648 -459 5683 -447
rect 5317 -461 5479 -459
rect 5335 -479 5348 -461
rect 5363 -463 5378 -461
rect 5212 -489 5253 -481
rect 5336 -485 5348 -479
rect 5412 -479 5479 -461
rect 5511 -461 5683 -459
rect 5511 -479 5591 -461
rect 5612 -463 5627 -461
rect 5175 -499 5176 -489
rect 5191 -499 5204 -489
rect 5218 -499 5219 -489
rect 5234 -499 5247 -489
rect 5262 -499 5292 -485
rect 5336 -499 5378 -485
rect 5402 -488 5409 -481
rect 5412 -489 5591 -479
rect 5385 -499 5415 -489
rect 5417 -499 5570 -489
rect 5578 -499 5608 -489
rect 5612 -499 5642 -485
rect 5670 -499 5683 -461
rect 5755 -455 5790 -447
rect 5755 -481 5756 -455
rect 5763 -481 5790 -455
rect 5698 -499 5728 -485
rect 5755 -489 5790 -481
rect 5792 -455 5833 -447
rect 5792 -481 5807 -455
rect 5814 -481 5833 -455
rect 5897 -459 5959 -447
rect 5971 -459 6046 -447
rect 6104 -459 6179 -447
rect 6191 -459 6222 -447
rect 6228 -459 6263 -447
rect 5897 -461 6059 -459
rect 5915 -479 5928 -461
rect 5943 -463 5958 -461
rect 5792 -489 5833 -481
rect 5916 -485 5928 -479
rect 5992 -479 6059 -461
rect 6091 -461 6263 -459
rect 6091 -479 6171 -461
rect 6192 -463 6207 -461
rect 5755 -499 5756 -489
rect 5771 -499 5784 -489
rect 5798 -499 5799 -489
rect 5814 -499 5827 -489
rect 5842 -499 5872 -485
rect 5916 -499 5958 -485
rect 5982 -488 5989 -481
rect 5992 -489 6171 -479
rect 5965 -499 5995 -489
rect 5997 -499 6150 -489
rect 6158 -499 6188 -489
rect 6192 -499 6222 -485
rect 6250 -499 6263 -461
rect 6335 -455 6370 -447
rect 6335 -481 6336 -455
rect 6343 -481 6370 -455
rect 6278 -499 6308 -485
rect 6335 -489 6370 -481
rect 6372 -455 6413 -447
rect 6372 -481 6387 -455
rect 6394 -481 6413 -455
rect 6477 -459 6539 -447
rect 6551 -459 6626 -447
rect 6684 -459 6759 -447
rect 6771 -459 6802 -447
rect 6808 -459 6843 -447
rect 6477 -461 6639 -459
rect 6495 -479 6508 -461
rect 6523 -463 6538 -461
rect 6372 -489 6413 -481
rect 6496 -485 6508 -479
rect 6572 -479 6639 -461
rect 6671 -461 6843 -459
rect 6671 -479 6751 -461
rect 6772 -463 6787 -461
rect 6335 -499 6336 -489
rect 6351 -499 6364 -489
rect 6378 -499 6379 -489
rect 6394 -499 6407 -489
rect 6422 -499 6452 -485
rect 6496 -499 6538 -485
rect 6562 -488 6569 -481
rect 6572 -489 6751 -479
rect 6545 -499 6575 -489
rect 6577 -499 6730 -489
rect 6738 -499 6768 -489
rect 6772 -499 6802 -485
rect 6830 -499 6843 -461
rect 6915 -455 6950 -447
rect 6915 -481 6916 -455
rect 6923 -481 6950 -455
rect 6858 -499 6888 -485
rect 6915 -489 6950 -481
rect 6915 -499 6916 -489
rect 6931 -499 6944 -489
rect -2 -504 6944 -499
rect -1 -512 6944 -504
rect 14 -542 27 -512
rect 42 -530 72 -512
rect 115 -526 129 -512
rect 165 -526 385 -512
rect 116 -528 129 -526
rect 82 -540 97 -528
rect 79 -542 101 -540
rect 106 -542 136 -528
rect 197 -530 350 -526
rect 179 -542 371 -530
rect 414 -542 444 -528
rect 450 -542 463 -512
rect 478 -530 508 -512
rect 551 -542 564 -512
rect 594 -542 607 -512
rect 622 -530 652 -512
rect 695 -526 709 -512
rect 745 -526 965 -512
rect 696 -528 709 -526
rect 662 -540 677 -528
rect 659 -542 681 -540
rect 686 -542 716 -528
rect 777 -530 930 -526
rect 759 -542 951 -530
rect 994 -542 1024 -528
rect 1030 -542 1043 -512
rect 1058 -530 1088 -512
rect 1131 -542 1144 -512
rect 1174 -542 1187 -512
rect 1202 -530 1232 -512
rect 1275 -526 1289 -512
rect 1325 -526 1545 -512
rect 1276 -528 1289 -526
rect 1242 -540 1257 -528
rect 1239 -542 1261 -540
rect 1266 -542 1296 -528
rect 1357 -530 1510 -526
rect 1339 -542 1531 -530
rect 1574 -542 1604 -528
rect 1610 -542 1623 -512
rect 1638 -530 1668 -512
rect 1711 -542 1724 -512
rect 1754 -542 1767 -512
rect 1782 -530 1812 -512
rect 1855 -526 1869 -512
rect 1905 -526 2125 -512
rect 1856 -528 1869 -526
rect 1822 -540 1837 -528
rect 1819 -542 1841 -540
rect 1846 -542 1876 -528
rect 1937 -530 2090 -526
rect 1919 -542 2111 -530
rect 2154 -542 2184 -528
rect 2190 -542 2203 -512
rect 2218 -530 2248 -512
rect 2291 -542 2304 -512
rect 2334 -542 2347 -512
rect 2362 -530 2392 -512
rect 2435 -526 2449 -512
rect 2485 -526 2705 -512
rect 2436 -528 2449 -526
rect 2402 -540 2417 -528
rect 2399 -542 2421 -540
rect 2426 -542 2456 -528
rect 2517 -530 2670 -526
rect 2499 -542 2691 -530
rect 2734 -542 2764 -528
rect 2770 -542 2783 -512
rect 2798 -530 2828 -512
rect 2871 -542 2884 -512
rect 2914 -542 2927 -512
rect 2942 -530 2972 -512
rect 3015 -526 3029 -512
rect 3065 -526 3285 -512
rect 3016 -528 3029 -526
rect 2982 -540 2997 -528
rect 2979 -542 3001 -540
rect 3006 -542 3036 -528
rect 3097 -530 3250 -526
rect 3079 -542 3271 -530
rect 3314 -542 3344 -528
rect 3350 -542 3363 -512
rect 3378 -530 3408 -512
rect 3451 -542 3464 -512
rect 3494 -542 3507 -512
rect 3522 -530 3552 -512
rect 3595 -526 3609 -512
rect 3645 -526 3865 -512
rect 3596 -528 3609 -526
rect 3562 -540 3577 -528
rect 3559 -542 3581 -540
rect 3586 -542 3616 -528
rect 3677 -530 3830 -526
rect 3659 -542 3851 -530
rect 3894 -542 3924 -528
rect 3930 -542 3943 -512
rect 3958 -530 3988 -512
rect 4031 -542 4044 -512
rect 4074 -542 4087 -512
rect 4102 -530 4132 -512
rect 4175 -526 4189 -512
rect 4225 -526 4445 -512
rect 4176 -528 4189 -526
rect 4142 -540 4157 -528
rect 4139 -542 4161 -540
rect 4166 -542 4196 -528
rect 4257 -530 4410 -526
rect 4239 -542 4431 -530
rect 4474 -542 4504 -528
rect 4510 -542 4523 -512
rect 4538 -530 4568 -512
rect 4611 -513 6944 -512
rect 4611 -542 4624 -513
rect -1 -543 4624 -542
rect 4654 -543 4667 -513
rect 4682 -531 4712 -513
rect 4756 -529 4769 -513
rect 4805 -527 5025 -513
rect 4722 -541 4737 -529
rect 4719 -543 4741 -541
rect 4746 -543 4776 -529
rect 4837 -531 4990 -527
rect 4819 -543 5011 -531
rect 5054 -543 5084 -529
rect 5090 -543 5103 -513
rect 5118 -531 5148 -513
rect 5191 -543 5204 -513
rect 5234 -543 5247 -513
rect 5262 -531 5292 -513
rect 5336 -529 5349 -513
rect 5385 -527 5605 -513
rect 5302 -541 5317 -529
rect 5299 -543 5321 -541
rect 5326 -543 5356 -529
rect 5417 -531 5570 -527
rect 5399 -543 5591 -531
rect 5634 -543 5664 -529
rect 5670 -543 5683 -513
rect 5698 -531 5728 -513
rect 5771 -543 5784 -513
rect 5814 -543 5827 -513
rect 5842 -531 5872 -513
rect 5916 -529 5929 -513
rect 5965 -527 6185 -513
rect 5882 -541 5897 -529
rect 5879 -543 5901 -541
rect 5906 -543 5936 -529
rect 5997 -531 6150 -527
rect 5979 -543 6171 -531
rect 6214 -543 6244 -529
rect 6250 -543 6263 -513
rect 6278 -531 6308 -513
rect 6351 -543 6364 -513
rect 6394 -543 6407 -513
rect 6422 -531 6452 -513
rect 6496 -529 6509 -513
rect 6545 -527 6765 -513
rect 6462 -541 6477 -529
rect 6459 -543 6481 -541
rect 6486 -543 6516 -529
rect 6577 -531 6730 -527
rect 6559 -543 6751 -531
rect 6794 -543 6824 -529
rect 6830 -543 6843 -513
rect 6858 -531 6888 -513
rect 6931 -543 6944 -513
rect -1 -556 6944 -543
rect 14 -660 27 -556
rect 72 -578 73 -568
rect 88 -578 101 -568
rect 72 -582 101 -578
rect 106 -582 136 -556
rect 154 -570 170 -568
rect 242 -570 295 -556
rect 243 -572 307 -570
rect 350 -572 365 -556
rect 414 -559 444 -556
rect 414 -562 450 -559
rect 380 -570 396 -568
rect 154 -582 169 -578
rect 72 -584 169 -582
rect 197 -584 365 -572
rect 381 -582 396 -578
rect 414 -581 453 -562
rect 472 -568 479 -567
rect 478 -575 479 -568
rect 462 -578 463 -575
rect 478 -578 491 -575
rect 414 -582 444 -581
rect 453 -582 459 -581
rect 462 -582 491 -578
rect 381 -583 491 -582
rect 381 -584 497 -583
rect 56 -592 107 -584
rect 56 -604 81 -592
rect 88 -604 107 -592
rect 138 -592 188 -584
rect 138 -600 154 -592
rect 161 -594 188 -592
rect 197 -594 418 -584
rect 161 -604 418 -594
rect 447 -592 497 -584
rect 447 -601 463 -592
rect 56 -612 107 -604
rect 154 -612 418 -604
rect 444 -604 463 -601
rect 470 -604 497 -592
rect 444 -612 497 -604
rect 72 -620 73 -612
rect 88 -620 101 -612
rect 72 -628 88 -620
rect 69 -635 88 -632
rect 69 -644 91 -635
rect 42 -654 91 -644
rect 42 -660 72 -654
rect 91 -659 96 -654
rect 14 -676 88 -660
rect 106 -668 136 -612
rect 171 -622 379 -612
rect 414 -616 459 -612
rect 462 -613 463 -612
rect 478 -613 491 -612
rect 197 -652 386 -622
rect 212 -655 386 -652
rect 205 -658 386 -655
rect 14 -678 27 -676
rect 42 -678 76 -676
rect 14 -694 88 -678
rect 115 -682 128 -668
rect 143 -682 159 -666
rect 205 -671 216 -658
rect -2 -716 -1 -700
rect 14 -716 27 -694
rect 42 -716 72 -694
rect 115 -698 177 -682
rect 205 -689 216 -673
rect 221 -678 231 -658
rect 241 -678 255 -658
rect 258 -671 267 -658
rect 283 -671 292 -658
rect 221 -689 255 -678
rect 258 -689 267 -673
rect 283 -689 292 -673
rect 299 -678 309 -658
rect 319 -678 333 -658
rect 334 -671 345 -658
rect 299 -689 333 -678
rect 334 -689 345 -673
rect 391 -682 407 -666
rect 414 -668 444 -616
rect 478 -620 479 -613
rect 463 -628 479 -620
rect 450 -660 463 -641
rect 478 -660 508 -644
rect 450 -676 524 -660
rect 450 -678 463 -676
rect 478 -678 512 -676
rect 115 -700 128 -698
rect 143 -700 177 -698
rect 115 -716 177 -700
rect 221 -705 237 -702
rect 299 -705 329 -694
rect 377 -698 423 -682
rect 450 -694 524 -678
rect 377 -700 411 -698
rect 376 -716 423 -700
rect 450 -716 463 -694
rect 478 -716 508 -694
rect 535 -716 536 -700
rect 551 -716 564 -556
rect 594 -660 607 -556
rect 652 -578 653 -568
rect 668 -578 681 -568
rect 652 -582 681 -578
rect 686 -582 716 -556
rect 734 -570 750 -568
rect 822 -570 875 -556
rect 823 -572 887 -570
rect 930 -572 945 -556
rect 994 -559 1024 -556
rect 994 -562 1030 -559
rect 960 -570 976 -568
rect 734 -582 749 -578
rect 652 -584 749 -582
rect 777 -584 945 -572
rect 961 -582 976 -578
rect 994 -581 1033 -562
rect 1052 -568 1059 -567
rect 1058 -575 1059 -568
rect 1042 -578 1043 -575
rect 1058 -578 1071 -575
rect 994 -582 1024 -581
rect 1033 -582 1039 -581
rect 1042 -582 1071 -578
rect 961 -583 1071 -582
rect 961 -584 1077 -583
rect 636 -592 687 -584
rect 636 -604 661 -592
rect 668 -604 687 -592
rect 718 -592 768 -584
rect 718 -600 734 -592
rect 741 -594 768 -592
rect 777 -594 998 -584
rect 741 -604 998 -594
rect 1027 -592 1077 -584
rect 1027 -601 1043 -592
rect 636 -612 687 -604
rect 734 -612 998 -604
rect 1024 -604 1043 -601
rect 1050 -604 1077 -592
rect 1024 -612 1077 -604
rect 652 -620 653 -612
rect 668 -620 681 -612
rect 652 -628 668 -620
rect 649 -635 668 -632
rect 649 -644 671 -635
rect 622 -654 671 -644
rect 622 -660 652 -654
rect 671 -659 676 -654
rect 594 -676 668 -660
rect 686 -668 716 -612
rect 751 -622 959 -612
rect 994 -616 1039 -612
rect 1042 -613 1043 -612
rect 1058 -613 1071 -612
rect 777 -652 966 -622
rect 792 -655 966 -652
rect 785 -658 966 -655
rect 594 -678 607 -676
rect 622 -678 656 -676
rect 594 -694 668 -678
rect 695 -682 708 -668
rect 723 -682 739 -666
rect 785 -671 796 -658
rect 578 -716 579 -700
rect 594 -716 607 -694
rect 622 -716 652 -694
rect 695 -698 757 -682
rect 785 -689 796 -673
rect 801 -678 811 -658
rect 821 -678 835 -658
rect 838 -671 847 -658
rect 863 -671 872 -658
rect 801 -689 835 -678
rect 838 -689 847 -673
rect 863 -689 872 -673
rect 879 -678 889 -658
rect 899 -678 913 -658
rect 914 -671 925 -658
rect 879 -689 913 -678
rect 914 -689 925 -673
rect 971 -682 987 -666
rect 994 -668 1024 -616
rect 1058 -620 1059 -613
rect 1043 -628 1059 -620
rect 1030 -660 1043 -641
rect 1058 -660 1088 -644
rect 1030 -676 1104 -660
rect 1030 -678 1043 -676
rect 1058 -678 1092 -676
rect 695 -700 708 -698
rect 723 -700 757 -698
rect 695 -716 757 -700
rect 801 -705 817 -702
rect 879 -705 909 -694
rect 957 -698 1003 -682
rect 1030 -694 1104 -678
rect 957 -700 991 -698
rect 956 -716 1003 -700
rect 1030 -716 1043 -694
rect 1058 -716 1088 -694
rect 1115 -716 1116 -700
rect 1131 -716 1144 -556
rect 1174 -660 1187 -556
rect 1232 -578 1233 -568
rect 1248 -578 1261 -568
rect 1232 -582 1261 -578
rect 1266 -582 1296 -556
rect 1314 -570 1330 -568
rect 1402 -570 1455 -556
rect 1403 -572 1467 -570
rect 1510 -572 1525 -556
rect 1574 -559 1604 -556
rect 1574 -562 1610 -559
rect 1540 -570 1556 -568
rect 1314 -582 1329 -578
rect 1232 -584 1329 -582
rect 1357 -584 1525 -572
rect 1541 -582 1556 -578
rect 1574 -581 1613 -562
rect 1632 -568 1639 -567
rect 1638 -575 1639 -568
rect 1622 -578 1623 -575
rect 1638 -578 1651 -575
rect 1574 -582 1604 -581
rect 1613 -582 1619 -581
rect 1622 -582 1651 -578
rect 1541 -583 1651 -582
rect 1541 -584 1657 -583
rect 1216 -592 1267 -584
rect 1216 -604 1241 -592
rect 1248 -604 1267 -592
rect 1298 -592 1348 -584
rect 1298 -600 1314 -592
rect 1321 -594 1348 -592
rect 1357 -594 1578 -584
rect 1321 -604 1578 -594
rect 1607 -592 1657 -584
rect 1607 -601 1623 -592
rect 1216 -612 1267 -604
rect 1314 -612 1578 -604
rect 1604 -604 1623 -601
rect 1630 -604 1657 -592
rect 1604 -612 1657 -604
rect 1232 -620 1233 -612
rect 1248 -620 1261 -612
rect 1232 -628 1248 -620
rect 1229 -635 1248 -632
rect 1229 -644 1251 -635
rect 1202 -654 1251 -644
rect 1202 -660 1232 -654
rect 1251 -659 1256 -654
rect 1174 -676 1248 -660
rect 1266 -668 1296 -612
rect 1331 -622 1539 -612
rect 1574 -616 1619 -612
rect 1622 -613 1623 -612
rect 1638 -613 1651 -612
rect 1357 -652 1546 -622
rect 1372 -655 1546 -652
rect 1365 -658 1546 -655
rect 1174 -678 1187 -676
rect 1202 -678 1236 -676
rect 1174 -694 1248 -678
rect 1275 -682 1288 -668
rect 1303 -682 1319 -666
rect 1365 -671 1376 -658
rect 1158 -716 1159 -700
rect 1174 -716 1187 -694
rect 1202 -716 1232 -694
rect 1275 -698 1337 -682
rect 1365 -689 1376 -673
rect 1381 -678 1391 -658
rect 1401 -678 1415 -658
rect 1418 -671 1427 -658
rect 1443 -671 1452 -658
rect 1381 -689 1415 -678
rect 1418 -689 1427 -673
rect 1443 -689 1452 -673
rect 1459 -678 1469 -658
rect 1479 -678 1493 -658
rect 1494 -671 1505 -658
rect 1459 -689 1493 -678
rect 1494 -689 1505 -673
rect 1551 -682 1567 -666
rect 1574 -668 1604 -616
rect 1638 -620 1639 -613
rect 1623 -628 1639 -620
rect 1610 -660 1623 -641
rect 1638 -660 1668 -644
rect 1610 -676 1684 -660
rect 1610 -678 1623 -676
rect 1638 -678 1672 -676
rect 1275 -700 1288 -698
rect 1303 -700 1337 -698
rect 1275 -716 1337 -700
rect 1381 -705 1397 -702
rect 1459 -705 1489 -694
rect 1537 -698 1583 -682
rect 1610 -694 1684 -678
rect 1537 -700 1571 -698
rect 1536 -716 1583 -700
rect 1610 -716 1623 -694
rect 1638 -716 1668 -694
rect 1695 -716 1696 -700
rect 1711 -716 1724 -556
rect 1754 -660 1767 -556
rect 1812 -578 1813 -568
rect 1828 -578 1841 -568
rect 1812 -582 1841 -578
rect 1846 -582 1876 -556
rect 1894 -570 1910 -568
rect 1982 -570 2035 -556
rect 1983 -572 2047 -570
rect 2090 -572 2105 -556
rect 2154 -559 2184 -556
rect 2154 -562 2190 -559
rect 2120 -570 2136 -568
rect 1894 -582 1909 -578
rect 1812 -584 1909 -582
rect 1937 -584 2105 -572
rect 2121 -582 2136 -578
rect 2154 -581 2193 -562
rect 2212 -568 2219 -567
rect 2218 -575 2219 -568
rect 2202 -578 2203 -575
rect 2218 -578 2231 -575
rect 2154 -582 2184 -581
rect 2193 -582 2199 -581
rect 2202 -582 2231 -578
rect 2121 -583 2231 -582
rect 2121 -584 2237 -583
rect 1796 -592 1847 -584
rect 1796 -604 1821 -592
rect 1828 -604 1847 -592
rect 1878 -592 1928 -584
rect 1878 -600 1894 -592
rect 1901 -594 1928 -592
rect 1937 -594 2158 -584
rect 1901 -604 2158 -594
rect 2187 -592 2237 -584
rect 2187 -601 2203 -592
rect 1796 -612 1847 -604
rect 1894 -612 2158 -604
rect 2184 -604 2203 -601
rect 2210 -604 2237 -592
rect 2184 -612 2237 -604
rect 1812 -620 1813 -612
rect 1828 -620 1841 -612
rect 1812 -628 1828 -620
rect 1809 -635 1828 -632
rect 1809 -644 1831 -635
rect 1782 -654 1831 -644
rect 1782 -660 1812 -654
rect 1831 -659 1836 -654
rect 1754 -676 1828 -660
rect 1846 -668 1876 -612
rect 1911 -622 2119 -612
rect 2154 -616 2199 -612
rect 2202 -613 2203 -612
rect 2218 -613 2231 -612
rect 1937 -652 2126 -622
rect 1952 -655 2126 -652
rect 1945 -658 2126 -655
rect 1754 -678 1767 -676
rect 1782 -678 1816 -676
rect 1754 -694 1828 -678
rect 1855 -682 1868 -668
rect 1883 -682 1899 -666
rect 1945 -671 1956 -658
rect 1738 -716 1739 -700
rect 1754 -716 1767 -694
rect 1782 -716 1812 -694
rect 1855 -698 1917 -682
rect 1945 -689 1956 -673
rect 1961 -678 1971 -658
rect 1981 -678 1995 -658
rect 1998 -671 2007 -658
rect 2023 -671 2032 -658
rect 1961 -689 1995 -678
rect 1998 -689 2007 -673
rect 2023 -689 2032 -673
rect 2039 -678 2049 -658
rect 2059 -678 2073 -658
rect 2074 -671 2085 -658
rect 2039 -689 2073 -678
rect 2074 -689 2085 -673
rect 2131 -682 2147 -666
rect 2154 -668 2184 -616
rect 2218 -620 2219 -613
rect 2203 -628 2219 -620
rect 2190 -660 2203 -641
rect 2218 -660 2248 -644
rect 2190 -676 2264 -660
rect 2190 -678 2203 -676
rect 2218 -678 2252 -676
rect 1855 -700 1868 -698
rect 1883 -700 1917 -698
rect 1855 -716 1917 -700
rect 1961 -705 1977 -702
rect 2039 -705 2069 -694
rect 2117 -698 2163 -682
rect 2190 -694 2264 -678
rect 2117 -700 2151 -698
rect 2116 -716 2163 -700
rect 2190 -716 2203 -694
rect 2218 -716 2248 -694
rect 2275 -716 2276 -700
rect 2291 -716 2304 -556
rect 2334 -660 2347 -556
rect 2392 -578 2393 -568
rect 2408 -578 2421 -568
rect 2392 -582 2421 -578
rect 2426 -582 2456 -556
rect 2474 -570 2490 -568
rect 2562 -570 2615 -556
rect 2563 -572 2627 -570
rect 2670 -572 2685 -556
rect 2734 -559 2764 -556
rect 2734 -562 2770 -559
rect 2700 -570 2716 -568
rect 2474 -582 2489 -578
rect 2392 -584 2489 -582
rect 2517 -584 2685 -572
rect 2701 -582 2716 -578
rect 2734 -581 2773 -562
rect 2792 -568 2799 -567
rect 2798 -575 2799 -568
rect 2782 -578 2783 -575
rect 2798 -578 2811 -575
rect 2734 -582 2764 -581
rect 2773 -582 2779 -581
rect 2782 -582 2811 -578
rect 2701 -583 2811 -582
rect 2701 -584 2817 -583
rect 2376 -592 2427 -584
rect 2376 -604 2401 -592
rect 2408 -604 2427 -592
rect 2458 -592 2508 -584
rect 2458 -600 2474 -592
rect 2481 -594 2508 -592
rect 2517 -594 2738 -584
rect 2481 -604 2738 -594
rect 2767 -592 2817 -584
rect 2767 -601 2783 -592
rect 2376 -612 2427 -604
rect 2474 -612 2738 -604
rect 2764 -604 2783 -601
rect 2790 -604 2817 -592
rect 2764 -612 2817 -604
rect 2392 -620 2393 -612
rect 2408 -620 2421 -612
rect 2392 -628 2408 -620
rect 2389 -635 2408 -632
rect 2389 -644 2411 -635
rect 2362 -654 2411 -644
rect 2362 -660 2392 -654
rect 2411 -659 2416 -654
rect 2334 -676 2408 -660
rect 2426 -668 2456 -612
rect 2491 -622 2699 -612
rect 2734 -616 2779 -612
rect 2782 -613 2783 -612
rect 2798 -613 2811 -612
rect 2517 -652 2706 -622
rect 2532 -655 2706 -652
rect 2525 -658 2706 -655
rect 2334 -678 2347 -676
rect 2362 -678 2396 -676
rect 2334 -694 2408 -678
rect 2435 -682 2448 -668
rect 2463 -682 2479 -666
rect 2525 -671 2536 -658
rect 2318 -716 2319 -700
rect 2334 -716 2347 -694
rect 2362 -716 2392 -694
rect 2435 -698 2497 -682
rect 2525 -689 2536 -673
rect 2541 -678 2551 -658
rect 2561 -678 2575 -658
rect 2578 -671 2587 -658
rect 2603 -671 2612 -658
rect 2541 -689 2575 -678
rect 2578 -689 2587 -673
rect 2603 -689 2612 -673
rect 2619 -678 2629 -658
rect 2639 -678 2653 -658
rect 2654 -671 2665 -658
rect 2619 -689 2653 -678
rect 2654 -689 2665 -673
rect 2711 -682 2727 -666
rect 2734 -668 2764 -616
rect 2798 -620 2799 -613
rect 2783 -628 2799 -620
rect 2770 -660 2783 -641
rect 2798 -660 2828 -644
rect 2770 -676 2844 -660
rect 2770 -678 2783 -676
rect 2798 -678 2832 -676
rect 2435 -700 2448 -698
rect 2463 -700 2497 -698
rect 2435 -716 2497 -700
rect 2541 -705 2557 -702
rect 2619 -705 2649 -694
rect 2697 -698 2743 -682
rect 2770 -694 2844 -678
rect 2697 -700 2731 -698
rect 2696 -716 2743 -700
rect 2770 -716 2783 -694
rect 2798 -716 2828 -694
rect 2855 -716 2856 -700
rect 2871 -716 2884 -556
rect 2914 -660 2927 -556
rect 2972 -578 2973 -568
rect 2988 -578 3001 -568
rect 2972 -582 3001 -578
rect 3006 -582 3036 -556
rect 3054 -570 3070 -568
rect 3142 -570 3195 -556
rect 3143 -572 3205 -570
rect 3250 -572 3265 -556
rect 3314 -559 3344 -556
rect 3314 -562 3350 -559
rect 3280 -570 3296 -568
rect 3054 -582 3069 -578
rect 2972 -584 3069 -582
rect 3097 -584 3265 -572
rect 3281 -582 3296 -578
rect 3314 -581 3353 -562
rect 3372 -568 3379 -567
rect 3378 -575 3379 -568
rect 3362 -578 3363 -575
rect 3378 -578 3391 -575
rect 3314 -582 3344 -581
rect 3353 -582 3359 -581
rect 3362 -582 3391 -578
rect 3281 -583 3391 -582
rect 3281 -584 3397 -583
rect 2956 -592 3007 -584
rect 2956 -604 2981 -592
rect 2988 -604 3007 -592
rect 3038 -592 3088 -584
rect 3038 -600 3054 -592
rect 3061 -594 3088 -592
rect 3097 -594 3318 -584
rect 3061 -604 3318 -594
rect 3347 -592 3397 -584
rect 3347 -601 3363 -592
rect 2956 -612 3007 -604
rect 3054 -612 3318 -604
rect 3344 -604 3363 -601
rect 3370 -604 3397 -592
rect 3344 -612 3397 -604
rect 2972 -620 2973 -612
rect 2988 -620 3001 -612
rect 2972 -628 2988 -620
rect 2969 -635 2988 -632
rect 2969 -644 2991 -635
rect 2942 -654 2991 -644
rect 2942 -660 2972 -654
rect 2991 -659 2996 -654
rect 2914 -676 2988 -660
rect 3006 -668 3036 -612
rect 3071 -622 3279 -612
rect 3314 -616 3359 -612
rect 3362 -613 3363 -612
rect 3378 -613 3391 -612
rect 3097 -652 3286 -622
rect 3112 -655 3286 -652
rect 3105 -658 3286 -655
rect 2914 -678 2927 -676
rect 2942 -678 2976 -676
rect 2914 -694 2988 -678
rect 3015 -682 3028 -668
rect 3043 -682 3059 -666
rect 3105 -671 3116 -658
rect 2898 -716 2899 -700
rect 2914 -716 2927 -694
rect 2942 -716 2972 -694
rect 3015 -698 3077 -682
rect 3105 -689 3116 -673
rect 3121 -678 3131 -658
rect 3141 -678 3155 -658
rect 3158 -671 3167 -658
rect 3183 -671 3192 -658
rect 3121 -689 3155 -678
rect 3158 -689 3167 -673
rect 3183 -689 3192 -673
rect 3199 -678 3209 -658
rect 3219 -678 3233 -658
rect 3234 -671 3245 -658
rect 3199 -689 3233 -678
rect 3234 -689 3245 -673
rect 3291 -682 3307 -666
rect 3314 -668 3344 -616
rect 3378 -620 3379 -613
rect 3363 -628 3379 -620
rect 3350 -660 3363 -641
rect 3378 -660 3408 -644
rect 3350 -676 3424 -660
rect 3350 -678 3363 -676
rect 3378 -678 3412 -676
rect 3015 -700 3028 -698
rect 3043 -700 3077 -698
rect 3015 -716 3077 -700
rect 3121 -705 3137 -702
rect 3199 -705 3229 -694
rect 3277 -698 3323 -682
rect 3350 -694 3424 -678
rect 3277 -700 3311 -698
rect 3276 -716 3323 -700
rect 3350 -716 3363 -694
rect 3378 -716 3408 -694
rect 3435 -716 3436 -700
rect 3451 -716 3464 -556
rect 3494 -660 3507 -556
rect 3552 -578 3553 -568
rect 3568 -578 3581 -568
rect 3552 -582 3581 -578
rect 3586 -582 3616 -556
rect 3634 -570 3650 -568
rect 3722 -570 3775 -556
rect 3723 -572 3787 -570
rect 3830 -572 3845 -556
rect 3894 -559 3924 -556
rect 3894 -562 3930 -559
rect 3860 -570 3876 -568
rect 3634 -582 3649 -578
rect 3552 -584 3649 -582
rect 3677 -584 3845 -572
rect 3861 -582 3876 -578
rect 3894 -581 3933 -562
rect 3952 -568 3959 -567
rect 3958 -575 3959 -568
rect 3942 -578 3943 -575
rect 3958 -578 3971 -575
rect 3894 -582 3924 -581
rect 3933 -582 3939 -581
rect 3942 -582 3971 -578
rect 3861 -583 3971 -582
rect 3861 -584 3977 -583
rect 3536 -592 3587 -584
rect 3536 -604 3561 -592
rect 3568 -604 3587 -592
rect 3618 -592 3668 -584
rect 3618 -600 3634 -592
rect 3641 -594 3668 -592
rect 3677 -594 3898 -584
rect 3641 -604 3898 -594
rect 3927 -592 3977 -584
rect 3927 -601 3943 -592
rect 3536 -612 3587 -604
rect 3634 -612 3898 -604
rect 3924 -604 3943 -601
rect 3950 -604 3977 -592
rect 3924 -612 3977 -604
rect 3552 -620 3553 -612
rect 3568 -620 3581 -612
rect 3552 -628 3568 -620
rect 3549 -635 3568 -632
rect 3549 -644 3571 -635
rect 3522 -654 3571 -644
rect 3522 -660 3552 -654
rect 3571 -659 3576 -654
rect 3494 -676 3568 -660
rect 3586 -668 3616 -612
rect 3651 -622 3859 -612
rect 3894 -616 3939 -612
rect 3942 -613 3943 -612
rect 3958 -613 3971 -612
rect 3677 -652 3866 -622
rect 3692 -655 3866 -652
rect 3685 -658 3866 -655
rect 3494 -678 3507 -676
rect 3522 -678 3556 -676
rect 3494 -694 3568 -678
rect 3595 -682 3608 -668
rect 3623 -682 3639 -666
rect 3685 -671 3696 -658
rect 3478 -716 3479 -700
rect 3494 -716 3507 -694
rect 3522 -716 3552 -694
rect 3595 -698 3657 -682
rect 3685 -689 3696 -673
rect 3701 -678 3711 -658
rect 3721 -678 3735 -658
rect 3738 -671 3747 -658
rect 3763 -671 3772 -658
rect 3701 -689 3735 -678
rect 3738 -689 3747 -673
rect 3763 -689 3772 -673
rect 3779 -678 3789 -658
rect 3799 -678 3813 -658
rect 3814 -671 3825 -658
rect 3779 -689 3813 -678
rect 3814 -689 3825 -673
rect 3871 -682 3887 -666
rect 3894 -668 3924 -616
rect 3958 -620 3959 -613
rect 3943 -628 3959 -620
rect 3930 -660 3943 -641
rect 3958 -660 3988 -644
rect 3930 -676 4004 -660
rect 3930 -678 3943 -676
rect 3958 -678 3992 -676
rect 3595 -700 3608 -698
rect 3623 -700 3657 -698
rect 3595 -716 3657 -700
rect 3701 -705 3717 -702
rect 3779 -705 3809 -694
rect 3857 -698 3903 -682
rect 3930 -694 4004 -678
rect 3857 -700 3891 -698
rect 3856 -716 3903 -700
rect 3930 -716 3943 -694
rect 3958 -716 3988 -694
rect 4015 -716 4016 -700
rect 4031 -716 4044 -556
rect 4074 -660 4087 -556
rect 4132 -578 4133 -568
rect 4148 -578 4161 -568
rect 4132 -582 4161 -578
rect 4166 -582 4196 -556
rect 4214 -570 4230 -568
rect 4302 -570 4355 -556
rect 4303 -572 4367 -570
rect 4410 -572 4425 -556
rect 4474 -559 4504 -556
rect 4611 -557 6944 -556
rect 4474 -562 4510 -559
rect 4440 -570 4456 -568
rect 4214 -582 4229 -578
rect 4132 -584 4229 -582
rect 4257 -584 4425 -572
rect 4441 -582 4456 -578
rect 4474 -581 4513 -562
rect 4532 -568 4539 -567
rect 4538 -575 4539 -568
rect 4522 -578 4523 -575
rect 4538 -578 4551 -575
rect 4474 -582 4504 -581
rect 4513 -582 4519 -581
rect 4522 -582 4551 -578
rect 4441 -583 4551 -582
rect 4441 -584 4557 -583
rect 4116 -592 4167 -584
rect 4116 -604 4141 -592
rect 4148 -604 4167 -592
rect 4198 -592 4248 -584
rect 4198 -600 4214 -592
rect 4221 -594 4248 -592
rect 4257 -594 4478 -584
rect 4221 -604 4478 -594
rect 4507 -592 4557 -584
rect 4507 -601 4523 -592
rect 4116 -612 4167 -604
rect 4214 -612 4478 -604
rect 4504 -604 4523 -601
rect 4530 -604 4557 -592
rect 4504 -612 4557 -604
rect 4132 -620 4133 -612
rect 4148 -620 4161 -612
rect 4132 -628 4148 -620
rect 4129 -635 4148 -632
rect 4129 -644 4151 -635
rect 4102 -654 4151 -644
rect 4102 -660 4132 -654
rect 4151 -659 4156 -654
rect 4074 -676 4148 -660
rect 4166 -668 4196 -612
rect 4231 -622 4439 -612
rect 4474 -616 4519 -612
rect 4522 -613 4523 -612
rect 4538 -613 4551 -612
rect 4257 -652 4446 -622
rect 4272 -655 4446 -652
rect 4265 -658 4446 -655
rect 4074 -678 4087 -676
rect 4102 -678 4136 -676
rect 4074 -694 4148 -678
rect 4175 -682 4188 -668
rect 4203 -682 4219 -666
rect 4265 -671 4276 -658
rect 4058 -716 4059 -700
rect 4074 -716 4087 -694
rect 4102 -716 4132 -694
rect 4175 -698 4237 -682
rect 4265 -689 4276 -673
rect 4281 -678 4291 -658
rect 4301 -678 4315 -658
rect 4318 -671 4327 -658
rect 4343 -671 4352 -658
rect 4281 -689 4315 -678
rect 4318 -689 4327 -673
rect 4343 -689 4352 -673
rect 4359 -678 4369 -658
rect 4379 -678 4393 -658
rect 4394 -671 4405 -658
rect 4359 -689 4393 -678
rect 4394 -689 4405 -673
rect 4451 -682 4467 -666
rect 4474 -668 4504 -616
rect 4538 -620 4539 -613
rect 4523 -628 4539 -620
rect 4510 -660 4523 -641
rect 4538 -660 4568 -644
rect 4510 -676 4584 -660
rect 4510 -678 4523 -676
rect 4538 -678 4572 -676
rect 4175 -700 4188 -698
rect 4203 -700 4237 -698
rect 4175 -716 4237 -700
rect 4281 -705 4297 -702
rect 4359 -705 4389 -694
rect 4437 -698 4483 -682
rect 4510 -694 4584 -678
rect 4437 -700 4471 -698
rect 4436 -716 4483 -700
rect 4510 -716 4523 -694
rect 4538 -716 4568 -694
rect 4595 -716 4596 -700
rect 4611 -716 4624 -557
rect 4654 -661 4667 -557
rect 4712 -579 4713 -569
rect 4733 -571 4741 -569
rect 4731 -573 4741 -571
rect 4729 -575 4741 -573
rect 4728 -579 4741 -575
rect 4712 -583 4741 -579
rect 4746 -583 4776 -557
rect 4794 -571 4810 -569
rect 4882 -571 4933 -557
rect 4883 -573 4947 -571
rect 4990 -573 5005 -557
rect 5054 -560 5084 -557
rect 5054 -563 5090 -560
rect 5020 -571 5036 -569
rect 4794 -583 4809 -579
rect 4712 -585 4809 -583
rect 4837 -585 5005 -573
rect 5021 -583 5036 -579
rect 5054 -582 5093 -563
rect 5112 -569 5119 -568
rect 5118 -576 5119 -569
rect 5102 -579 5103 -576
rect 5118 -579 5131 -576
rect 5054 -583 5084 -582
rect 5093 -583 5099 -582
rect 5102 -583 5131 -579
rect 5021 -584 5131 -583
rect 5021 -585 5137 -584
rect 4696 -593 4747 -585
rect 4696 -605 4721 -593
rect 4728 -605 4747 -593
rect 4778 -593 4828 -585
rect 4778 -601 4794 -593
rect 4801 -595 4828 -593
rect 4837 -595 5058 -585
rect 4801 -605 5058 -595
rect 5087 -593 5137 -585
rect 5087 -602 5103 -593
rect 4696 -613 4747 -605
rect 4794 -613 5058 -605
rect 5084 -605 5103 -602
rect 5110 -605 5137 -593
rect 5084 -613 5137 -605
rect 4712 -621 4713 -613
rect 4728 -621 4741 -613
rect 4712 -629 4728 -621
rect 4709 -636 4728 -633
rect 4709 -645 4731 -636
rect 4682 -655 4731 -645
rect 4682 -661 4712 -655
rect 4731 -660 4736 -655
rect 4654 -677 4728 -661
rect 4746 -669 4776 -613
rect 4811 -623 5019 -613
rect 5054 -617 5099 -613
rect 5102 -614 5103 -613
rect 5118 -614 5131 -613
rect 4837 -653 5026 -623
rect 4852 -656 5026 -653
rect 4845 -659 5026 -656
rect 4654 -679 4667 -677
rect 4682 -679 4716 -677
rect 4654 -695 4728 -679
rect 4755 -683 4768 -669
rect 4783 -683 4799 -667
rect 4845 -672 4856 -659
rect -8 -724 33 -716
rect -8 -750 7 -724
rect 14 -750 33 -724
rect 97 -728 159 -716
rect 171 -728 246 -716
rect 304 -728 379 -716
rect 391 -728 422 -716
rect 428 -728 463 -716
rect 97 -730 259 -728
rect -8 -758 33 -750
rect 115 -754 128 -730
rect 143 -732 158 -730
rect -2 -768 -1 -758
rect 14 -768 27 -758
rect 42 -768 72 -754
rect 115 -768 158 -754
rect 182 -757 189 -750
rect 192 -754 259 -730
rect 291 -730 463 -728
rect 261 -752 289 -748
rect 291 -752 371 -730
rect 392 -732 407 -730
rect 261 -754 371 -752
rect 192 -758 371 -754
rect 165 -768 195 -758
rect 197 -768 350 -758
rect 358 -768 388 -758
rect 392 -768 422 -754
rect 450 -768 463 -730
rect 535 -724 570 -716
rect 535 -750 536 -724
rect 543 -750 570 -724
rect 478 -768 508 -754
rect 535 -758 570 -750
rect 572 -724 613 -716
rect 572 -750 587 -724
rect 594 -750 613 -724
rect 677 -728 739 -716
rect 751 -728 826 -716
rect 884 -728 959 -716
rect 971 -728 1002 -716
rect 1008 -728 1043 -716
rect 677 -730 839 -728
rect 572 -758 613 -750
rect 695 -754 708 -730
rect 723 -732 738 -730
rect 535 -768 536 -758
rect 551 -768 564 -758
rect 578 -768 579 -758
rect 594 -768 607 -758
rect 622 -768 652 -754
rect 695 -768 738 -754
rect 762 -757 769 -750
rect 772 -754 839 -730
rect 871 -730 1043 -728
rect 841 -752 869 -748
rect 871 -752 951 -730
rect 972 -732 987 -730
rect 841 -754 951 -752
rect 772 -758 951 -754
rect 745 -768 775 -758
rect 777 -768 930 -758
rect 938 -768 968 -758
rect 972 -768 1002 -754
rect 1030 -768 1043 -730
rect 1115 -724 1150 -716
rect 1115 -750 1116 -724
rect 1123 -750 1150 -724
rect 1058 -768 1088 -754
rect 1115 -758 1150 -750
rect 1152 -724 1193 -716
rect 1152 -750 1167 -724
rect 1174 -750 1193 -724
rect 1257 -728 1319 -716
rect 1331 -728 1406 -716
rect 1464 -728 1539 -716
rect 1551 -728 1582 -716
rect 1588 -728 1623 -716
rect 1257 -730 1419 -728
rect 1152 -758 1193 -750
rect 1275 -754 1288 -730
rect 1303 -732 1318 -730
rect 1115 -768 1116 -758
rect 1131 -768 1144 -758
rect 1158 -768 1159 -758
rect 1174 -768 1187 -758
rect 1202 -768 1232 -754
rect 1275 -768 1318 -754
rect 1342 -757 1349 -750
rect 1352 -754 1419 -730
rect 1451 -730 1623 -728
rect 1421 -752 1449 -748
rect 1451 -752 1531 -730
rect 1552 -732 1567 -730
rect 1421 -754 1531 -752
rect 1352 -758 1531 -754
rect 1325 -768 1355 -758
rect 1357 -768 1510 -758
rect 1518 -768 1548 -758
rect 1552 -768 1582 -754
rect 1610 -768 1623 -730
rect 1695 -724 1730 -716
rect 1695 -750 1696 -724
rect 1703 -750 1730 -724
rect 1638 -768 1668 -754
rect 1695 -758 1730 -750
rect 1732 -724 1773 -716
rect 1732 -750 1747 -724
rect 1754 -750 1773 -724
rect 1837 -728 1899 -716
rect 1911 -728 1986 -716
rect 2044 -728 2119 -716
rect 2131 -728 2162 -716
rect 2168 -728 2203 -716
rect 1837 -730 1999 -728
rect 1732 -758 1773 -750
rect 1855 -754 1868 -730
rect 1883 -732 1898 -730
rect 1695 -768 1696 -758
rect 1711 -768 1724 -758
rect 1738 -768 1739 -758
rect 1754 -768 1767 -758
rect 1782 -768 1812 -754
rect 1855 -768 1898 -754
rect 1922 -757 1929 -750
rect 1932 -754 1999 -730
rect 2031 -730 2203 -728
rect 2001 -752 2029 -748
rect 2031 -752 2111 -730
rect 2132 -732 2147 -730
rect 2001 -754 2111 -752
rect 1932 -758 2111 -754
rect 1905 -768 1935 -758
rect 1937 -768 2090 -758
rect 2098 -768 2128 -758
rect 2132 -768 2162 -754
rect 2190 -768 2203 -730
rect 2275 -724 2310 -716
rect 2275 -750 2276 -724
rect 2283 -750 2310 -724
rect 2218 -768 2248 -754
rect 2275 -758 2310 -750
rect 2312 -724 2353 -716
rect 2312 -750 2327 -724
rect 2334 -750 2353 -724
rect 2417 -728 2479 -716
rect 2491 -728 2566 -716
rect 2624 -728 2699 -716
rect 2711 -728 2742 -716
rect 2748 -728 2783 -716
rect 2417 -730 2579 -728
rect 2312 -758 2353 -750
rect 2435 -754 2448 -730
rect 2463 -732 2478 -730
rect 2275 -768 2276 -758
rect 2291 -768 2304 -758
rect 2318 -768 2319 -758
rect 2334 -768 2347 -758
rect 2362 -768 2392 -754
rect 2435 -768 2478 -754
rect 2502 -757 2509 -750
rect 2512 -754 2579 -730
rect 2611 -730 2783 -728
rect 2581 -752 2609 -748
rect 2611 -752 2691 -730
rect 2712 -732 2727 -730
rect 2581 -754 2691 -752
rect 2512 -758 2691 -754
rect 2485 -768 2515 -758
rect 2517 -768 2670 -758
rect 2678 -768 2708 -758
rect 2712 -768 2742 -754
rect 2770 -768 2783 -730
rect 2855 -724 2890 -716
rect 2855 -750 2856 -724
rect 2863 -750 2890 -724
rect 2798 -768 2828 -754
rect 2855 -758 2890 -750
rect 2892 -724 2933 -716
rect 2892 -750 2907 -724
rect 2914 -750 2933 -724
rect 2997 -728 3059 -716
rect 3071 -728 3146 -716
rect 3204 -728 3279 -716
rect 3291 -728 3322 -716
rect 3328 -728 3363 -716
rect 2997 -730 3159 -728
rect 2892 -758 2933 -750
rect 3015 -754 3028 -730
rect 3043 -732 3058 -730
rect 2855 -768 2856 -758
rect 2871 -768 2884 -758
rect 2898 -768 2899 -758
rect 2914 -768 2927 -758
rect 2942 -768 2972 -754
rect 3015 -768 3058 -754
rect 3082 -757 3089 -750
rect 3092 -754 3159 -730
rect 3191 -730 3363 -728
rect 3161 -752 3189 -748
rect 3191 -752 3271 -730
rect 3292 -732 3307 -730
rect 3161 -754 3271 -752
rect 3092 -758 3271 -754
rect 3065 -768 3095 -758
rect 3097 -768 3250 -758
rect 3258 -768 3288 -758
rect 3292 -768 3322 -754
rect 3350 -768 3363 -730
rect 3435 -724 3470 -716
rect 3435 -750 3436 -724
rect 3443 -750 3470 -724
rect 3378 -768 3408 -754
rect 3435 -758 3470 -750
rect 3472 -724 3513 -716
rect 3472 -750 3487 -724
rect 3494 -750 3513 -724
rect 3577 -728 3639 -716
rect 3651 -728 3726 -716
rect 3784 -728 3859 -716
rect 3871 -728 3902 -716
rect 3908 -728 3943 -716
rect 3577 -730 3739 -728
rect 3472 -758 3513 -750
rect 3595 -754 3608 -730
rect 3623 -732 3638 -730
rect 3435 -768 3436 -758
rect 3451 -768 3464 -758
rect 3478 -768 3479 -758
rect 3494 -768 3507 -758
rect 3522 -768 3552 -754
rect 3595 -768 3638 -754
rect 3662 -757 3669 -750
rect 3672 -754 3739 -730
rect 3771 -730 3943 -728
rect 3741 -752 3769 -748
rect 3771 -752 3851 -730
rect 3872 -732 3887 -730
rect 3741 -754 3851 -752
rect 3672 -758 3851 -754
rect 3645 -768 3675 -758
rect 3677 -768 3830 -758
rect 3838 -768 3868 -758
rect 3872 -768 3902 -754
rect 3930 -768 3943 -730
rect 4015 -724 4050 -716
rect 4015 -750 4016 -724
rect 4023 -750 4050 -724
rect 3958 -768 3988 -754
rect 4015 -758 4050 -750
rect 4052 -724 4093 -716
rect 4052 -750 4067 -724
rect 4074 -750 4093 -724
rect 4157 -728 4219 -716
rect 4231 -728 4306 -716
rect 4364 -728 4439 -716
rect 4451 -728 4482 -716
rect 4488 -728 4523 -716
rect 4157 -730 4319 -728
rect 4052 -758 4093 -750
rect 4175 -754 4188 -730
rect 4203 -732 4218 -730
rect 4015 -768 4016 -758
rect 4031 -768 4044 -758
rect 4058 -768 4059 -758
rect 4074 -768 4087 -758
rect 4102 -768 4132 -754
rect 4175 -768 4218 -754
rect 4242 -757 4249 -750
rect 4252 -754 4319 -730
rect 4351 -730 4523 -728
rect 4321 -752 4349 -748
rect 4351 -752 4431 -730
rect 4452 -732 4467 -730
rect 4321 -754 4431 -752
rect 4252 -758 4431 -754
rect 4225 -768 4255 -758
rect 4257 -768 4410 -758
rect 4418 -768 4448 -758
rect 4452 -768 4482 -754
rect 4510 -768 4523 -730
rect 4595 -724 4630 -716
rect 4638 -717 4639 -701
rect 4654 -717 4667 -695
rect 4682 -717 4712 -695
rect 4755 -699 4817 -683
rect 4845 -690 4856 -674
rect 4861 -679 4871 -659
rect 4881 -679 4895 -659
rect 4898 -672 4907 -659
rect 4923 -672 4932 -659
rect 4861 -690 4895 -679
rect 4898 -690 4907 -674
rect 4923 -690 4932 -674
rect 4939 -679 4949 -659
rect 4959 -679 4973 -659
rect 4974 -672 4985 -659
rect 4939 -690 4973 -679
rect 4974 -690 4985 -674
rect 5031 -683 5047 -667
rect 5054 -669 5084 -617
rect 5118 -621 5119 -614
rect 5103 -629 5119 -621
rect 5090 -661 5103 -642
rect 5118 -661 5148 -645
rect 5090 -677 5164 -661
rect 5090 -679 5103 -677
rect 5118 -679 5152 -677
rect 4755 -701 4768 -699
rect 4783 -701 4817 -699
rect 4755 -717 4817 -701
rect 4861 -706 4877 -703
rect 4939 -706 4969 -695
rect 5017 -699 5063 -683
rect 5090 -695 5164 -679
rect 5017 -701 5051 -699
rect 5016 -717 5063 -701
rect 5090 -717 5103 -695
rect 5118 -717 5148 -695
rect 5175 -717 5176 -701
rect 5191 -717 5204 -557
rect 5234 -661 5247 -557
rect 5292 -579 5293 -569
rect 5313 -571 5321 -569
rect 5311 -573 5321 -571
rect 5309 -575 5321 -573
rect 5308 -579 5321 -575
rect 5292 -583 5321 -579
rect 5326 -583 5356 -557
rect 5374 -571 5390 -569
rect 5462 -571 5513 -557
rect 5463 -573 5527 -571
rect 5570 -573 5585 -557
rect 5634 -560 5664 -557
rect 5634 -563 5670 -560
rect 5600 -571 5616 -569
rect 5374 -583 5389 -579
rect 5292 -585 5389 -583
rect 5417 -585 5585 -573
rect 5601 -583 5616 -579
rect 5634 -582 5673 -563
rect 5692 -569 5699 -568
rect 5698 -576 5699 -569
rect 5682 -579 5683 -576
rect 5698 -579 5711 -576
rect 5634 -583 5664 -582
rect 5673 -583 5679 -582
rect 5682 -583 5711 -579
rect 5601 -584 5711 -583
rect 5601 -585 5717 -584
rect 5276 -593 5327 -585
rect 5276 -605 5301 -593
rect 5308 -605 5327 -593
rect 5358 -593 5408 -585
rect 5358 -601 5374 -593
rect 5381 -595 5408 -593
rect 5417 -595 5638 -585
rect 5381 -605 5638 -595
rect 5667 -593 5717 -585
rect 5667 -602 5683 -593
rect 5276 -613 5327 -605
rect 5374 -613 5638 -605
rect 5664 -605 5683 -602
rect 5690 -605 5717 -593
rect 5664 -613 5717 -605
rect 5292 -621 5293 -613
rect 5308 -621 5321 -613
rect 5292 -629 5308 -621
rect 5289 -636 5308 -633
rect 5289 -645 5311 -636
rect 5262 -655 5311 -645
rect 5262 -661 5292 -655
rect 5311 -660 5316 -655
rect 5234 -677 5308 -661
rect 5326 -669 5356 -613
rect 5391 -623 5599 -613
rect 5634 -617 5679 -613
rect 5682 -614 5683 -613
rect 5698 -614 5711 -613
rect 5417 -653 5606 -623
rect 5432 -656 5606 -653
rect 5425 -659 5606 -656
rect 5234 -679 5247 -677
rect 5262 -679 5296 -677
rect 5234 -695 5308 -679
rect 5335 -683 5348 -669
rect 5363 -683 5379 -667
rect 5425 -672 5436 -659
rect 5218 -717 5219 -701
rect 5234 -717 5247 -695
rect 5262 -717 5292 -695
rect 5335 -699 5397 -683
rect 5425 -690 5436 -674
rect 5441 -679 5451 -659
rect 5461 -679 5475 -659
rect 5478 -672 5487 -659
rect 5503 -672 5512 -659
rect 5441 -690 5475 -679
rect 5478 -690 5487 -674
rect 5503 -690 5512 -674
rect 5519 -679 5529 -659
rect 5539 -679 5553 -659
rect 5554 -672 5565 -659
rect 5519 -690 5553 -679
rect 5554 -690 5565 -674
rect 5611 -683 5627 -667
rect 5634 -669 5664 -617
rect 5698 -621 5699 -614
rect 5683 -629 5699 -621
rect 5670 -661 5683 -642
rect 5698 -661 5728 -645
rect 5670 -677 5744 -661
rect 5670 -679 5683 -677
rect 5698 -679 5732 -677
rect 5335 -701 5348 -699
rect 5363 -701 5397 -699
rect 5335 -717 5397 -701
rect 5441 -706 5457 -703
rect 5519 -706 5549 -695
rect 5597 -699 5643 -683
rect 5670 -695 5744 -679
rect 5597 -701 5631 -699
rect 5596 -717 5643 -701
rect 5670 -717 5683 -695
rect 5698 -717 5728 -695
rect 5755 -717 5756 -701
rect 5771 -717 5784 -557
rect 5814 -661 5827 -557
rect 5872 -579 5873 -569
rect 5893 -571 5901 -569
rect 5891 -573 5901 -571
rect 5889 -575 5901 -573
rect 5888 -579 5901 -575
rect 5872 -583 5901 -579
rect 5906 -583 5936 -557
rect 5954 -571 5970 -569
rect 6042 -571 6093 -557
rect 6043 -573 6107 -571
rect 6150 -573 6165 -557
rect 6214 -560 6244 -557
rect 6214 -563 6250 -560
rect 6180 -571 6196 -569
rect 5954 -583 5969 -579
rect 5872 -585 5969 -583
rect 5997 -585 6165 -573
rect 6181 -583 6196 -579
rect 6214 -582 6253 -563
rect 6272 -569 6279 -568
rect 6278 -576 6279 -569
rect 6262 -579 6263 -576
rect 6278 -579 6291 -576
rect 6214 -583 6244 -582
rect 6253 -583 6259 -582
rect 6262 -583 6291 -579
rect 6181 -584 6291 -583
rect 6181 -585 6297 -584
rect 5856 -593 5907 -585
rect 5856 -605 5881 -593
rect 5888 -605 5907 -593
rect 5938 -593 5988 -585
rect 5938 -601 5954 -593
rect 5961 -595 5988 -593
rect 5997 -595 6218 -585
rect 5961 -605 6218 -595
rect 6247 -593 6297 -585
rect 6247 -602 6263 -593
rect 5856 -613 5907 -605
rect 5954 -613 6218 -605
rect 6244 -605 6263 -602
rect 6270 -605 6297 -593
rect 6244 -613 6297 -605
rect 5872 -621 5873 -613
rect 5888 -621 5901 -613
rect 5872 -629 5888 -621
rect 5869 -636 5888 -633
rect 5869 -645 5891 -636
rect 5842 -655 5891 -645
rect 5842 -661 5872 -655
rect 5891 -660 5896 -655
rect 5814 -677 5888 -661
rect 5906 -669 5936 -613
rect 5971 -623 6179 -613
rect 6214 -617 6259 -613
rect 6262 -614 6263 -613
rect 6278 -614 6291 -613
rect 5997 -653 6186 -623
rect 6012 -656 6186 -653
rect 6005 -659 6186 -656
rect 5814 -679 5827 -677
rect 5842 -679 5876 -677
rect 5814 -695 5888 -679
rect 5915 -683 5928 -669
rect 5943 -683 5959 -667
rect 6005 -672 6016 -659
rect 5798 -717 5799 -701
rect 5814 -717 5827 -695
rect 5842 -717 5872 -695
rect 5915 -699 5977 -683
rect 6005 -690 6016 -674
rect 6021 -679 6031 -659
rect 6041 -679 6055 -659
rect 6058 -672 6067 -659
rect 6083 -672 6092 -659
rect 6021 -690 6055 -679
rect 6058 -690 6067 -674
rect 6083 -690 6092 -674
rect 6099 -679 6109 -659
rect 6119 -679 6133 -659
rect 6134 -672 6145 -659
rect 6099 -690 6133 -679
rect 6134 -690 6145 -674
rect 6191 -683 6207 -667
rect 6214 -669 6244 -617
rect 6278 -621 6279 -614
rect 6263 -629 6279 -621
rect 6250 -661 6263 -642
rect 6278 -661 6308 -645
rect 6250 -677 6324 -661
rect 6250 -679 6263 -677
rect 6278 -679 6312 -677
rect 5915 -701 5928 -699
rect 5943 -701 5977 -699
rect 5915 -717 5977 -701
rect 6021 -706 6037 -703
rect 6099 -706 6129 -695
rect 6177 -699 6223 -683
rect 6250 -695 6324 -679
rect 6177 -701 6211 -699
rect 6176 -717 6223 -701
rect 6250 -717 6263 -695
rect 6278 -717 6308 -695
rect 6335 -717 6336 -701
rect 6351 -717 6364 -557
rect 6394 -661 6407 -557
rect 6452 -579 6453 -569
rect 6473 -571 6481 -569
rect 6471 -573 6481 -571
rect 6469 -575 6481 -573
rect 6468 -579 6481 -575
rect 6452 -583 6481 -579
rect 6486 -583 6516 -557
rect 6534 -571 6550 -569
rect 6622 -571 6673 -557
rect 6623 -573 6687 -571
rect 6730 -573 6745 -557
rect 6794 -560 6824 -557
rect 6794 -563 6830 -560
rect 6760 -571 6776 -569
rect 6534 -583 6549 -579
rect 6452 -585 6549 -583
rect 6577 -585 6745 -573
rect 6761 -583 6776 -579
rect 6794 -582 6833 -563
rect 6852 -569 6859 -568
rect 6858 -576 6859 -569
rect 6842 -579 6843 -576
rect 6858 -579 6871 -576
rect 6794 -583 6824 -582
rect 6833 -583 6839 -582
rect 6842 -583 6871 -579
rect 6761 -584 6871 -583
rect 6761 -585 6877 -584
rect 6436 -593 6487 -585
rect 6436 -605 6461 -593
rect 6468 -605 6487 -593
rect 6518 -593 6568 -585
rect 6518 -601 6534 -593
rect 6541 -595 6568 -593
rect 6577 -595 6798 -585
rect 6541 -605 6798 -595
rect 6827 -593 6877 -585
rect 6827 -602 6843 -593
rect 6436 -613 6487 -605
rect 6534 -613 6798 -605
rect 6824 -605 6843 -602
rect 6850 -605 6877 -593
rect 6824 -613 6877 -605
rect 6452 -621 6453 -613
rect 6468 -621 6481 -613
rect 6452 -629 6468 -621
rect 6449 -636 6468 -633
rect 6449 -645 6471 -636
rect 6422 -655 6471 -645
rect 6422 -661 6452 -655
rect 6471 -660 6476 -655
rect 6394 -677 6468 -661
rect 6486 -669 6516 -613
rect 6551 -623 6759 -613
rect 6794 -617 6839 -613
rect 6842 -614 6843 -613
rect 6858 -614 6871 -613
rect 6577 -653 6766 -623
rect 6592 -656 6766 -653
rect 6585 -659 6766 -656
rect 6394 -679 6407 -677
rect 6422 -679 6456 -677
rect 6394 -695 6468 -679
rect 6495 -683 6508 -669
rect 6523 -683 6539 -667
rect 6585 -672 6596 -659
rect 6378 -717 6379 -701
rect 6394 -717 6407 -695
rect 6422 -717 6452 -695
rect 6495 -699 6557 -683
rect 6585 -690 6596 -674
rect 6601 -679 6611 -659
rect 6621 -679 6635 -659
rect 6638 -672 6647 -659
rect 6663 -672 6672 -659
rect 6601 -690 6635 -679
rect 6638 -690 6647 -674
rect 6663 -690 6672 -674
rect 6679 -679 6689 -659
rect 6699 -679 6713 -659
rect 6714 -672 6725 -659
rect 6679 -690 6713 -679
rect 6714 -690 6725 -674
rect 6771 -683 6787 -667
rect 6794 -669 6824 -617
rect 6858 -621 6859 -614
rect 6843 -629 6859 -621
rect 6830 -661 6843 -642
rect 6858 -661 6888 -645
rect 6830 -677 6904 -661
rect 6830 -679 6843 -677
rect 6858 -679 6892 -677
rect 6495 -701 6508 -699
rect 6523 -701 6557 -699
rect 6495 -717 6557 -701
rect 6601 -706 6617 -703
rect 6679 -706 6709 -695
rect 6757 -699 6803 -683
rect 6830 -695 6904 -679
rect 6757 -701 6791 -699
rect 6756 -717 6803 -701
rect 6830 -717 6843 -695
rect 6858 -717 6888 -695
rect 6915 -717 6916 -701
rect 6931 -717 6944 -557
rect 4595 -750 4596 -724
rect 4603 -750 4630 -724
rect 4538 -768 4568 -754
rect 4595 -758 4630 -750
rect 4632 -725 4673 -717
rect 4632 -751 4647 -725
rect 4654 -751 4673 -725
rect 4737 -729 4799 -717
rect 4811 -729 4886 -717
rect 4944 -729 5019 -717
rect 5031 -729 5062 -717
rect 5068 -729 5103 -717
rect 4737 -731 4899 -729
rect 4595 -768 4596 -758
rect 4611 -768 4624 -758
rect 4632 -759 4673 -751
rect 4755 -755 4768 -731
rect 4783 -733 4798 -731
rect 4832 -749 4899 -731
rect 4931 -731 5103 -729
rect 4931 -749 5011 -731
rect 5032 -733 5047 -731
rect -2 -769 4624 -768
rect 4638 -769 4639 -759
rect 4654 -769 4667 -759
rect 4682 -769 4712 -755
rect 4755 -769 4798 -755
rect 4822 -758 4829 -751
rect 4832 -759 5011 -749
rect 4805 -769 4835 -759
rect 4837 -769 4990 -759
rect 4998 -769 5028 -759
rect 5032 -769 5062 -755
rect 5090 -769 5103 -731
rect 5175 -725 5210 -717
rect 5175 -751 5176 -725
rect 5183 -751 5210 -725
rect 5118 -769 5148 -755
rect 5175 -759 5210 -751
rect 5212 -725 5253 -717
rect 5212 -751 5227 -725
rect 5234 -751 5253 -725
rect 5317 -729 5379 -717
rect 5391 -729 5466 -717
rect 5524 -729 5599 -717
rect 5611 -729 5642 -717
rect 5648 -729 5683 -717
rect 5317 -731 5479 -729
rect 5212 -759 5253 -751
rect 5335 -755 5348 -731
rect 5363 -733 5378 -731
rect 5412 -749 5479 -731
rect 5511 -731 5683 -729
rect 5511 -749 5591 -731
rect 5612 -733 5627 -731
rect 5175 -769 5176 -759
rect 5191 -769 5204 -759
rect 5218 -769 5219 -759
rect 5234 -769 5247 -759
rect 5262 -769 5292 -755
rect 5335 -769 5378 -755
rect 5402 -758 5409 -751
rect 5412 -759 5591 -749
rect 5385 -769 5415 -759
rect 5417 -769 5570 -759
rect 5578 -769 5608 -759
rect 5612 -769 5642 -755
rect 5670 -769 5683 -731
rect 5755 -725 5790 -717
rect 5755 -751 5756 -725
rect 5763 -751 5790 -725
rect 5698 -769 5728 -755
rect 5755 -759 5790 -751
rect 5792 -725 5833 -717
rect 5792 -751 5807 -725
rect 5814 -751 5833 -725
rect 5897 -729 5959 -717
rect 5971 -729 6046 -717
rect 6104 -729 6179 -717
rect 6191 -729 6222 -717
rect 6228 -729 6263 -717
rect 5897 -731 6059 -729
rect 5792 -759 5833 -751
rect 5915 -755 5928 -731
rect 5943 -733 5958 -731
rect 5992 -749 6059 -731
rect 6091 -731 6263 -729
rect 6091 -749 6171 -731
rect 6192 -733 6207 -731
rect 5755 -769 5756 -759
rect 5771 -769 5784 -759
rect 5798 -769 5799 -759
rect 5814 -769 5827 -759
rect 5842 -769 5872 -755
rect 5915 -769 5958 -755
rect 5982 -758 5989 -751
rect 5992 -759 6171 -749
rect 5965 -769 5995 -759
rect 5997 -769 6150 -759
rect 6158 -769 6188 -759
rect 6192 -769 6222 -755
rect 6250 -769 6263 -731
rect 6335 -725 6370 -717
rect 6335 -751 6336 -725
rect 6343 -751 6370 -725
rect 6278 -769 6308 -755
rect 6335 -759 6370 -751
rect 6372 -725 6413 -717
rect 6372 -751 6387 -725
rect 6394 -751 6413 -725
rect 6477 -729 6539 -717
rect 6551 -729 6626 -717
rect 6684 -729 6759 -717
rect 6771 -729 6802 -717
rect 6808 -729 6843 -717
rect 6477 -731 6639 -729
rect 6372 -759 6413 -751
rect 6495 -755 6508 -731
rect 6523 -733 6538 -731
rect 6572 -749 6639 -731
rect 6671 -731 6843 -729
rect 6671 -749 6751 -731
rect 6772 -733 6787 -731
rect 6335 -769 6336 -759
rect 6351 -769 6364 -759
rect 6378 -769 6379 -759
rect 6394 -769 6407 -759
rect 6422 -769 6452 -755
rect 6495 -769 6538 -755
rect 6562 -758 6569 -751
rect 6572 -759 6751 -749
rect 6545 -769 6575 -759
rect 6577 -769 6730 -759
rect 6738 -769 6768 -759
rect 6772 -769 6802 -755
rect 6830 -769 6843 -731
rect 6915 -725 6950 -717
rect 6915 -751 6916 -725
rect 6923 -751 6950 -725
rect 6858 -769 6888 -755
rect 6915 -759 6950 -751
rect 6915 -769 6916 -759
rect 6931 -769 6944 -759
rect -2 -774 6944 -769
rect -1 -782 6944 -774
rect 14 -812 27 -782
rect 42 -800 72 -782
rect 115 -796 129 -782
rect 165 -796 385 -782
rect 116 -798 129 -796
rect 82 -810 97 -798
rect 79 -812 101 -810
rect 106 -812 136 -798
rect 197 -800 350 -796
rect 179 -812 371 -800
rect 414 -812 444 -798
rect 450 -812 463 -782
rect 478 -800 508 -782
rect 551 -812 564 -782
rect 594 -812 607 -782
rect 622 -800 652 -782
rect 695 -796 709 -782
rect 745 -796 965 -782
rect 696 -798 709 -796
rect 662 -810 677 -798
rect 659 -812 681 -810
rect 686 -812 716 -798
rect 777 -800 930 -796
rect 759 -812 951 -800
rect 994 -812 1024 -798
rect 1030 -812 1043 -782
rect 1058 -800 1088 -782
rect 1131 -812 1144 -782
rect 1174 -812 1187 -782
rect 1202 -800 1232 -782
rect 1275 -796 1289 -782
rect 1325 -796 1545 -782
rect 1276 -798 1289 -796
rect 1242 -810 1257 -798
rect 1239 -812 1261 -810
rect 1266 -812 1296 -798
rect 1357 -800 1510 -796
rect 1339 -812 1531 -800
rect 1574 -812 1604 -798
rect 1610 -812 1623 -782
rect 1638 -800 1668 -782
rect 1711 -812 1724 -782
rect 1754 -812 1767 -782
rect 1782 -800 1812 -782
rect 1855 -796 1869 -782
rect 1905 -796 2125 -782
rect 1856 -798 1869 -796
rect 1822 -810 1837 -798
rect 1819 -812 1841 -810
rect 1846 -812 1876 -798
rect 1937 -800 2090 -796
rect 1919 -812 2111 -800
rect 2154 -812 2184 -798
rect 2190 -812 2203 -782
rect 2218 -800 2248 -782
rect 2291 -812 2304 -782
rect 2334 -812 2347 -782
rect 2362 -800 2392 -782
rect 2435 -796 2449 -782
rect 2485 -796 2705 -782
rect 2436 -798 2449 -796
rect 2402 -810 2417 -798
rect 2399 -812 2421 -810
rect 2426 -812 2456 -798
rect 2517 -800 2670 -796
rect 2499 -812 2691 -800
rect 2734 -812 2764 -798
rect 2770 -812 2783 -782
rect 2798 -800 2828 -782
rect 2871 -812 2884 -782
rect 2914 -812 2927 -782
rect 2942 -800 2972 -782
rect 3015 -796 3029 -782
rect 3065 -796 3285 -782
rect 3016 -798 3029 -796
rect 2982 -810 2997 -798
rect 2979 -812 3001 -810
rect 3006 -812 3036 -798
rect 3097 -800 3250 -796
rect 3079 -812 3271 -800
rect 3314 -812 3344 -798
rect 3350 -812 3363 -782
rect 3378 -800 3408 -782
rect 3451 -812 3464 -782
rect 3494 -812 3507 -782
rect 3522 -800 3552 -782
rect 3595 -796 3609 -782
rect 3645 -796 3865 -782
rect 3596 -798 3609 -796
rect 3562 -810 3577 -798
rect 3559 -812 3581 -810
rect 3586 -812 3616 -798
rect 3677 -800 3830 -796
rect 3659 -812 3851 -800
rect 3894 -812 3924 -798
rect 3930 -812 3943 -782
rect 3958 -800 3988 -782
rect 4031 -812 4044 -782
rect 4074 -812 4087 -782
rect 4102 -800 4132 -782
rect 4175 -796 4189 -782
rect 4225 -796 4445 -782
rect 4176 -798 4189 -796
rect 4142 -810 4157 -798
rect 4139 -812 4161 -810
rect 4166 -812 4196 -798
rect 4257 -800 4410 -796
rect 4239 -812 4431 -800
rect 4474 -812 4504 -798
rect 4510 -812 4523 -782
rect 4538 -800 4568 -782
rect 4611 -783 6944 -782
rect 4611 -812 4624 -783
rect -1 -813 4624 -812
rect 4654 -813 4667 -783
rect 4682 -801 4712 -783
rect 4755 -797 4769 -783
rect 4805 -797 5025 -783
rect 4756 -799 4769 -797
rect 4722 -811 4737 -799
rect 4719 -813 4741 -811
rect 4746 -813 4776 -799
rect 4837 -801 4990 -797
rect 4819 -813 5011 -801
rect 5054 -813 5084 -799
rect 5090 -813 5103 -783
rect 5118 -801 5148 -783
rect 5191 -813 5204 -783
rect 5234 -813 5247 -783
rect 5262 -801 5292 -783
rect 5335 -797 5349 -783
rect 5385 -797 5605 -783
rect 5336 -799 5349 -797
rect 5302 -811 5317 -799
rect 5299 -813 5321 -811
rect 5326 -813 5356 -799
rect 5417 -801 5570 -797
rect 5399 -813 5591 -801
rect 5634 -813 5664 -799
rect 5670 -813 5683 -783
rect 5698 -801 5728 -783
rect 5771 -813 5784 -783
rect 5814 -813 5827 -783
rect 5842 -801 5872 -783
rect 5915 -797 5929 -783
rect 5965 -797 6185 -783
rect 5916 -799 5929 -797
rect 5882 -811 5897 -799
rect 5879 -813 5901 -811
rect 5906 -813 5936 -799
rect 5997 -801 6150 -797
rect 5979 -813 6171 -801
rect 6214 -813 6244 -799
rect 6250 -813 6263 -783
rect 6278 -801 6308 -783
rect 6351 -813 6364 -783
rect 6394 -813 6407 -783
rect 6422 -801 6452 -783
rect 6495 -797 6509 -783
rect 6545 -797 6765 -783
rect 6496 -799 6509 -797
rect 6462 -811 6477 -799
rect 6459 -813 6481 -811
rect 6486 -813 6516 -799
rect 6577 -801 6730 -797
rect 6559 -813 6751 -801
rect 6794 -813 6824 -799
rect 6830 -813 6843 -783
rect 6858 -801 6888 -783
rect 6931 -813 6944 -783
rect -1 -826 6944 -813
rect 14 -930 27 -826
rect 72 -848 73 -838
rect 88 -848 101 -838
rect 72 -852 101 -848
rect 106 -852 136 -826
rect 154 -840 170 -838
rect 242 -840 295 -826
rect 243 -842 307 -840
rect 350 -842 365 -826
rect 414 -829 444 -826
rect 414 -832 450 -829
rect 380 -840 396 -838
rect 154 -852 169 -848
rect 72 -854 169 -852
rect 197 -854 365 -842
rect 381 -852 396 -848
rect 414 -851 453 -832
rect 472 -838 479 -837
rect 478 -845 479 -838
rect 462 -848 463 -845
rect 478 -848 491 -845
rect 414 -852 444 -851
rect 453 -852 459 -851
rect 462 -852 491 -848
rect 381 -853 491 -852
rect 381 -854 497 -853
rect 56 -862 107 -854
rect 56 -874 81 -862
rect 88 -874 107 -862
rect 138 -862 188 -854
rect 138 -870 154 -862
rect 161 -864 188 -862
rect 197 -864 418 -854
rect 161 -874 418 -864
rect 447 -862 497 -854
rect 447 -871 463 -862
rect 56 -882 107 -874
rect 154 -882 418 -874
rect 444 -874 463 -871
rect 470 -874 497 -862
rect 444 -882 497 -874
rect 72 -890 73 -882
rect 88 -890 101 -882
rect 72 -898 88 -890
rect 69 -905 88 -902
rect 69 -914 91 -905
rect 42 -924 91 -914
rect 42 -930 72 -924
rect 91 -929 96 -924
rect 14 -946 88 -930
rect 106 -938 136 -882
rect 171 -892 379 -882
rect 414 -886 459 -882
rect 462 -883 463 -882
rect 478 -883 491 -882
rect 197 -922 386 -892
rect 212 -925 386 -922
rect 205 -928 386 -925
rect 14 -948 27 -946
rect 42 -948 76 -946
rect 14 -964 88 -948
rect 115 -952 128 -938
rect 143 -952 159 -936
rect 205 -941 216 -928
rect -2 -986 -1 -970
rect 14 -986 27 -964
rect 42 -986 72 -964
rect 115 -968 177 -952
rect 205 -959 216 -943
rect 221 -948 231 -928
rect 241 -948 255 -928
rect 258 -941 267 -928
rect 283 -941 292 -928
rect 221 -959 255 -948
rect 258 -959 267 -943
rect 283 -959 292 -943
rect 299 -948 309 -928
rect 319 -948 333 -928
rect 334 -941 345 -928
rect 299 -959 333 -948
rect 334 -959 345 -943
rect 391 -952 407 -936
rect 414 -938 444 -886
rect 478 -890 479 -883
rect 463 -898 479 -890
rect 450 -930 463 -911
rect 478 -930 508 -914
rect 450 -946 524 -930
rect 450 -948 463 -946
rect 478 -948 512 -946
rect 115 -970 128 -968
rect 143 -970 177 -968
rect 115 -986 177 -970
rect 221 -975 237 -972
rect 299 -975 329 -964
rect 377 -968 423 -952
rect 450 -964 524 -948
rect 377 -970 411 -968
rect 376 -986 423 -970
rect 450 -986 463 -964
rect 478 -986 508 -964
rect 535 -986 536 -970
rect 551 -986 564 -826
rect 594 -930 607 -826
rect 652 -848 653 -838
rect 668 -848 681 -838
rect 652 -852 681 -848
rect 686 -852 716 -826
rect 734 -840 750 -838
rect 822 -840 875 -826
rect 823 -842 887 -840
rect 930 -842 945 -826
rect 994 -829 1024 -826
rect 994 -832 1030 -829
rect 960 -840 976 -838
rect 734 -852 749 -848
rect 652 -854 749 -852
rect 777 -854 945 -842
rect 961 -852 976 -848
rect 994 -851 1033 -832
rect 1052 -838 1059 -837
rect 1058 -845 1059 -838
rect 1042 -848 1043 -845
rect 1058 -848 1071 -845
rect 994 -852 1024 -851
rect 1033 -852 1039 -851
rect 1042 -852 1071 -848
rect 961 -853 1071 -852
rect 961 -854 1077 -853
rect 636 -862 687 -854
rect 636 -874 661 -862
rect 668 -874 687 -862
rect 718 -862 768 -854
rect 718 -870 734 -862
rect 741 -864 768 -862
rect 777 -864 998 -854
rect 741 -874 998 -864
rect 1027 -862 1077 -854
rect 1027 -871 1043 -862
rect 636 -882 687 -874
rect 734 -882 998 -874
rect 1024 -874 1043 -871
rect 1050 -874 1077 -862
rect 1024 -882 1077 -874
rect 652 -890 653 -882
rect 668 -890 681 -882
rect 652 -898 668 -890
rect 649 -905 668 -902
rect 649 -914 671 -905
rect 622 -924 671 -914
rect 622 -930 652 -924
rect 671 -929 676 -924
rect 594 -946 668 -930
rect 686 -938 716 -882
rect 751 -892 959 -882
rect 994 -886 1039 -882
rect 1042 -883 1043 -882
rect 1058 -883 1071 -882
rect 777 -922 966 -892
rect 792 -925 966 -922
rect 785 -928 966 -925
rect 594 -948 607 -946
rect 622 -948 656 -946
rect 594 -964 668 -948
rect 695 -952 708 -938
rect 723 -952 739 -936
rect 785 -941 796 -928
rect 578 -986 579 -970
rect 594 -986 607 -964
rect 622 -986 652 -964
rect 695 -968 757 -952
rect 785 -959 796 -943
rect 801 -948 811 -928
rect 821 -948 835 -928
rect 838 -941 847 -928
rect 863 -941 872 -928
rect 801 -959 835 -948
rect 838 -959 847 -943
rect 863 -959 872 -943
rect 879 -948 889 -928
rect 899 -948 913 -928
rect 914 -941 925 -928
rect 879 -959 913 -948
rect 914 -959 925 -943
rect 971 -952 987 -936
rect 994 -938 1024 -886
rect 1058 -890 1059 -883
rect 1043 -898 1059 -890
rect 1030 -930 1043 -911
rect 1058 -930 1088 -914
rect 1030 -946 1104 -930
rect 1030 -948 1043 -946
rect 1058 -948 1092 -946
rect 695 -970 708 -968
rect 723 -970 757 -968
rect 695 -986 757 -970
rect 801 -975 817 -972
rect 879 -975 909 -964
rect 957 -968 1003 -952
rect 1030 -964 1104 -948
rect 957 -970 991 -968
rect 956 -986 1003 -970
rect 1030 -986 1043 -964
rect 1058 -986 1088 -964
rect 1115 -986 1116 -970
rect 1131 -986 1144 -826
rect 1174 -930 1187 -826
rect 1232 -848 1233 -838
rect 1248 -848 1261 -838
rect 1232 -852 1261 -848
rect 1266 -852 1296 -826
rect 1314 -840 1330 -838
rect 1402 -840 1455 -826
rect 1403 -842 1467 -840
rect 1510 -842 1525 -826
rect 1574 -829 1604 -826
rect 1574 -832 1610 -829
rect 1540 -840 1556 -838
rect 1314 -852 1329 -848
rect 1232 -854 1329 -852
rect 1357 -854 1525 -842
rect 1541 -852 1556 -848
rect 1574 -851 1613 -832
rect 1632 -838 1639 -837
rect 1638 -845 1639 -838
rect 1622 -848 1623 -845
rect 1638 -848 1651 -845
rect 1574 -852 1604 -851
rect 1613 -852 1619 -851
rect 1622 -852 1651 -848
rect 1541 -853 1651 -852
rect 1541 -854 1657 -853
rect 1216 -862 1267 -854
rect 1216 -874 1241 -862
rect 1248 -874 1267 -862
rect 1298 -862 1348 -854
rect 1298 -870 1314 -862
rect 1321 -864 1348 -862
rect 1357 -864 1578 -854
rect 1321 -874 1578 -864
rect 1607 -862 1657 -854
rect 1607 -871 1623 -862
rect 1216 -882 1267 -874
rect 1314 -882 1578 -874
rect 1604 -874 1623 -871
rect 1630 -874 1657 -862
rect 1604 -882 1657 -874
rect 1232 -890 1233 -882
rect 1248 -890 1261 -882
rect 1232 -898 1248 -890
rect 1229 -905 1248 -902
rect 1229 -914 1251 -905
rect 1202 -924 1251 -914
rect 1202 -930 1232 -924
rect 1251 -929 1256 -924
rect 1174 -946 1248 -930
rect 1266 -938 1296 -882
rect 1331 -892 1539 -882
rect 1574 -886 1619 -882
rect 1622 -883 1623 -882
rect 1638 -883 1651 -882
rect 1357 -922 1546 -892
rect 1372 -925 1546 -922
rect 1365 -928 1546 -925
rect 1174 -948 1187 -946
rect 1202 -948 1236 -946
rect 1174 -964 1248 -948
rect 1275 -952 1288 -938
rect 1303 -952 1319 -936
rect 1365 -941 1376 -928
rect 1158 -986 1159 -970
rect 1174 -986 1187 -964
rect 1202 -986 1232 -964
rect 1275 -968 1337 -952
rect 1365 -959 1376 -943
rect 1381 -948 1391 -928
rect 1401 -948 1415 -928
rect 1418 -941 1427 -928
rect 1443 -941 1452 -928
rect 1381 -959 1415 -948
rect 1418 -959 1427 -943
rect 1443 -959 1452 -943
rect 1459 -948 1469 -928
rect 1479 -948 1493 -928
rect 1494 -941 1505 -928
rect 1459 -959 1493 -948
rect 1494 -959 1505 -943
rect 1551 -952 1567 -936
rect 1574 -938 1604 -886
rect 1638 -890 1639 -883
rect 1623 -898 1639 -890
rect 1610 -930 1623 -911
rect 1638 -930 1668 -914
rect 1610 -946 1684 -930
rect 1610 -948 1623 -946
rect 1638 -948 1672 -946
rect 1275 -970 1288 -968
rect 1303 -970 1337 -968
rect 1275 -986 1337 -970
rect 1381 -975 1397 -972
rect 1459 -975 1489 -964
rect 1537 -968 1583 -952
rect 1610 -964 1684 -948
rect 1537 -970 1571 -968
rect 1536 -986 1583 -970
rect 1610 -986 1623 -964
rect 1638 -986 1668 -964
rect 1695 -986 1696 -970
rect 1711 -986 1724 -826
rect 1754 -930 1767 -826
rect 1812 -848 1813 -838
rect 1828 -848 1841 -838
rect 1812 -852 1841 -848
rect 1846 -852 1876 -826
rect 1894 -840 1910 -838
rect 1982 -840 2035 -826
rect 1983 -842 2047 -840
rect 2090 -842 2105 -826
rect 2154 -829 2184 -826
rect 2154 -832 2190 -829
rect 2120 -840 2136 -838
rect 1894 -852 1909 -848
rect 1812 -854 1909 -852
rect 1937 -854 2105 -842
rect 2121 -852 2136 -848
rect 2154 -851 2193 -832
rect 2212 -838 2219 -837
rect 2218 -845 2219 -838
rect 2202 -848 2203 -845
rect 2218 -848 2231 -845
rect 2154 -852 2184 -851
rect 2193 -852 2199 -851
rect 2202 -852 2231 -848
rect 2121 -853 2231 -852
rect 2121 -854 2237 -853
rect 1796 -862 1847 -854
rect 1796 -874 1821 -862
rect 1828 -874 1847 -862
rect 1878 -862 1928 -854
rect 1878 -870 1894 -862
rect 1901 -864 1928 -862
rect 1937 -864 2158 -854
rect 1901 -874 2158 -864
rect 2187 -862 2237 -854
rect 2187 -871 2203 -862
rect 1796 -882 1847 -874
rect 1894 -882 2158 -874
rect 2184 -874 2203 -871
rect 2210 -874 2237 -862
rect 2184 -882 2237 -874
rect 1812 -890 1813 -882
rect 1828 -890 1841 -882
rect 1812 -898 1828 -890
rect 1809 -905 1828 -902
rect 1809 -914 1831 -905
rect 1782 -924 1831 -914
rect 1782 -930 1812 -924
rect 1831 -929 1836 -924
rect 1754 -946 1828 -930
rect 1846 -938 1876 -882
rect 1911 -892 2119 -882
rect 2154 -886 2199 -882
rect 2202 -883 2203 -882
rect 2218 -883 2231 -882
rect 1937 -922 2126 -892
rect 1952 -925 2126 -922
rect 1945 -928 2126 -925
rect 1754 -948 1767 -946
rect 1782 -948 1816 -946
rect 1754 -964 1828 -948
rect 1855 -952 1868 -938
rect 1883 -952 1899 -936
rect 1945 -941 1956 -928
rect 1738 -986 1739 -970
rect 1754 -986 1767 -964
rect 1782 -986 1812 -964
rect 1855 -968 1917 -952
rect 1945 -959 1956 -943
rect 1961 -948 1971 -928
rect 1981 -948 1995 -928
rect 1998 -941 2007 -928
rect 2023 -941 2032 -928
rect 1961 -959 1995 -948
rect 1998 -959 2007 -943
rect 2023 -959 2032 -943
rect 2039 -948 2049 -928
rect 2059 -948 2073 -928
rect 2074 -941 2085 -928
rect 2039 -959 2073 -948
rect 2074 -959 2085 -943
rect 2131 -952 2147 -936
rect 2154 -938 2184 -886
rect 2218 -890 2219 -883
rect 2203 -898 2219 -890
rect 2190 -930 2203 -911
rect 2218 -930 2248 -914
rect 2190 -946 2264 -930
rect 2190 -948 2203 -946
rect 2218 -948 2252 -946
rect 1855 -970 1868 -968
rect 1883 -970 1917 -968
rect 1855 -986 1917 -970
rect 1961 -975 1977 -972
rect 2039 -975 2069 -964
rect 2117 -968 2163 -952
rect 2190 -964 2264 -948
rect 2117 -970 2151 -968
rect 2116 -986 2163 -970
rect 2190 -986 2203 -964
rect 2218 -986 2248 -964
rect 2275 -986 2276 -970
rect 2291 -986 2304 -826
rect 2334 -930 2347 -826
rect 2392 -848 2393 -838
rect 2408 -848 2421 -838
rect 2392 -852 2421 -848
rect 2426 -852 2456 -826
rect 2474 -840 2490 -838
rect 2562 -840 2615 -826
rect 2563 -842 2627 -840
rect 2670 -842 2685 -826
rect 2734 -829 2764 -826
rect 2734 -832 2770 -829
rect 2700 -840 2716 -838
rect 2474 -852 2489 -848
rect 2392 -854 2489 -852
rect 2517 -854 2685 -842
rect 2701 -852 2716 -848
rect 2734 -851 2773 -832
rect 2792 -838 2799 -837
rect 2798 -845 2799 -838
rect 2782 -848 2783 -845
rect 2798 -848 2811 -845
rect 2734 -852 2764 -851
rect 2773 -852 2779 -851
rect 2782 -852 2811 -848
rect 2701 -853 2811 -852
rect 2701 -854 2817 -853
rect 2376 -862 2427 -854
rect 2376 -874 2401 -862
rect 2408 -874 2427 -862
rect 2458 -862 2508 -854
rect 2458 -870 2474 -862
rect 2481 -864 2508 -862
rect 2517 -864 2738 -854
rect 2481 -874 2738 -864
rect 2767 -862 2817 -854
rect 2767 -871 2783 -862
rect 2376 -882 2427 -874
rect 2474 -882 2738 -874
rect 2764 -874 2783 -871
rect 2790 -874 2817 -862
rect 2764 -882 2817 -874
rect 2392 -890 2393 -882
rect 2408 -890 2421 -882
rect 2392 -898 2408 -890
rect 2389 -905 2408 -902
rect 2389 -914 2411 -905
rect 2362 -924 2411 -914
rect 2362 -930 2392 -924
rect 2411 -929 2416 -924
rect 2334 -946 2408 -930
rect 2426 -938 2456 -882
rect 2491 -892 2699 -882
rect 2734 -886 2779 -882
rect 2782 -883 2783 -882
rect 2798 -883 2811 -882
rect 2517 -922 2706 -892
rect 2532 -925 2706 -922
rect 2525 -928 2706 -925
rect 2334 -948 2347 -946
rect 2362 -948 2396 -946
rect 2334 -964 2408 -948
rect 2435 -952 2448 -938
rect 2463 -952 2479 -936
rect 2525 -941 2536 -928
rect 2318 -986 2319 -970
rect 2334 -986 2347 -964
rect 2362 -986 2392 -964
rect 2435 -968 2497 -952
rect 2525 -959 2536 -943
rect 2541 -948 2551 -928
rect 2561 -948 2575 -928
rect 2578 -941 2587 -928
rect 2603 -941 2612 -928
rect 2541 -959 2575 -948
rect 2578 -959 2587 -943
rect 2603 -959 2612 -943
rect 2619 -948 2629 -928
rect 2639 -948 2653 -928
rect 2654 -941 2665 -928
rect 2619 -959 2653 -948
rect 2654 -959 2665 -943
rect 2711 -952 2727 -936
rect 2734 -938 2764 -886
rect 2798 -890 2799 -883
rect 2783 -898 2799 -890
rect 2770 -930 2783 -911
rect 2798 -930 2828 -914
rect 2770 -946 2844 -930
rect 2770 -948 2783 -946
rect 2798 -948 2832 -946
rect 2435 -970 2448 -968
rect 2463 -970 2497 -968
rect 2435 -986 2497 -970
rect 2541 -975 2557 -972
rect 2619 -975 2649 -964
rect 2697 -968 2743 -952
rect 2770 -964 2844 -948
rect 2697 -970 2731 -968
rect 2696 -986 2743 -970
rect 2770 -986 2783 -964
rect 2798 -986 2828 -964
rect 2855 -986 2856 -970
rect 2871 -986 2884 -826
rect 2914 -930 2927 -826
rect 2972 -848 2973 -838
rect 2988 -848 3001 -838
rect 2972 -852 3001 -848
rect 3006 -852 3036 -826
rect 3054 -840 3070 -838
rect 3142 -840 3195 -826
rect 3143 -842 3205 -840
rect 3250 -842 3265 -826
rect 3314 -829 3344 -826
rect 3314 -832 3350 -829
rect 3280 -840 3296 -838
rect 3054 -852 3069 -848
rect 2972 -854 3069 -852
rect 3097 -854 3265 -842
rect 3281 -852 3296 -848
rect 3314 -851 3353 -832
rect 3372 -838 3379 -837
rect 3378 -845 3379 -838
rect 3362 -848 3363 -845
rect 3378 -848 3391 -845
rect 3314 -852 3344 -851
rect 3353 -852 3359 -851
rect 3362 -852 3391 -848
rect 3281 -853 3391 -852
rect 3281 -854 3397 -853
rect 2956 -862 3007 -854
rect 2956 -874 2981 -862
rect 2988 -874 3007 -862
rect 3038 -862 3088 -854
rect 3038 -870 3054 -862
rect 3061 -864 3088 -862
rect 3097 -864 3318 -854
rect 3061 -874 3318 -864
rect 3347 -862 3397 -854
rect 3347 -871 3363 -862
rect 2956 -882 3007 -874
rect 3054 -882 3318 -874
rect 3344 -874 3363 -871
rect 3370 -874 3397 -862
rect 3344 -882 3397 -874
rect 2972 -890 2973 -882
rect 2988 -890 3001 -882
rect 2972 -898 2988 -890
rect 2969 -905 2988 -902
rect 2969 -914 2991 -905
rect 2942 -924 2991 -914
rect 2942 -930 2972 -924
rect 2991 -929 2996 -924
rect 2914 -946 2988 -930
rect 3006 -938 3036 -882
rect 3071 -892 3279 -882
rect 3314 -886 3359 -882
rect 3362 -883 3363 -882
rect 3378 -883 3391 -882
rect 3097 -922 3286 -892
rect 3112 -925 3286 -922
rect 3105 -928 3286 -925
rect 2914 -948 2927 -946
rect 2942 -948 2976 -946
rect 2914 -964 2988 -948
rect 3015 -952 3028 -938
rect 3043 -952 3059 -936
rect 3105 -941 3116 -928
rect 2898 -986 2899 -970
rect 2914 -986 2927 -964
rect 2942 -986 2972 -964
rect 3015 -968 3077 -952
rect 3105 -959 3116 -943
rect 3121 -948 3131 -928
rect 3141 -948 3155 -928
rect 3158 -941 3167 -928
rect 3183 -941 3192 -928
rect 3121 -959 3155 -948
rect 3158 -959 3167 -943
rect 3183 -959 3192 -943
rect 3199 -948 3209 -928
rect 3219 -948 3233 -928
rect 3234 -941 3245 -928
rect 3199 -959 3233 -948
rect 3234 -959 3245 -943
rect 3291 -952 3307 -936
rect 3314 -938 3344 -886
rect 3378 -890 3379 -883
rect 3363 -898 3379 -890
rect 3350 -930 3363 -911
rect 3378 -930 3408 -914
rect 3350 -946 3424 -930
rect 3350 -948 3363 -946
rect 3378 -948 3412 -946
rect 3015 -970 3028 -968
rect 3043 -970 3077 -968
rect 3015 -986 3077 -970
rect 3121 -975 3137 -972
rect 3199 -975 3229 -964
rect 3277 -968 3323 -952
rect 3350 -964 3424 -948
rect 3277 -970 3311 -968
rect 3276 -986 3323 -970
rect 3350 -986 3363 -964
rect 3378 -986 3408 -964
rect 3435 -986 3436 -970
rect 3451 -986 3464 -826
rect 3494 -930 3507 -826
rect 3552 -848 3553 -838
rect 3568 -848 3581 -838
rect 3552 -852 3581 -848
rect 3586 -852 3616 -826
rect 3634 -840 3650 -838
rect 3722 -840 3775 -826
rect 3723 -842 3787 -840
rect 3830 -842 3845 -826
rect 3894 -829 3924 -826
rect 3894 -832 3930 -829
rect 3860 -840 3876 -838
rect 3634 -852 3649 -848
rect 3552 -854 3649 -852
rect 3677 -854 3845 -842
rect 3861 -852 3876 -848
rect 3894 -851 3933 -832
rect 3952 -838 3959 -837
rect 3958 -845 3959 -838
rect 3942 -848 3943 -845
rect 3958 -848 3971 -845
rect 3894 -852 3924 -851
rect 3933 -852 3939 -851
rect 3942 -852 3971 -848
rect 3861 -853 3971 -852
rect 3861 -854 3977 -853
rect 3536 -862 3587 -854
rect 3536 -874 3561 -862
rect 3568 -874 3587 -862
rect 3618 -862 3668 -854
rect 3618 -870 3634 -862
rect 3641 -864 3668 -862
rect 3677 -864 3898 -854
rect 3641 -874 3898 -864
rect 3927 -862 3977 -854
rect 3927 -871 3943 -862
rect 3536 -882 3587 -874
rect 3634 -882 3898 -874
rect 3924 -874 3943 -871
rect 3950 -874 3977 -862
rect 3924 -882 3977 -874
rect 3552 -890 3553 -882
rect 3568 -890 3581 -882
rect 3552 -898 3568 -890
rect 3549 -905 3568 -902
rect 3549 -914 3571 -905
rect 3522 -924 3571 -914
rect 3522 -930 3552 -924
rect 3571 -929 3576 -924
rect 3494 -946 3568 -930
rect 3586 -938 3616 -882
rect 3651 -892 3859 -882
rect 3894 -886 3939 -882
rect 3942 -883 3943 -882
rect 3958 -883 3971 -882
rect 3677 -922 3866 -892
rect 3692 -925 3866 -922
rect 3685 -928 3866 -925
rect 3494 -948 3507 -946
rect 3522 -948 3556 -946
rect 3494 -964 3568 -948
rect 3595 -952 3608 -938
rect 3623 -952 3639 -936
rect 3685 -941 3696 -928
rect 3478 -986 3479 -970
rect 3494 -986 3507 -964
rect 3522 -986 3552 -964
rect 3595 -968 3657 -952
rect 3685 -959 3696 -943
rect 3701 -948 3711 -928
rect 3721 -948 3735 -928
rect 3738 -941 3747 -928
rect 3763 -941 3772 -928
rect 3701 -959 3735 -948
rect 3738 -959 3747 -943
rect 3763 -959 3772 -943
rect 3779 -948 3789 -928
rect 3799 -948 3813 -928
rect 3814 -941 3825 -928
rect 3779 -959 3813 -948
rect 3814 -959 3825 -943
rect 3871 -952 3887 -936
rect 3894 -938 3924 -886
rect 3958 -890 3959 -883
rect 3943 -898 3959 -890
rect 3930 -930 3943 -911
rect 3958 -930 3988 -914
rect 3930 -946 4004 -930
rect 3930 -948 3943 -946
rect 3958 -948 3992 -946
rect 3595 -970 3608 -968
rect 3623 -970 3657 -968
rect 3595 -986 3657 -970
rect 3701 -975 3717 -972
rect 3779 -975 3809 -964
rect 3857 -968 3903 -952
rect 3930 -964 4004 -948
rect 3857 -970 3891 -968
rect 3856 -986 3903 -970
rect 3930 -986 3943 -964
rect 3958 -986 3988 -964
rect 4015 -986 4016 -970
rect 4031 -986 4044 -826
rect 4074 -930 4087 -826
rect 4132 -848 4133 -838
rect 4148 -848 4161 -838
rect 4132 -852 4161 -848
rect 4166 -852 4196 -826
rect 4214 -840 4230 -838
rect 4302 -840 4355 -826
rect 4303 -842 4367 -840
rect 4410 -842 4425 -826
rect 4474 -829 4504 -826
rect 4611 -827 6944 -826
rect 4474 -832 4510 -829
rect 4440 -840 4456 -838
rect 4214 -852 4229 -848
rect 4132 -854 4229 -852
rect 4257 -854 4425 -842
rect 4441 -852 4456 -848
rect 4474 -851 4513 -832
rect 4532 -838 4539 -837
rect 4538 -845 4539 -838
rect 4522 -848 4523 -845
rect 4538 -848 4551 -845
rect 4474 -852 4504 -851
rect 4513 -852 4519 -851
rect 4522 -852 4551 -848
rect 4441 -853 4551 -852
rect 4441 -854 4557 -853
rect 4116 -862 4167 -854
rect 4116 -874 4141 -862
rect 4148 -874 4167 -862
rect 4198 -862 4248 -854
rect 4198 -870 4214 -862
rect 4221 -864 4248 -862
rect 4257 -864 4478 -854
rect 4221 -874 4478 -864
rect 4507 -862 4557 -854
rect 4507 -871 4523 -862
rect 4116 -882 4167 -874
rect 4214 -882 4478 -874
rect 4504 -874 4523 -871
rect 4530 -874 4557 -862
rect 4504 -882 4557 -874
rect 4132 -890 4133 -882
rect 4148 -890 4161 -882
rect 4132 -898 4148 -890
rect 4129 -905 4148 -902
rect 4129 -914 4151 -905
rect 4102 -924 4151 -914
rect 4102 -930 4132 -924
rect 4151 -929 4156 -924
rect 4074 -946 4148 -930
rect 4166 -938 4196 -882
rect 4231 -892 4439 -882
rect 4474 -886 4519 -882
rect 4522 -883 4523 -882
rect 4538 -883 4551 -882
rect 4257 -922 4446 -892
rect 4272 -925 4446 -922
rect 4265 -928 4446 -925
rect 4074 -948 4087 -946
rect 4102 -948 4136 -946
rect 4074 -964 4148 -948
rect 4175 -952 4188 -938
rect 4203 -952 4219 -936
rect 4265 -941 4276 -928
rect 4058 -986 4059 -970
rect 4074 -986 4087 -964
rect 4102 -986 4132 -964
rect 4175 -968 4237 -952
rect 4265 -959 4276 -943
rect 4281 -948 4291 -928
rect 4301 -948 4315 -928
rect 4318 -941 4327 -928
rect 4343 -941 4352 -928
rect 4281 -959 4315 -948
rect 4318 -959 4327 -943
rect 4343 -959 4352 -943
rect 4359 -948 4369 -928
rect 4379 -948 4393 -928
rect 4394 -941 4405 -928
rect 4359 -959 4393 -948
rect 4394 -959 4405 -943
rect 4451 -952 4467 -936
rect 4474 -938 4504 -886
rect 4538 -890 4539 -883
rect 4523 -898 4539 -890
rect 4510 -930 4523 -911
rect 4538 -930 4568 -914
rect 4510 -946 4584 -930
rect 4510 -948 4523 -946
rect 4538 -948 4572 -946
rect 4175 -970 4188 -968
rect 4203 -970 4237 -968
rect 4175 -986 4237 -970
rect 4281 -975 4297 -972
rect 4359 -975 4389 -964
rect 4437 -968 4483 -952
rect 4510 -964 4584 -948
rect 4437 -970 4471 -968
rect 4436 -986 4483 -970
rect 4510 -986 4523 -964
rect 4538 -986 4568 -964
rect 4595 -986 4596 -970
rect 4611 -986 4624 -827
rect 4654 -931 4667 -827
rect 4712 -849 4713 -839
rect 4733 -841 4741 -839
rect 4731 -843 4741 -841
rect 4728 -849 4741 -843
rect 4712 -853 4741 -849
rect 4746 -853 4776 -827
rect 4794 -841 4810 -839
rect 4882 -841 4933 -827
rect 4883 -843 4947 -841
rect 4990 -843 5005 -827
rect 5054 -830 5084 -827
rect 5054 -833 5090 -830
rect 5020 -841 5036 -839
rect 4794 -853 4809 -849
rect 4712 -855 4809 -853
rect 4837 -855 5005 -843
rect 5021 -853 5036 -849
rect 5054 -852 5093 -833
rect 5112 -839 5119 -838
rect 5118 -846 5119 -839
rect 5102 -849 5103 -846
rect 5118 -849 5131 -846
rect 5054 -853 5084 -852
rect 5093 -853 5099 -852
rect 5102 -853 5131 -849
rect 5021 -854 5131 -853
rect 5021 -855 5137 -854
rect 4696 -863 4747 -855
rect 4696 -875 4721 -863
rect 4728 -875 4747 -863
rect 4778 -863 4828 -855
rect 4778 -871 4794 -863
rect 4801 -865 4828 -863
rect 4837 -865 5058 -855
rect 4801 -875 5058 -865
rect 5087 -863 5137 -855
rect 5087 -872 5103 -863
rect 4696 -883 4747 -875
rect 4794 -883 5058 -875
rect 5084 -875 5103 -872
rect 5110 -875 5137 -863
rect 5084 -883 5137 -875
rect 4712 -891 4713 -883
rect 4728 -891 4741 -883
rect 4712 -899 4728 -891
rect 4709 -906 4728 -903
rect 4709 -915 4731 -906
rect 4682 -925 4731 -915
rect 4682 -931 4712 -925
rect 4731 -930 4736 -925
rect 4654 -947 4728 -931
rect 4746 -939 4776 -883
rect 4811 -893 5019 -883
rect 5054 -887 5099 -883
rect 5102 -884 5103 -883
rect 5118 -884 5131 -883
rect 4837 -923 5026 -893
rect 4852 -926 5026 -923
rect 4845 -929 5026 -926
rect 4654 -949 4667 -947
rect 4682 -949 4716 -947
rect 4654 -965 4728 -949
rect 4755 -953 4768 -939
rect 4783 -953 4799 -937
rect 4845 -942 4856 -929
rect -8 -994 33 -986
rect -8 -1020 7 -994
rect 14 -1020 33 -994
rect 97 -998 159 -986
rect 171 -998 246 -986
rect 304 -998 379 -986
rect 391 -998 422 -986
rect 428 -998 463 -986
rect 97 -1000 259 -998
rect -8 -1028 33 -1020
rect 115 -1024 128 -1000
rect 143 -1002 158 -1000
rect -2 -1038 -1 -1028
rect 14 -1038 27 -1028
rect 42 -1038 72 -1024
rect 115 -1038 158 -1024
rect 182 -1027 189 -1020
rect 192 -1024 259 -1000
rect 291 -1000 463 -998
rect 261 -1022 289 -1018
rect 291 -1022 371 -1000
rect 392 -1002 407 -1000
rect 261 -1024 371 -1022
rect 192 -1028 371 -1024
rect 165 -1038 195 -1028
rect 197 -1038 350 -1028
rect 358 -1038 388 -1028
rect 392 -1038 422 -1024
rect 450 -1038 463 -1000
rect 535 -994 570 -986
rect 535 -1020 536 -994
rect 543 -1020 570 -994
rect 478 -1038 508 -1024
rect 535 -1028 570 -1020
rect 572 -994 613 -986
rect 572 -1020 587 -994
rect 594 -1020 613 -994
rect 677 -998 739 -986
rect 751 -998 826 -986
rect 884 -998 959 -986
rect 971 -998 1002 -986
rect 1008 -998 1043 -986
rect 677 -1000 839 -998
rect 572 -1028 613 -1020
rect 695 -1024 708 -1000
rect 723 -1002 738 -1000
rect 535 -1038 536 -1028
rect 551 -1038 564 -1028
rect 578 -1038 579 -1028
rect 594 -1038 607 -1028
rect 622 -1038 652 -1024
rect 695 -1038 738 -1024
rect 762 -1027 769 -1020
rect 772 -1024 839 -1000
rect 871 -1000 1043 -998
rect 841 -1022 869 -1018
rect 871 -1022 951 -1000
rect 972 -1002 987 -1000
rect 841 -1024 951 -1022
rect 772 -1028 951 -1024
rect 745 -1038 775 -1028
rect 777 -1038 930 -1028
rect 938 -1038 968 -1028
rect 972 -1038 1002 -1024
rect 1030 -1038 1043 -1000
rect 1115 -994 1150 -986
rect 1115 -1020 1116 -994
rect 1123 -1020 1150 -994
rect 1058 -1038 1088 -1024
rect 1115 -1028 1150 -1020
rect 1152 -994 1193 -986
rect 1152 -1020 1167 -994
rect 1174 -1020 1193 -994
rect 1257 -998 1319 -986
rect 1331 -998 1406 -986
rect 1464 -998 1539 -986
rect 1551 -998 1582 -986
rect 1588 -998 1623 -986
rect 1257 -1000 1419 -998
rect 1152 -1028 1193 -1020
rect 1275 -1024 1288 -1000
rect 1303 -1002 1318 -1000
rect 1115 -1038 1116 -1028
rect 1131 -1038 1144 -1028
rect 1158 -1038 1159 -1028
rect 1174 -1038 1187 -1028
rect 1202 -1038 1232 -1024
rect 1275 -1038 1318 -1024
rect 1342 -1027 1349 -1020
rect 1352 -1024 1419 -1000
rect 1451 -1000 1623 -998
rect 1421 -1022 1449 -1018
rect 1451 -1022 1531 -1000
rect 1552 -1002 1567 -1000
rect 1421 -1024 1531 -1022
rect 1352 -1028 1531 -1024
rect 1325 -1038 1355 -1028
rect 1357 -1038 1510 -1028
rect 1518 -1038 1548 -1028
rect 1552 -1038 1582 -1024
rect 1610 -1038 1623 -1000
rect 1695 -994 1730 -986
rect 1695 -1020 1696 -994
rect 1703 -1020 1730 -994
rect 1638 -1038 1668 -1024
rect 1695 -1028 1730 -1020
rect 1732 -994 1773 -986
rect 1732 -1020 1747 -994
rect 1754 -1020 1773 -994
rect 1837 -998 1899 -986
rect 1911 -998 1986 -986
rect 2044 -998 2119 -986
rect 2131 -998 2162 -986
rect 2168 -998 2203 -986
rect 1837 -1000 1999 -998
rect 1732 -1028 1773 -1020
rect 1855 -1024 1868 -1000
rect 1883 -1002 1898 -1000
rect 1695 -1038 1696 -1028
rect 1711 -1038 1724 -1028
rect 1738 -1038 1739 -1028
rect 1754 -1038 1767 -1028
rect 1782 -1038 1812 -1024
rect 1855 -1038 1898 -1024
rect 1922 -1027 1929 -1020
rect 1932 -1024 1999 -1000
rect 2031 -1000 2203 -998
rect 2001 -1022 2029 -1018
rect 2031 -1022 2111 -1000
rect 2132 -1002 2147 -1000
rect 2001 -1024 2111 -1022
rect 1932 -1028 2111 -1024
rect 1905 -1038 1935 -1028
rect 1937 -1038 2090 -1028
rect 2098 -1038 2128 -1028
rect 2132 -1038 2162 -1024
rect 2190 -1038 2203 -1000
rect 2275 -994 2310 -986
rect 2275 -1020 2276 -994
rect 2283 -1020 2310 -994
rect 2218 -1038 2248 -1024
rect 2275 -1028 2310 -1020
rect 2312 -994 2353 -986
rect 2312 -1020 2327 -994
rect 2334 -1020 2353 -994
rect 2417 -998 2479 -986
rect 2491 -998 2566 -986
rect 2624 -998 2699 -986
rect 2711 -998 2742 -986
rect 2748 -998 2783 -986
rect 2417 -1000 2579 -998
rect 2312 -1028 2353 -1020
rect 2435 -1024 2448 -1000
rect 2463 -1002 2478 -1000
rect 2275 -1038 2276 -1028
rect 2291 -1038 2304 -1028
rect 2318 -1038 2319 -1028
rect 2334 -1038 2347 -1028
rect 2362 -1038 2392 -1024
rect 2435 -1038 2478 -1024
rect 2502 -1027 2509 -1020
rect 2512 -1024 2579 -1000
rect 2611 -1000 2783 -998
rect 2581 -1022 2609 -1018
rect 2611 -1022 2691 -1000
rect 2712 -1002 2727 -1000
rect 2581 -1024 2691 -1022
rect 2512 -1028 2691 -1024
rect 2485 -1038 2515 -1028
rect 2517 -1038 2670 -1028
rect 2678 -1038 2708 -1028
rect 2712 -1038 2742 -1024
rect 2770 -1038 2783 -1000
rect 2855 -994 2890 -986
rect 2855 -1020 2856 -994
rect 2863 -1020 2890 -994
rect 2798 -1038 2828 -1024
rect 2855 -1028 2890 -1020
rect 2892 -994 2933 -986
rect 2892 -1020 2907 -994
rect 2914 -1020 2933 -994
rect 2997 -998 3059 -986
rect 3071 -998 3146 -986
rect 3204 -998 3279 -986
rect 3291 -998 3322 -986
rect 3328 -998 3363 -986
rect 2997 -1000 3159 -998
rect 2892 -1028 2933 -1020
rect 3015 -1024 3028 -1000
rect 3043 -1002 3058 -1000
rect 2855 -1038 2856 -1028
rect 2871 -1038 2884 -1028
rect 2898 -1038 2899 -1028
rect 2914 -1038 2927 -1028
rect 2942 -1038 2972 -1024
rect 3015 -1038 3058 -1024
rect 3082 -1027 3089 -1020
rect 3092 -1024 3159 -1000
rect 3191 -1000 3363 -998
rect 3161 -1022 3189 -1018
rect 3191 -1022 3271 -1000
rect 3292 -1002 3307 -1000
rect 3161 -1024 3271 -1022
rect 3092 -1028 3271 -1024
rect 3065 -1038 3095 -1028
rect 3097 -1038 3250 -1028
rect 3258 -1038 3288 -1028
rect 3292 -1038 3322 -1024
rect 3350 -1038 3363 -1000
rect 3435 -994 3470 -986
rect 3435 -1020 3436 -994
rect 3443 -1020 3470 -994
rect 3378 -1038 3408 -1024
rect 3435 -1028 3470 -1020
rect 3472 -994 3513 -986
rect 3472 -1020 3487 -994
rect 3494 -1020 3513 -994
rect 3577 -998 3639 -986
rect 3651 -998 3726 -986
rect 3784 -998 3859 -986
rect 3871 -998 3902 -986
rect 3908 -998 3943 -986
rect 3577 -1000 3739 -998
rect 3472 -1028 3513 -1020
rect 3595 -1024 3608 -1000
rect 3623 -1002 3638 -1000
rect 3435 -1038 3436 -1028
rect 3451 -1038 3464 -1028
rect 3478 -1038 3479 -1028
rect 3494 -1038 3507 -1028
rect 3522 -1038 3552 -1024
rect 3595 -1038 3638 -1024
rect 3662 -1027 3669 -1020
rect 3672 -1024 3739 -1000
rect 3771 -1000 3943 -998
rect 3741 -1022 3769 -1018
rect 3771 -1022 3851 -1000
rect 3872 -1002 3887 -1000
rect 3741 -1024 3851 -1022
rect 3672 -1028 3851 -1024
rect 3645 -1038 3675 -1028
rect 3677 -1038 3830 -1028
rect 3838 -1038 3868 -1028
rect 3872 -1038 3902 -1024
rect 3930 -1038 3943 -1000
rect 4015 -994 4050 -986
rect 4015 -1020 4016 -994
rect 4023 -1020 4050 -994
rect 3958 -1038 3988 -1024
rect 4015 -1028 4050 -1020
rect 4052 -994 4093 -986
rect 4052 -1020 4067 -994
rect 4074 -1020 4093 -994
rect 4157 -998 4219 -986
rect 4231 -998 4306 -986
rect 4364 -998 4439 -986
rect 4451 -998 4482 -986
rect 4488 -998 4523 -986
rect 4157 -1000 4319 -998
rect 4052 -1028 4093 -1020
rect 4175 -1024 4188 -1000
rect 4203 -1002 4218 -1000
rect 4015 -1038 4016 -1028
rect 4031 -1038 4044 -1028
rect 4058 -1038 4059 -1028
rect 4074 -1038 4087 -1028
rect 4102 -1038 4132 -1024
rect 4175 -1038 4218 -1024
rect 4242 -1027 4249 -1020
rect 4252 -1024 4319 -1000
rect 4351 -1000 4523 -998
rect 4321 -1022 4349 -1018
rect 4351 -1022 4431 -1000
rect 4452 -1002 4467 -1000
rect 4321 -1024 4431 -1022
rect 4252 -1028 4431 -1024
rect 4225 -1038 4255 -1028
rect 4257 -1038 4410 -1028
rect 4418 -1038 4448 -1028
rect 4452 -1038 4482 -1024
rect 4510 -1038 4523 -1000
rect 4595 -994 4630 -986
rect 4638 -987 4639 -971
rect 4654 -987 4667 -965
rect 4682 -987 4712 -965
rect 4755 -969 4817 -953
rect 4845 -960 4856 -944
rect 4861 -949 4871 -929
rect 4881 -949 4895 -929
rect 4898 -942 4907 -929
rect 4923 -942 4932 -929
rect 4861 -960 4895 -949
rect 4898 -960 4907 -944
rect 4923 -960 4932 -944
rect 4939 -949 4949 -929
rect 4959 -949 4973 -929
rect 4974 -942 4985 -929
rect 4939 -960 4973 -949
rect 4974 -960 4985 -944
rect 5031 -953 5047 -937
rect 5054 -939 5084 -887
rect 5118 -891 5119 -884
rect 5103 -899 5119 -891
rect 5090 -931 5103 -912
rect 5118 -931 5148 -915
rect 5090 -947 5164 -931
rect 5090 -949 5103 -947
rect 5118 -949 5152 -947
rect 4755 -971 4768 -969
rect 4783 -971 4817 -969
rect 4755 -987 4817 -971
rect 4861 -976 4877 -973
rect 4939 -976 4969 -965
rect 5017 -969 5063 -953
rect 5090 -965 5164 -949
rect 5017 -971 5051 -969
rect 5016 -987 5063 -971
rect 5090 -987 5103 -965
rect 5118 -987 5148 -965
rect 5175 -987 5176 -971
rect 5191 -987 5204 -827
rect 5234 -931 5247 -827
rect 5292 -849 5293 -839
rect 5313 -841 5321 -839
rect 5311 -843 5321 -841
rect 5308 -849 5321 -843
rect 5292 -853 5321 -849
rect 5326 -853 5356 -827
rect 5374 -841 5390 -839
rect 5462 -841 5513 -827
rect 5463 -843 5527 -841
rect 5570 -843 5585 -827
rect 5634 -830 5664 -827
rect 5634 -833 5670 -830
rect 5600 -841 5616 -839
rect 5374 -853 5389 -849
rect 5292 -855 5389 -853
rect 5417 -855 5585 -843
rect 5601 -853 5616 -849
rect 5634 -852 5673 -833
rect 5692 -839 5699 -838
rect 5698 -846 5699 -839
rect 5682 -849 5683 -846
rect 5698 -849 5711 -846
rect 5634 -853 5664 -852
rect 5673 -853 5679 -852
rect 5682 -853 5711 -849
rect 5601 -854 5711 -853
rect 5601 -855 5717 -854
rect 5276 -863 5327 -855
rect 5276 -875 5301 -863
rect 5308 -875 5327 -863
rect 5358 -863 5408 -855
rect 5358 -871 5374 -863
rect 5381 -865 5408 -863
rect 5417 -865 5638 -855
rect 5381 -875 5638 -865
rect 5667 -863 5717 -855
rect 5667 -872 5683 -863
rect 5276 -883 5327 -875
rect 5374 -883 5638 -875
rect 5664 -875 5683 -872
rect 5690 -875 5717 -863
rect 5664 -883 5717 -875
rect 5292 -891 5293 -883
rect 5308 -891 5321 -883
rect 5292 -899 5308 -891
rect 5289 -906 5308 -903
rect 5289 -915 5311 -906
rect 5262 -925 5311 -915
rect 5262 -931 5292 -925
rect 5311 -930 5316 -925
rect 5234 -947 5308 -931
rect 5326 -939 5356 -883
rect 5391 -893 5599 -883
rect 5634 -887 5679 -883
rect 5682 -884 5683 -883
rect 5698 -884 5711 -883
rect 5417 -923 5606 -893
rect 5432 -926 5606 -923
rect 5425 -929 5606 -926
rect 5234 -949 5247 -947
rect 5262 -949 5296 -947
rect 5234 -965 5308 -949
rect 5335 -953 5348 -939
rect 5363 -953 5379 -937
rect 5425 -942 5436 -929
rect 5218 -987 5219 -971
rect 5234 -987 5247 -965
rect 5262 -987 5292 -965
rect 5335 -969 5397 -953
rect 5425 -960 5436 -944
rect 5441 -949 5451 -929
rect 5461 -949 5475 -929
rect 5478 -942 5487 -929
rect 5503 -942 5512 -929
rect 5441 -960 5475 -949
rect 5478 -960 5487 -944
rect 5503 -960 5512 -944
rect 5519 -949 5529 -929
rect 5539 -949 5553 -929
rect 5554 -942 5565 -929
rect 5519 -960 5553 -949
rect 5554 -960 5565 -944
rect 5611 -953 5627 -937
rect 5634 -939 5664 -887
rect 5698 -891 5699 -884
rect 5683 -899 5699 -891
rect 5670 -931 5683 -912
rect 5698 -931 5728 -915
rect 5670 -947 5744 -931
rect 5670 -949 5683 -947
rect 5698 -949 5732 -947
rect 5335 -971 5348 -969
rect 5363 -971 5397 -969
rect 5335 -987 5397 -971
rect 5441 -976 5457 -973
rect 5519 -976 5549 -965
rect 5597 -969 5643 -953
rect 5670 -965 5744 -949
rect 5597 -971 5631 -969
rect 5596 -987 5643 -971
rect 5670 -987 5683 -965
rect 5698 -987 5728 -965
rect 5755 -987 5756 -971
rect 5771 -987 5784 -827
rect 5814 -931 5827 -827
rect 5872 -849 5873 -839
rect 5893 -841 5901 -839
rect 5891 -843 5901 -841
rect 5888 -849 5901 -843
rect 5872 -853 5901 -849
rect 5906 -853 5936 -827
rect 5954 -841 5970 -839
rect 6042 -841 6093 -827
rect 6043 -843 6107 -841
rect 6150 -843 6165 -827
rect 6214 -830 6244 -827
rect 6214 -833 6250 -830
rect 6180 -841 6196 -839
rect 5954 -853 5969 -849
rect 5872 -855 5969 -853
rect 5997 -855 6165 -843
rect 6181 -853 6196 -849
rect 6214 -852 6253 -833
rect 6272 -839 6279 -838
rect 6278 -846 6279 -839
rect 6262 -849 6263 -846
rect 6278 -849 6291 -846
rect 6214 -853 6244 -852
rect 6253 -853 6259 -852
rect 6262 -853 6291 -849
rect 6181 -854 6291 -853
rect 6181 -855 6297 -854
rect 5856 -863 5907 -855
rect 5856 -875 5881 -863
rect 5888 -875 5907 -863
rect 5938 -863 5988 -855
rect 5938 -871 5954 -863
rect 5961 -865 5988 -863
rect 5997 -865 6218 -855
rect 5961 -875 6218 -865
rect 6247 -863 6297 -855
rect 6247 -872 6263 -863
rect 5856 -883 5907 -875
rect 5954 -883 6218 -875
rect 6244 -875 6263 -872
rect 6270 -875 6297 -863
rect 6244 -883 6297 -875
rect 5872 -891 5873 -883
rect 5888 -891 5901 -883
rect 5872 -899 5888 -891
rect 5869 -906 5888 -903
rect 5869 -915 5891 -906
rect 5842 -925 5891 -915
rect 5842 -931 5872 -925
rect 5891 -930 5896 -925
rect 5814 -947 5888 -931
rect 5906 -939 5936 -883
rect 5971 -893 6179 -883
rect 6214 -887 6259 -883
rect 6262 -884 6263 -883
rect 6278 -884 6291 -883
rect 5997 -923 6186 -893
rect 6012 -926 6186 -923
rect 6005 -929 6186 -926
rect 5814 -949 5827 -947
rect 5842 -949 5876 -947
rect 5814 -965 5888 -949
rect 5915 -953 5928 -939
rect 5943 -953 5959 -937
rect 6005 -942 6016 -929
rect 5798 -987 5799 -971
rect 5814 -987 5827 -965
rect 5842 -987 5872 -965
rect 5915 -969 5977 -953
rect 6005 -960 6016 -944
rect 6021 -949 6031 -929
rect 6041 -949 6055 -929
rect 6058 -942 6067 -929
rect 6083 -942 6092 -929
rect 6021 -960 6055 -949
rect 6058 -960 6067 -944
rect 6083 -960 6092 -944
rect 6099 -949 6109 -929
rect 6119 -949 6133 -929
rect 6134 -942 6145 -929
rect 6099 -960 6133 -949
rect 6134 -960 6145 -944
rect 6191 -953 6207 -937
rect 6214 -939 6244 -887
rect 6278 -891 6279 -884
rect 6263 -899 6279 -891
rect 6250 -931 6263 -912
rect 6278 -931 6308 -915
rect 6250 -947 6324 -931
rect 6250 -949 6263 -947
rect 6278 -949 6312 -947
rect 5915 -971 5928 -969
rect 5943 -971 5977 -969
rect 5915 -987 5977 -971
rect 6021 -976 6037 -973
rect 6099 -976 6129 -965
rect 6177 -969 6223 -953
rect 6250 -965 6324 -949
rect 6177 -971 6211 -969
rect 6176 -987 6223 -971
rect 6250 -987 6263 -965
rect 6278 -987 6308 -965
rect 6335 -987 6336 -971
rect 6351 -987 6364 -827
rect 6394 -931 6407 -827
rect 6452 -849 6453 -839
rect 6473 -841 6481 -839
rect 6471 -843 6481 -841
rect 6468 -849 6481 -843
rect 6452 -853 6481 -849
rect 6486 -853 6516 -827
rect 6534 -841 6550 -839
rect 6622 -841 6673 -827
rect 6623 -843 6687 -841
rect 6730 -843 6745 -827
rect 6794 -830 6824 -827
rect 6794 -833 6830 -830
rect 6760 -841 6776 -839
rect 6534 -853 6549 -849
rect 6452 -855 6549 -853
rect 6577 -855 6745 -843
rect 6761 -853 6776 -849
rect 6794 -852 6833 -833
rect 6852 -839 6859 -838
rect 6858 -846 6859 -839
rect 6842 -849 6843 -846
rect 6858 -849 6871 -846
rect 6794 -853 6824 -852
rect 6833 -853 6839 -852
rect 6842 -853 6871 -849
rect 6761 -854 6871 -853
rect 6761 -855 6877 -854
rect 6436 -863 6487 -855
rect 6436 -875 6461 -863
rect 6468 -875 6487 -863
rect 6518 -863 6568 -855
rect 6518 -871 6534 -863
rect 6541 -865 6568 -863
rect 6577 -865 6798 -855
rect 6541 -875 6798 -865
rect 6827 -863 6877 -855
rect 6827 -872 6843 -863
rect 6436 -883 6487 -875
rect 6534 -883 6798 -875
rect 6824 -875 6843 -872
rect 6850 -875 6877 -863
rect 6824 -883 6877 -875
rect 6452 -891 6453 -883
rect 6468 -891 6481 -883
rect 6452 -899 6468 -891
rect 6449 -906 6468 -903
rect 6449 -915 6471 -906
rect 6422 -925 6471 -915
rect 6422 -931 6452 -925
rect 6471 -930 6476 -925
rect 6394 -947 6468 -931
rect 6486 -939 6516 -883
rect 6551 -893 6759 -883
rect 6794 -887 6839 -883
rect 6842 -884 6843 -883
rect 6858 -884 6871 -883
rect 6577 -923 6766 -893
rect 6592 -926 6766 -923
rect 6585 -929 6766 -926
rect 6394 -949 6407 -947
rect 6422 -949 6456 -947
rect 6394 -965 6468 -949
rect 6495 -953 6508 -939
rect 6523 -953 6539 -937
rect 6585 -942 6596 -929
rect 6378 -987 6379 -971
rect 6394 -987 6407 -965
rect 6422 -987 6452 -965
rect 6495 -969 6557 -953
rect 6585 -960 6596 -944
rect 6601 -949 6611 -929
rect 6621 -949 6635 -929
rect 6638 -942 6647 -929
rect 6663 -942 6672 -929
rect 6601 -960 6635 -949
rect 6638 -960 6647 -944
rect 6663 -960 6672 -944
rect 6679 -949 6689 -929
rect 6699 -949 6713 -929
rect 6714 -942 6725 -929
rect 6679 -960 6713 -949
rect 6714 -960 6725 -944
rect 6771 -953 6787 -937
rect 6794 -939 6824 -887
rect 6858 -891 6859 -884
rect 6843 -899 6859 -891
rect 6830 -931 6843 -912
rect 6858 -931 6888 -915
rect 6830 -947 6904 -931
rect 6830 -949 6843 -947
rect 6858 -949 6892 -947
rect 6495 -971 6508 -969
rect 6523 -971 6557 -969
rect 6495 -987 6557 -971
rect 6601 -976 6617 -973
rect 6679 -976 6709 -965
rect 6757 -969 6803 -953
rect 6830 -965 6904 -949
rect 6757 -971 6791 -969
rect 6756 -987 6803 -971
rect 6830 -987 6843 -965
rect 6858 -987 6888 -965
rect 6915 -987 6916 -971
rect 6931 -987 6944 -827
rect 4595 -1020 4596 -994
rect 4603 -1020 4630 -994
rect 4538 -1038 4568 -1024
rect 4595 -1028 4630 -1020
rect 4632 -995 4673 -987
rect 4632 -1021 4647 -995
rect 4654 -1021 4673 -995
rect 4737 -999 4799 -987
rect 4811 -999 4886 -987
rect 4944 -999 5019 -987
rect 5031 -999 5062 -987
rect 5068 -999 5103 -987
rect 4737 -1001 4899 -999
rect 4755 -1019 4768 -1001
rect 4783 -1003 4798 -1001
rect 4595 -1038 4596 -1028
rect 4611 -1038 4624 -1028
rect 4632 -1029 4673 -1021
rect 4756 -1025 4768 -1019
rect 4832 -1019 4899 -1001
rect 4931 -1001 5103 -999
rect 4931 -1019 5011 -1001
rect 5032 -1003 5047 -1001
rect -2 -1039 4624 -1038
rect 4638 -1039 4639 -1029
rect 4654 -1039 4667 -1029
rect 4682 -1039 4712 -1025
rect 4756 -1039 4798 -1025
rect 4822 -1028 4829 -1021
rect 4832 -1029 5011 -1019
rect 4805 -1039 4835 -1029
rect 4837 -1039 4990 -1029
rect 4998 -1039 5028 -1029
rect 5032 -1039 5062 -1025
rect 5090 -1039 5103 -1001
rect 5175 -995 5210 -987
rect 5175 -1021 5176 -995
rect 5183 -1021 5210 -995
rect 5118 -1039 5148 -1025
rect 5175 -1029 5210 -1021
rect 5212 -995 5253 -987
rect 5212 -1021 5227 -995
rect 5234 -1021 5253 -995
rect 5317 -999 5379 -987
rect 5391 -999 5466 -987
rect 5524 -999 5599 -987
rect 5611 -999 5642 -987
rect 5648 -999 5683 -987
rect 5317 -1001 5479 -999
rect 5335 -1019 5348 -1001
rect 5363 -1003 5378 -1001
rect 5212 -1029 5253 -1021
rect 5336 -1025 5348 -1019
rect 5412 -1019 5479 -1001
rect 5511 -1001 5683 -999
rect 5511 -1019 5591 -1001
rect 5612 -1003 5627 -1001
rect 5175 -1039 5176 -1029
rect 5191 -1039 5204 -1029
rect 5218 -1039 5219 -1029
rect 5234 -1039 5247 -1029
rect 5262 -1039 5292 -1025
rect 5336 -1039 5378 -1025
rect 5402 -1028 5409 -1021
rect 5412 -1029 5591 -1019
rect 5385 -1039 5415 -1029
rect 5417 -1039 5570 -1029
rect 5578 -1039 5608 -1029
rect 5612 -1039 5642 -1025
rect 5670 -1039 5683 -1001
rect 5755 -995 5790 -987
rect 5755 -1021 5756 -995
rect 5763 -1021 5790 -995
rect 5698 -1039 5728 -1025
rect 5755 -1029 5790 -1021
rect 5792 -995 5833 -987
rect 5792 -1021 5807 -995
rect 5814 -1021 5833 -995
rect 5897 -999 5959 -987
rect 5971 -999 6046 -987
rect 6104 -999 6179 -987
rect 6191 -999 6222 -987
rect 6228 -999 6263 -987
rect 5897 -1001 6059 -999
rect 5915 -1019 5928 -1001
rect 5943 -1003 5958 -1001
rect 5792 -1029 5833 -1021
rect 5916 -1025 5928 -1019
rect 5992 -1019 6059 -1001
rect 6091 -1001 6263 -999
rect 6091 -1019 6171 -1001
rect 6192 -1003 6207 -1001
rect 5755 -1039 5756 -1029
rect 5771 -1039 5784 -1029
rect 5798 -1039 5799 -1029
rect 5814 -1039 5827 -1029
rect 5842 -1039 5872 -1025
rect 5916 -1039 5958 -1025
rect 5982 -1028 5989 -1021
rect 5992 -1029 6171 -1019
rect 5965 -1039 5995 -1029
rect 5997 -1039 6150 -1029
rect 6158 -1039 6188 -1029
rect 6192 -1039 6222 -1025
rect 6250 -1039 6263 -1001
rect 6335 -995 6370 -987
rect 6335 -1021 6336 -995
rect 6343 -1021 6370 -995
rect 6278 -1039 6308 -1025
rect 6335 -1029 6370 -1021
rect 6372 -995 6413 -987
rect 6372 -1021 6387 -995
rect 6394 -1021 6413 -995
rect 6477 -999 6539 -987
rect 6551 -999 6626 -987
rect 6684 -999 6759 -987
rect 6771 -999 6802 -987
rect 6808 -999 6843 -987
rect 6477 -1001 6639 -999
rect 6495 -1019 6508 -1001
rect 6523 -1003 6538 -1001
rect 6372 -1029 6413 -1021
rect 6496 -1025 6508 -1019
rect 6572 -1019 6639 -1001
rect 6671 -1001 6843 -999
rect 6671 -1019 6751 -1001
rect 6772 -1003 6787 -1001
rect 6335 -1039 6336 -1029
rect 6351 -1039 6364 -1029
rect 6378 -1039 6379 -1029
rect 6394 -1039 6407 -1029
rect 6422 -1039 6452 -1025
rect 6496 -1039 6538 -1025
rect 6562 -1028 6569 -1021
rect 6572 -1029 6751 -1019
rect 6545 -1039 6575 -1029
rect 6577 -1039 6730 -1029
rect 6738 -1039 6768 -1029
rect 6772 -1039 6802 -1025
rect 6830 -1039 6843 -1001
rect 6915 -995 6950 -987
rect 6915 -1021 6916 -995
rect 6923 -1021 6950 -995
rect 6858 -1039 6888 -1025
rect 6915 -1029 6950 -1021
rect 6915 -1039 6916 -1029
rect 6931 -1039 6944 -1029
rect -2 -1044 6944 -1039
rect -1 -1052 6944 -1044
rect 14 -1082 27 -1052
rect 42 -1070 72 -1052
rect 115 -1066 129 -1052
rect 165 -1066 385 -1052
rect 116 -1068 129 -1066
rect 82 -1080 97 -1068
rect 79 -1082 101 -1080
rect 106 -1082 136 -1068
rect 197 -1070 350 -1066
rect 179 -1082 371 -1070
rect 414 -1082 444 -1068
rect 450 -1082 463 -1052
rect 478 -1070 508 -1052
rect 551 -1082 564 -1052
rect 594 -1082 607 -1052
rect 622 -1070 652 -1052
rect 695 -1066 709 -1052
rect 745 -1066 965 -1052
rect 696 -1068 709 -1066
rect 662 -1080 677 -1068
rect 659 -1082 681 -1080
rect 686 -1082 716 -1068
rect 777 -1070 930 -1066
rect 759 -1082 951 -1070
rect 994 -1082 1024 -1068
rect 1030 -1082 1043 -1052
rect 1058 -1070 1088 -1052
rect 1131 -1082 1144 -1052
rect 1174 -1082 1187 -1052
rect 1202 -1070 1232 -1052
rect 1275 -1066 1289 -1052
rect 1325 -1066 1545 -1052
rect 1276 -1068 1289 -1066
rect 1242 -1080 1257 -1068
rect 1239 -1082 1261 -1080
rect 1266 -1082 1296 -1068
rect 1357 -1070 1510 -1066
rect 1339 -1082 1531 -1070
rect 1574 -1082 1604 -1068
rect 1610 -1082 1623 -1052
rect 1638 -1070 1668 -1052
rect 1711 -1082 1724 -1052
rect 1754 -1082 1767 -1052
rect 1782 -1070 1812 -1052
rect 1855 -1066 1869 -1052
rect 1905 -1066 2125 -1052
rect 1856 -1068 1869 -1066
rect 1822 -1080 1837 -1068
rect 1819 -1082 1841 -1080
rect 1846 -1082 1876 -1068
rect 1937 -1070 2090 -1066
rect 1919 -1082 2111 -1070
rect 2154 -1082 2184 -1068
rect 2190 -1082 2203 -1052
rect 2218 -1070 2248 -1052
rect 2291 -1082 2304 -1052
rect 2334 -1082 2347 -1052
rect 2362 -1070 2392 -1052
rect 2435 -1066 2449 -1052
rect 2485 -1066 2705 -1052
rect 2436 -1068 2449 -1066
rect 2402 -1080 2417 -1068
rect 2399 -1082 2421 -1080
rect 2426 -1082 2456 -1068
rect 2517 -1070 2670 -1066
rect 2499 -1082 2691 -1070
rect 2734 -1082 2764 -1068
rect 2770 -1082 2783 -1052
rect 2798 -1070 2828 -1052
rect 2871 -1082 2884 -1052
rect 2914 -1082 2927 -1052
rect 2942 -1070 2972 -1052
rect 3015 -1066 3029 -1052
rect 3065 -1066 3285 -1052
rect 3016 -1068 3029 -1066
rect 2982 -1080 2997 -1068
rect 2979 -1082 3001 -1080
rect 3006 -1082 3036 -1068
rect 3097 -1070 3250 -1066
rect 3079 -1082 3271 -1070
rect 3314 -1082 3344 -1068
rect 3350 -1082 3363 -1052
rect 3378 -1070 3408 -1052
rect 3451 -1082 3464 -1052
rect 3494 -1082 3507 -1052
rect 3522 -1070 3552 -1052
rect 3595 -1066 3609 -1052
rect 3645 -1066 3865 -1052
rect 3596 -1068 3609 -1066
rect 3562 -1080 3577 -1068
rect 3559 -1082 3581 -1080
rect 3586 -1082 3616 -1068
rect 3677 -1070 3830 -1066
rect 3659 -1082 3851 -1070
rect 3894 -1082 3924 -1068
rect 3930 -1082 3943 -1052
rect 3958 -1070 3988 -1052
rect 4031 -1082 4044 -1052
rect 4074 -1082 4087 -1052
rect 4102 -1070 4132 -1052
rect 4175 -1066 4189 -1052
rect 4225 -1066 4445 -1052
rect 4176 -1068 4189 -1066
rect 4142 -1080 4157 -1068
rect 4139 -1082 4161 -1080
rect 4166 -1082 4196 -1068
rect 4257 -1070 4410 -1066
rect 4239 -1082 4431 -1070
rect 4474 -1082 4504 -1068
rect 4510 -1082 4523 -1052
rect 4538 -1070 4568 -1052
rect 4611 -1053 6944 -1052
rect 4611 -1082 4624 -1053
rect -1 -1083 4624 -1082
rect 4654 -1083 4667 -1053
rect 4682 -1071 4712 -1053
rect 4756 -1069 4769 -1053
rect 4805 -1067 5025 -1053
rect 4722 -1081 4737 -1069
rect 4719 -1083 4741 -1081
rect 4746 -1083 4776 -1069
rect 4837 -1071 4990 -1067
rect 4819 -1083 5011 -1071
rect 5054 -1083 5084 -1069
rect 5090 -1083 5103 -1053
rect 5118 -1071 5148 -1053
rect 5191 -1083 5204 -1053
rect 5234 -1083 5247 -1053
rect 5262 -1071 5292 -1053
rect 5336 -1069 5349 -1053
rect 5385 -1067 5605 -1053
rect 5302 -1081 5317 -1069
rect 5299 -1083 5321 -1081
rect 5326 -1083 5356 -1069
rect 5417 -1071 5570 -1067
rect 5399 -1083 5591 -1071
rect 5634 -1083 5664 -1069
rect 5670 -1083 5683 -1053
rect 5698 -1071 5728 -1053
rect 5771 -1083 5784 -1053
rect 5814 -1083 5827 -1053
rect 5842 -1071 5872 -1053
rect 5916 -1069 5929 -1053
rect 5965 -1067 6185 -1053
rect 5882 -1081 5897 -1069
rect 5879 -1083 5901 -1081
rect 5906 -1083 5936 -1069
rect 5997 -1071 6150 -1067
rect 5979 -1083 6171 -1071
rect 6214 -1083 6244 -1069
rect 6250 -1083 6263 -1053
rect 6278 -1071 6308 -1053
rect 6351 -1083 6364 -1053
rect 6394 -1083 6407 -1053
rect 6422 -1071 6452 -1053
rect 6496 -1069 6509 -1053
rect 6545 -1067 6765 -1053
rect 6462 -1081 6477 -1069
rect 6459 -1083 6481 -1081
rect 6486 -1083 6516 -1069
rect 6577 -1071 6730 -1067
rect 6559 -1083 6751 -1071
rect 6794 -1083 6824 -1069
rect 6830 -1083 6843 -1053
rect 6858 -1071 6888 -1053
rect 6931 -1083 6944 -1053
rect -1 -1096 6944 -1083
rect 14 -1200 27 -1096
rect 72 -1118 73 -1108
rect 88 -1118 101 -1108
rect 72 -1122 101 -1118
rect 106 -1122 136 -1096
rect 154 -1110 170 -1108
rect 242 -1110 295 -1096
rect 243 -1112 307 -1110
rect 350 -1112 365 -1096
rect 414 -1099 444 -1096
rect 414 -1102 450 -1099
rect 380 -1110 396 -1108
rect 154 -1122 169 -1118
rect 72 -1124 169 -1122
rect 197 -1124 365 -1112
rect 381 -1122 396 -1118
rect 414 -1121 453 -1102
rect 472 -1108 479 -1107
rect 478 -1115 479 -1108
rect 462 -1118 463 -1115
rect 478 -1118 491 -1115
rect 414 -1122 444 -1121
rect 453 -1122 459 -1121
rect 462 -1122 491 -1118
rect 381 -1123 491 -1122
rect 381 -1124 497 -1123
rect 56 -1132 107 -1124
rect 56 -1144 81 -1132
rect 88 -1144 107 -1132
rect 138 -1132 188 -1124
rect 138 -1140 154 -1132
rect 161 -1134 188 -1132
rect 197 -1134 418 -1124
rect 161 -1144 418 -1134
rect 447 -1132 497 -1124
rect 447 -1141 463 -1132
rect 56 -1152 107 -1144
rect 154 -1152 418 -1144
rect 444 -1144 463 -1141
rect 470 -1144 497 -1132
rect 444 -1152 497 -1144
rect 72 -1160 73 -1152
rect 88 -1160 101 -1152
rect 72 -1168 88 -1160
rect 69 -1175 88 -1172
rect 69 -1184 91 -1175
rect 42 -1194 91 -1184
rect 42 -1200 72 -1194
rect 91 -1199 96 -1194
rect 14 -1216 88 -1200
rect 106 -1208 136 -1152
rect 171 -1162 379 -1152
rect 414 -1156 459 -1152
rect 462 -1153 463 -1152
rect 478 -1153 491 -1152
rect 197 -1192 386 -1162
rect 212 -1195 386 -1192
rect 205 -1198 386 -1195
rect 14 -1218 27 -1216
rect 42 -1218 76 -1216
rect 14 -1234 88 -1218
rect 115 -1222 128 -1208
rect 143 -1222 159 -1206
rect 205 -1211 216 -1198
rect 14 -1256 27 -1234
rect 42 -1256 72 -1234
rect 115 -1238 177 -1222
rect 205 -1229 216 -1213
rect 221 -1218 231 -1198
rect 241 -1218 255 -1198
rect 258 -1211 267 -1198
rect 283 -1211 292 -1198
rect 221 -1229 255 -1218
rect 258 -1229 267 -1213
rect 283 -1229 292 -1213
rect 299 -1218 309 -1198
rect 319 -1218 333 -1198
rect 334 -1211 345 -1198
rect 299 -1229 333 -1218
rect 334 -1229 345 -1213
rect 391 -1222 407 -1206
rect 414 -1208 444 -1156
rect 478 -1160 479 -1153
rect 463 -1168 479 -1160
rect 450 -1200 463 -1181
rect 478 -1200 508 -1184
rect 450 -1216 524 -1200
rect 450 -1218 463 -1216
rect 478 -1218 512 -1216
rect 115 -1240 128 -1238
rect 143 -1240 177 -1238
rect 115 -1256 177 -1240
rect 221 -1245 237 -1242
rect 299 -1245 329 -1234
rect 377 -1238 423 -1222
rect 450 -1234 524 -1218
rect 377 -1240 411 -1238
rect 376 -1256 423 -1240
rect 450 -1256 463 -1234
rect 478 -1256 508 -1234
rect 535 -1256 536 -1240
rect 551 -1256 564 -1096
rect 594 -1200 607 -1096
rect 652 -1118 653 -1108
rect 668 -1118 681 -1108
rect 652 -1122 681 -1118
rect 686 -1122 716 -1096
rect 734 -1110 750 -1108
rect 822 -1110 875 -1096
rect 823 -1112 887 -1110
rect 930 -1112 945 -1096
rect 994 -1099 1024 -1096
rect 994 -1102 1030 -1099
rect 960 -1110 976 -1108
rect 734 -1122 749 -1118
rect 652 -1124 749 -1122
rect 777 -1124 945 -1112
rect 961 -1122 976 -1118
rect 994 -1121 1033 -1102
rect 1052 -1108 1059 -1107
rect 1058 -1115 1059 -1108
rect 1042 -1118 1043 -1115
rect 1058 -1118 1071 -1115
rect 994 -1122 1024 -1121
rect 1033 -1122 1039 -1121
rect 1042 -1122 1071 -1118
rect 961 -1123 1071 -1122
rect 961 -1124 1077 -1123
rect 636 -1132 687 -1124
rect 636 -1144 661 -1132
rect 668 -1144 687 -1132
rect 718 -1132 768 -1124
rect 718 -1140 734 -1132
rect 741 -1134 768 -1132
rect 777 -1134 998 -1124
rect 741 -1144 998 -1134
rect 1027 -1132 1077 -1124
rect 1027 -1141 1043 -1132
rect 636 -1152 687 -1144
rect 734 -1152 998 -1144
rect 1024 -1144 1043 -1141
rect 1050 -1144 1077 -1132
rect 1024 -1152 1077 -1144
rect 652 -1160 653 -1152
rect 668 -1160 681 -1152
rect 652 -1168 668 -1160
rect 649 -1175 668 -1172
rect 649 -1184 671 -1175
rect 622 -1194 671 -1184
rect 622 -1200 652 -1194
rect 671 -1199 676 -1194
rect 594 -1216 668 -1200
rect 686 -1208 716 -1152
rect 751 -1162 959 -1152
rect 994 -1156 1039 -1152
rect 1042 -1153 1043 -1152
rect 1058 -1153 1071 -1152
rect 777 -1192 966 -1162
rect 792 -1195 966 -1192
rect 785 -1198 966 -1195
rect 594 -1218 607 -1216
rect 622 -1218 656 -1216
rect 594 -1234 668 -1218
rect 695 -1222 708 -1208
rect 723 -1222 739 -1206
rect 785 -1211 796 -1198
rect 578 -1256 579 -1240
rect 594 -1256 607 -1234
rect 622 -1256 652 -1234
rect 695 -1238 757 -1222
rect 785 -1229 796 -1213
rect 801 -1218 811 -1198
rect 821 -1218 835 -1198
rect 838 -1211 847 -1198
rect 863 -1211 872 -1198
rect 801 -1229 835 -1218
rect 838 -1229 847 -1213
rect 863 -1229 872 -1213
rect 879 -1218 889 -1198
rect 899 -1218 913 -1198
rect 914 -1211 925 -1198
rect 879 -1229 913 -1218
rect 914 -1229 925 -1213
rect 971 -1222 987 -1206
rect 994 -1208 1024 -1156
rect 1058 -1160 1059 -1153
rect 1043 -1168 1059 -1160
rect 1030 -1200 1043 -1181
rect 1058 -1200 1088 -1184
rect 1030 -1216 1104 -1200
rect 1030 -1218 1043 -1216
rect 1058 -1218 1092 -1216
rect 695 -1240 708 -1238
rect 723 -1240 757 -1238
rect 695 -1256 757 -1240
rect 801 -1245 817 -1242
rect 879 -1245 909 -1234
rect 957 -1238 1003 -1222
rect 1030 -1234 1104 -1218
rect 957 -1240 991 -1238
rect 956 -1256 1003 -1240
rect 1030 -1256 1043 -1234
rect 1058 -1256 1088 -1234
rect 1115 -1256 1116 -1240
rect 1131 -1256 1144 -1096
rect 1174 -1200 1187 -1096
rect 1232 -1118 1233 -1108
rect 1248 -1118 1261 -1108
rect 1232 -1122 1261 -1118
rect 1266 -1122 1296 -1096
rect 1314 -1110 1330 -1108
rect 1402 -1110 1455 -1096
rect 1403 -1112 1467 -1110
rect 1510 -1112 1525 -1096
rect 1574 -1099 1604 -1096
rect 1574 -1102 1610 -1099
rect 1540 -1110 1556 -1108
rect 1314 -1122 1329 -1118
rect 1232 -1124 1329 -1122
rect 1357 -1124 1525 -1112
rect 1541 -1122 1556 -1118
rect 1574 -1121 1613 -1102
rect 1632 -1108 1639 -1107
rect 1638 -1115 1639 -1108
rect 1622 -1118 1623 -1115
rect 1638 -1118 1651 -1115
rect 1574 -1122 1604 -1121
rect 1613 -1122 1619 -1121
rect 1622 -1122 1651 -1118
rect 1541 -1123 1651 -1122
rect 1541 -1124 1657 -1123
rect 1216 -1132 1267 -1124
rect 1216 -1144 1241 -1132
rect 1248 -1144 1267 -1132
rect 1298 -1132 1348 -1124
rect 1298 -1140 1314 -1132
rect 1321 -1134 1348 -1132
rect 1357 -1134 1578 -1124
rect 1321 -1144 1578 -1134
rect 1607 -1132 1657 -1124
rect 1607 -1141 1623 -1132
rect 1216 -1152 1267 -1144
rect 1314 -1152 1578 -1144
rect 1604 -1144 1623 -1141
rect 1630 -1144 1657 -1132
rect 1604 -1152 1657 -1144
rect 1232 -1160 1233 -1152
rect 1248 -1160 1261 -1152
rect 1232 -1168 1248 -1160
rect 1229 -1175 1248 -1172
rect 1229 -1184 1251 -1175
rect 1202 -1194 1251 -1184
rect 1202 -1200 1232 -1194
rect 1251 -1199 1256 -1194
rect 1174 -1216 1248 -1200
rect 1266 -1208 1296 -1152
rect 1331 -1162 1539 -1152
rect 1574 -1156 1619 -1152
rect 1622 -1153 1623 -1152
rect 1638 -1153 1651 -1152
rect 1357 -1192 1546 -1162
rect 1372 -1195 1546 -1192
rect 1365 -1198 1546 -1195
rect 1174 -1218 1187 -1216
rect 1202 -1218 1236 -1216
rect 1174 -1234 1248 -1218
rect 1275 -1222 1288 -1208
rect 1303 -1222 1319 -1206
rect 1365 -1211 1376 -1198
rect 1158 -1256 1159 -1240
rect 1174 -1256 1187 -1234
rect 1202 -1256 1232 -1234
rect 1275 -1238 1337 -1222
rect 1365 -1229 1376 -1213
rect 1381 -1218 1391 -1198
rect 1401 -1218 1415 -1198
rect 1418 -1211 1427 -1198
rect 1443 -1211 1452 -1198
rect 1381 -1229 1415 -1218
rect 1418 -1229 1427 -1213
rect 1443 -1229 1452 -1213
rect 1459 -1218 1469 -1198
rect 1479 -1218 1493 -1198
rect 1494 -1211 1505 -1198
rect 1459 -1229 1493 -1218
rect 1494 -1229 1505 -1213
rect 1551 -1222 1567 -1206
rect 1574 -1208 1604 -1156
rect 1638 -1160 1639 -1153
rect 1623 -1168 1639 -1160
rect 1610 -1200 1623 -1181
rect 1638 -1200 1668 -1184
rect 1610 -1216 1684 -1200
rect 1610 -1218 1623 -1216
rect 1638 -1218 1672 -1216
rect 1275 -1240 1288 -1238
rect 1303 -1240 1337 -1238
rect 1275 -1256 1337 -1240
rect 1381 -1245 1397 -1242
rect 1459 -1245 1489 -1234
rect 1537 -1238 1583 -1222
rect 1610 -1234 1684 -1218
rect 1537 -1240 1571 -1238
rect 1536 -1256 1583 -1240
rect 1610 -1256 1623 -1234
rect 1638 -1256 1668 -1234
rect 1695 -1256 1696 -1240
rect 1711 -1256 1724 -1096
rect 1754 -1200 1767 -1096
rect 1812 -1118 1813 -1108
rect 1828 -1118 1841 -1108
rect 1812 -1122 1841 -1118
rect 1846 -1122 1876 -1096
rect 1894 -1110 1910 -1108
rect 1982 -1110 2035 -1096
rect 1983 -1112 2047 -1110
rect 2090 -1112 2105 -1096
rect 2154 -1099 2184 -1096
rect 2154 -1102 2190 -1099
rect 2120 -1110 2136 -1108
rect 1894 -1122 1909 -1118
rect 1812 -1124 1909 -1122
rect 1937 -1124 2105 -1112
rect 2121 -1122 2136 -1118
rect 2154 -1121 2193 -1102
rect 2212 -1108 2219 -1107
rect 2218 -1115 2219 -1108
rect 2202 -1118 2203 -1115
rect 2218 -1118 2231 -1115
rect 2154 -1122 2184 -1121
rect 2193 -1122 2199 -1121
rect 2202 -1122 2231 -1118
rect 2121 -1123 2231 -1122
rect 2121 -1124 2237 -1123
rect 1796 -1132 1847 -1124
rect 1796 -1144 1821 -1132
rect 1828 -1144 1847 -1132
rect 1878 -1132 1928 -1124
rect 1878 -1140 1894 -1132
rect 1901 -1134 1928 -1132
rect 1937 -1134 2158 -1124
rect 1901 -1144 2158 -1134
rect 2187 -1132 2237 -1124
rect 2187 -1141 2203 -1132
rect 1796 -1152 1847 -1144
rect 1894 -1152 2158 -1144
rect 2184 -1144 2203 -1141
rect 2210 -1144 2237 -1132
rect 2184 -1152 2237 -1144
rect 1812 -1160 1813 -1152
rect 1828 -1160 1841 -1152
rect 1812 -1168 1828 -1160
rect 1809 -1175 1828 -1172
rect 1809 -1184 1831 -1175
rect 1782 -1194 1831 -1184
rect 1782 -1200 1812 -1194
rect 1831 -1199 1836 -1194
rect 1754 -1216 1828 -1200
rect 1846 -1208 1876 -1152
rect 1911 -1162 2119 -1152
rect 2154 -1156 2199 -1152
rect 2202 -1153 2203 -1152
rect 2218 -1153 2231 -1152
rect 1937 -1192 2126 -1162
rect 1952 -1195 2126 -1192
rect 1945 -1198 2126 -1195
rect 1754 -1218 1767 -1216
rect 1782 -1218 1816 -1216
rect 1754 -1234 1828 -1218
rect 1855 -1222 1868 -1208
rect 1883 -1222 1899 -1206
rect 1945 -1211 1956 -1198
rect 1738 -1256 1739 -1240
rect 1754 -1256 1767 -1234
rect 1782 -1256 1812 -1234
rect 1855 -1238 1917 -1222
rect 1945 -1229 1956 -1213
rect 1961 -1218 1971 -1198
rect 1981 -1218 1995 -1198
rect 1998 -1211 2007 -1198
rect 2023 -1211 2032 -1198
rect 1961 -1229 1995 -1218
rect 1998 -1229 2007 -1213
rect 2023 -1229 2032 -1213
rect 2039 -1218 2049 -1198
rect 2059 -1218 2073 -1198
rect 2074 -1211 2085 -1198
rect 2039 -1229 2073 -1218
rect 2074 -1229 2085 -1213
rect 2131 -1222 2147 -1206
rect 2154 -1208 2184 -1156
rect 2218 -1160 2219 -1153
rect 2203 -1168 2219 -1160
rect 2190 -1200 2203 -1181
rect 2218 -1200 2248 -1184
rect 2190 -1216 2264 -1200
rect 2190 -1218 2203 -1216
rect 2218 -1218 2252 -1216
rect 1855 -1240 1868 -1238
rect 1883 -1240 1917 -1238
rect 1855 -1256 1917 -1240
rect 1961 -1245 1977 -1242
rect 2039 -1245 2069 -1234
rect 2117 -1238 2163 -1222
rect 2190 -1234 2264 -1218
rect 2117 -1240 2151 -1238
rect 2116 -1256 2163 -1240
rect 2190 -1256 2203 -1234
rect 2218 -1256 2248 -1234
rect 2275 -1256 2276 -1240
rect 2291 -1256 2304 -1096
rect 2334 -1200 2347 -1096
rect 2392 -1118 2393 -1108
rect 2408 -1118 2421 -1108
rect 2392 -1122 2421 -1118
rect 2426 -1122 2456 -1096
rect 2474 -1110 2490 -1108
rect 2562 -1110 2615 -1096
rect 2563 -1112 2627 -1110
rect 2670 -1112 2685 -1096
rect 2734 -1099 2764 -1096
rect 2734 -1102 2770 -1099
rect 2700 -1110 2716 -1108
rect 2474 -1122 2489 -1118
rect 2392 -1124 2489 -1122
rect 2517 -1124 2685 -1112
rect 2701 -1122 2716 -1118
rect 2734 -1121 2773 -1102
rect 2792 -1108 2799 -1107
rect 2798 -1115 2799 -1108
rect 2782 -1118 2783 -1115
rect 2798 -1118 2811 -1115
rect 2734 -1122 2764 -1121
rect 2773 -1122 2779 -1121
rect 2782 -1122 2811 -1118
rect 2701 -1123 2811 -1122
rect 2701 -1124 2817 -1123
rect 2376 -1132 2427 -1124
rect 2376 -1144 2401 -1132
rect 2408 -1144 2427 -1132
rect 2458 -1132 2508 -1124
rect 2458 -1140 2474 -1132
rect 2481 -1134 2508 -1132
rect 2517 -1134 2738 -1124
rect 2481 -1144 2738 -1134
rect 2767 -1132 2817 -1124
rect 2767 -1141 2783 -1132
rect 2376 -1152 2427 -1144
rect 2474 -1152 2738 -1144
rect 2764 -1144 2783 -1141
rect 2790 -1144 2817 -1132
rect 2764 -1152 2817 -1144
rect 2392 -1160 2393 -1152
rect 2408 -1160 2421 -1152
rect 2392 -1168 2408 -1160
rect 2389 -1175 2408 -1172
rect 2389 -1184 2411 -1175
rect 2362 -1194 2411 -1184
rect 2362 -1200 2392 -1194
rect 2411 -1199 2416 -1194
rect 2334 -1216 2408 -1200
rect 2426 -1208 2456 -1152
rect 2491 -1162 2699 -1152
rect 2734 -1156 2779 -1152
rect 2782 -1153 2783 -1152
rect 2798 -1153 2811 -1152
rect 2517 -1192 2706 -1162
rect 2532 -1195 2706 -1192
rect 2525 -1198 2706 -1195
rect 2334 -1218 2347 -1216
rect 2362 -1218 2396 -1216
rect 2334 -1234 2408 -1218
rect 2435 -1222 2448 -1208
rect 2463 -1222 2479 -1206
rect 2525 -1211 2536 -1198
rect 2318 -1256 2319 -1240
rect 2334 -1256 2347 -1234
rect 2362 -1256 2392 -1234
rect 2435 -1238 2497 -1222
rect 2525 -1229 2536 -1213
rect 2541 -1218 2551 -1198
rect 2561 -1218 2575 -1198
rect 2578 -1211 2587 -1198
rect 2603 -1211 2612 -1198
rect 2541 -1229 2575 -1218
rect 2578 -1229 2587 -1213
rect 2603 -1229 2612 -1213
rect 2619 -1218 2629 -1198
rect 2639 -1218 2653 -1198
rect 2654 -1211 2665 -1198
rect 2619 -1229 2653 -1218
rect 2654 -1229 2665 -1213
rect 2711 -1222 2727 -1206
rect 2734 -1208 2764 -1156
rect 2798 -1160 2799 -1153
rect 2783 -1168 2799 -1160
rect 2770 -1200 2783 -1181
rect 2798 -1200 2828 -1184
rect 2770 -1216 2844 -1200
rect 2770 -1218 2783 -1216
rect 2798 -1218 2832 -1216
rect 2435 -1240 2448 -1238
rect 2463 -1240 2497 -1238
rect 2435 -1256 2497 -1240
rect 2541 -1245 2557 -1242
rect 2619 -1245 2649 -1234
rect 2697 -1238 2743 -1222
rect 2770 -1234 2844 -1218
rect 2697 -1240 2731 -1238
rect 2696 -1256 2743 -1240
rect 2770 -1256 2783 -1234
rect 2798 -1256 2828 -1234
rect 2855 -1256 2856 -1240
rect 2871 -1256 2884 -1096
rect 2914 -1200 2927 -1096
rect 2972 -1118 2973 -1108
rect 2988 -1118 3001 -1108
rect 2972 -1122 3001 -1118
rect 3006 -1122 3036 -1096
rect 3054 -1110 3070 -1108
rect 3142 -1110 3195 -1096
rect 3143 -1112 3205 -1110
rect 3250 -1112 3265 -1096
rect 3314 -1099 3344 -1096
rect 3314 -1102 3350 -1099
rect 3280 -1110 3296 -1108
rect 3054 -1122 3069 -1118
rect 2972 -1124 3069 -1122
rect 3097 -1124 3265 -1112
rect 3281 -1122 3296 -1118
rect 3314 -1121 3353 -1102
rect 3372 -1108 3379 -1107
rect 3378 -1115 3379 -1108
rect 3362 -1118 3363 -1115
rect 3378 -1118 3391 -1115
rect 3314 -1122 3344 -1121
rect 3353 -1122 3359 -1121
rect 3362 -1122 3391 -1118
rect 3281 -1123 3391 -1122
rect 3281 -1124 3397 -1123
rect 2956 -1132 3007 -1124
rect 2956 -1144 2981 -1132
rect 2988 -1144 3007 -1132
rect 3038 -1132 3088 -1124
rect 3038 -1140 3054 -1132
rect 3061 -1134 3088 -1132
rect 3097 -1134 3318 -1124
rect 3061 -1144 3318 -1134
rect 3347 -1132 3397 -1124
rect 3347 -1141 3363 -1132
rect 2956 -1152 3007 -1144
rect 3054 -1152 3318 -1144
rect 3344 -1144 3363 -1141
rect 3370 -1144 3397 -1132
rect 3344 -1152 3397 -1144
rect 2972 -1160 2973 -1152
rect 2988 -1160 3001 -1152
rect 2972 -1168 2988 -1160
rect 2969 -1175 2988 -1172
rect 2969 -1184 2991 -1175
rect 2942 -1194 2991 -1184
rect 2942 -1200 2972 -1194
rect 2991 -1199 2996 -1194
rect 2914 -1216 2988 -1200
rect 3006 -1208 3036 -1152
rect 3071 -1162 3279 -1152
rect 3314 -1156 3359 -1152
rect 3362 -1153 3363 -1152
rect 3378 -1153 3391 -1152
rect 3097 -1192 3286 -1162
rect 3112 -1195 3286 -1192
rect 3105 -1198 3286 -1195
rect 2914 -1218 2927 -1216
rect 2942 -1218 2976 -1216
rect 2914 -1234 2988 -1218
rect 3015 -1222 3028 -1208
rect 3043 -1222 3059 -1206
rect 3105 -1211 3116 -1198
rect 2898 -1256 2899 -1240
rect 2914 -1256 2927 -1234
rect 2942 -1256 2972 -1234
rect 3015 -1238 3077 -1222
rect 3105 -1229 3116 -1213
rect 3121 -1218 3131 -1198
rect 3141 -1218 3155 -1198
rect 3158 -1211 3167 -1198
rect 3183 -1211 3192 -1198
rect 3121 -1229 3155 -1218
rect 3158 -1229 3167 -1213
rect 3183 -1229 3192 -1213
rect 3199 -1218 3209 -1198
rect 3219 -1218 3233 -1198
rect 3234 -1211 3245 -1198
rect 3199 -1229 3233 -1218
rect 3234 -1229 3245 -1213
rect 3291 -1222 3307 -1206
rect 3314 -1208 3344 -1156
rect 3378 -1160 3379 -1153
rect 3363 -1168 3379 -1160
rect 3350 -1200 3363 -1181
rect 3378 -1200 3408 -1184
rect 3350 -1216 3424 -1200
rect 3350 -1218 3363 -1216
rect 3378 -1218 3412 -1216
rect 3015 -1240 3028 -1238
rect 3043 -1240 3077 -1238
rect 3015 -1256 3077 -1240
rect 3121 -1245 3137 -1242
rect 3199 -1245 3229 -1234
rect 3277 -1238 3323 -1222
rect 3350 -1234 3424 -1218
rect 3277 -1240 3311 -1238
rect 3276 -1256 3323 -1240
rect 3350 -1256 3363 -1234
rect 3378 -1256 3408 -1234
rect 3435 -1256 3436 -1240
rect 3451 -1256 3464 -1096
rect 3494 -1200 3507 -1096
rect 3552 -1118 3553 -1108
rect 3568 -1118 3581 -1108
rect 3552 -1122 3581 -1118
rect 3586 -1122 3616 -1096
rect 3634 -1110 3650 -1108
rect 3722 -1110 3775 -1096
rect 3723 -1112 3787 -1110
rect 3830 -1112 3845 -1096
rect 3894 -1099 3924 -1096
rect 3894 -1102 3930 -1099
rect 3860 -1110 3876 -1108
rect 3634 -1122 3649 -1118
rect 3552 -1124 3649 -1122
rect 3677 -1124 3845 -1112
rect 3861 -1122 3876 -1118
rect 3894 -1121 3933 -1102
rect 3952 -1108 3959 -1107
rect 3958 -1115 3959 -1108
rect 3942 -1118 3943 -1115
rect 3958 -1118 3971 -1115
rect 3894 -1122 3924 -1121
rect 3933 -1122 3939 -1121
rect 3942 -1122 3971 -1118
rect 3861 -1123 3971 -1122
rect 3861 -1124 3977 -1123
rect 3536 -1132 3587 -1124
rect 3536 -1144 3561 -1132
rect 3568 -1144 3587 -1132
rect 3618 -1132 3668 -1124
rect 3618 -1140 3634 -1132
rect 3641 -1134 3668 -1132
rect 3677 -1134 3898 -1124
rect 3641 -1144 3898 -1134
rect 3927 -1132 3977 -1124
rect 3927 -1141 3943 -1132
rect 3536 -1152 3587 -1144
rect 3634 -1152 3898 -1144
rect 3924 -1144 3943 -1141
rect 3950 -1144 3977 -1132
rect 3924 -1152 3977 -1144
rect 3552 -1160 3553 -1152
rect 3568 -1160 3581 -1152
rect 3552 -1168 3568 -1160
rect 3549 -1175 3568 -1172
rect 3549 -1184 3571 -1175
rect 3522 -1194 3571 -1184
rect 3522 -1200 3552 -1194
rect 3571 -1199 3576 -1194
rect 3494 -1216 3568 -1200
rect 3586 -1208 3616 -1152
rect 3651 -1162 3859 -1152
rect 3894 -1156 3939 -1152
rect 3942 -1153 3943 -1152
rect 3958 -1153 3971 -1152
rect 3677 -1192 3866 -1162
rect 3692 -1195 3866 -1192
rect 3685 -1198 3866 -1195
rect 3494 -1218 3507 -1216
rect 3522 -1218 3556 -1216
rect 3494 -1234 3568 -1218
rect 3595 -1222 3608 -1208
rect 3623 -1222 3639 -1206
rect 3685 -1211 3696 -1198
rect 3478 -1256 3479 -1240
rect 3494 -1256 3507 -1234
rect 3522 -1256 3552 -1234
rect 3595 -1238 3657 -1222
rect 3685 -1229 3696 -1213
rect 3701 -1218 3711 -1198
rect 3721 -1218 3735 -1198
rect 3738 -1211 3747 -1198
rect 3763 -1211 3772 -1198
rect 3701 -1229 3735 -1218
rect 3738 -1229 3747 -1213
rect 3763 -1229 3772 -1213
rect 3779 -1218 3789 -1198
rect 3799 -1218 3813 -1198
rect 3814 -1211 3825 -1198
rect 3779 -1229 3813 -1218
rect 3814 -1229 3825 -1213
rect 3871 -1222 3887 -1206
rect 3894 -1208 3924 -1156
rect 3958 -1160 3959 -1153
rect 3943 -1168 3959 -1160
rect 3930 -1200 3943 -1181
rect 3958 -1200 3988 -1184
rect 3930 -1216 4004 -1200
rect 3930 -1218 3943 -1216
rect 3958 -1218 3992 -1216
rect 3595 -1240 3608 -1238
rect 3623 -1240 3657 -1238
rect 3595 -1256 3657 -1240
rect 3701 -1245 3717 -1242
rect 3779 -1245 3809 -1234
rect 3857 -1238 3903 -1222
rect 3930 -1234 4004 -1218
rect 3857 -1240 3891 -1238
rect 3856 -1256 3903 -1240
rect 3930 -1256 3943 -1234
rect 3958 -1256 3988 -1234
rect 4015 -1256 4016 -1240
rect 4031 -1256 4044 -1096
rect 4074 -1200 4087 -1096
rect 4132 -1118 4133 -1108
rect 4148 -1118 4161 -1108
rect 4132 -1122 4161 -1118
rect 4166 -1122 4196 -1096
rect 4214 -1110 4230 -1108
rect 4302 -1110 4355 -1096
rect 4303 -1112 4367 -1110
rect 4410 -1112 4425 -1096
rect 4474 -1099 4504 -1096
rect 4611 -1097 6944 -1096
rect 4474 -1102 4510 -1099
rect 4440 -1110 4456 -1108
rect 4214 -1122 4229 -1118
rect 4132 -1124 4229 -1122
rect 4257 -1124 4425 -1112
rect 4441 -1122 4456 -1118
rect 4474 -1121 4513 -1102
rect 4532 -1108 4539 -1107
rect 4538 -1115 4539 -1108
rect 4522 -1118 4523 -1115
rect 4538 -1118 4551 -1115
rect 4474 -1122 4504 -1121
rect 4513 -1122 4519 -1121
rect 4522 -1122 4551 -1118
rect 4441 -1123 4551 -1122
rect 4441 -1124 4557 -1123
rect 4116 -1132 4167 -1124
rect 4116 -1144 4141 -1132
rect 4148 -1144 4167 -1132
rect 4198 -1132 4248 -1124
rect 4198 -1140 4214 -1132
rect 4221 -1134 4248 -1132
rect 4257 -1134 4478 -1124
rect 4221 -1144 4478 -1134
rect 4507 -1132 4557 -1124
rect 4507 -1141 4523 -1132
rect 4116 -1152 4167 -1144
rect 4214 -1152 4478 -1144
rect 4504 -1144 4523 -1141
rect 4530 -1144 4557 -1132
rect 4504 -1152 4557 -1144
rect 4132 -1160 4133 -1152
rect 4148 -1160 4161 -1152
rect 4132 -1168 4148 -1160
rect 4129 -1175 4148 -1172
rect 4129 -1184 4151 -1175
rect 4102 -1194 4151 -1184
rect 4102 -1200 4132 -1194
rect 4151 -1199 4156 -1194
rect 4074 -1216 4148 -1200
rect 4166 -1208 4196 -1152
rect 4231 -1162 4439 -1152
rect 4474 -1156 4519 -1152
rect 4522 -1153 4523 -1152
rect 4538 -1153 4551 -1152
rect 4257 -1192 4446 -1162
rect 4272 -1195 4446 -1192
rect 4265 -1198 4446 -1195
rect 4074 -1218 4087 -1216
rect 4102 -1218 4136 -1216
rect 4074 -1234 4148 -1218
rect 4175 -1222 4188 -1208
rect 4203 -1222 4219 -1206
rect 4265 -1211 4276 -1198
rect 4058 -1256 4059 -1240
rect 4074 -1256 4087 -1234
rect 4102 -1256 4132 -1234
rect 4175 -1238 4237 -1222
rect 4265 -1229 4276 -1213
rect 4281 -1218 4291 -1198
rect 4301 -1218 4315 -1198
rect 4318 -1211 4327 -1198
rect 4343 -1211 4352 -1198
rect 4281 -1229 4315 -1218
rect 4318 -1229 4327 -1213
rect 4343 -1229 4352 -1213
rect 4359 -1218 4369 -1198
rect 4379 -1218 4393 -1198
rect 4394 -1211 4405 -1198
rect 4359 -1229 4393 -1218
rect 4394 -1229 4405 -1213
rect 4451 -1222 4467 -1206
rect 4474 -1208 4504 -1156
rect 4538 -1160 4539 -1153
rect 4523 -1168 4539 -1160
rect 4510 -1200 4523 -1181
rect 4538 -1200 4568 -1184
rect 4510 -1216 4584 -1200
rect 4510 -1218 4523 -1216
rect 4538 -1218 4572 -1216
rect 4175 -1240 4188 -1238
rect 4203 -1240 4237 -1238
rect 4175 -1256 4237 -1240
rect 4281 -1245 4297 -1242
rect 4359 -1245 4389 -1234
rect 4437 -1238 4483 -1222
rect 4510 -1234 4584 -1218
rect 4437 -1240 4471 -1238
rect 4436 -1256 4483 -1240
rect 4510 -1256 4523 -1234
rect 4538 -1256 4568 -1234
rect 4595 -1256 4596 -1240
rect 4611 -1256 4624 -1097
rect 4654 -1201 4667 -1097
rect 4712 -1119 4713 -1109
rect 4733 -1111 4741 -1109
rect 4731 -1113 4741 -1111
rect 4729 -1115 4741 -1113
rect 4728 -1119 4741 -1115
rect 4712 -1123 4741 -1119
rect 4746 -1123 4776 -1097
rect 4794 -1111 4810 -1109
rect 4882 -1111 4933 -1097
rect 4883 -1113 4947 -1111
rect 4990 -1113 5005 -1097
rect 5054 -1100 5084 -1097
rect 5054 -1103 5090 -1100
rect 5020 -1111 5036 -1109
rect 4794 -1123 4809 -1119
rect 4712 -1125 4809 -1123
rect 4837 -1125 5005 -1113
rect 5021 -1123 5036 -1119
rect 5054 -1122 5093 -1103
rect 5112 -1109 5119 -1108
rect 5118 -1116 5119 -1109
rect 5102 -1119 5103 -1116
rect 5118 -1119 5131 -1116
rect 5054 -1123 5084 -1122
rect 5093 -1123 5099 -1122
rect 5102 -1123 5131 -1119
rect 5021 -1124 5131 -1123
rect 5021 -1125 5137 -1124
rect 4696 -1133 4747 -1125
rect 4696 -1145 4721 -1133
rect 4728 -1145 4747 -1133
rect 4778 -1133 4828 -1125
rect 4778 -1141 4794 -1133
rect 4801 -1135 4828 -1133
rect 4837 -1135 5058 -1125
rect 4801 -1145 5058 -1135
rect 5087 -1133 5137 -1125
rect 5087 -1142 5103 -1133
rect 4696 -1153 4747 -1145
rect 4794 -1153 5058 -1145
rect 5084 -1145 5103 -1142
rect 5110 -1145 5137 -1133
rect 5084 -1153 5137 -1145
rect 4712 -1161 4713 -1153
rect 4728 -1161 4741 -1153
rect 4712 -1169 4728 -1161
rect 4709 -1176 4728 -1173
rect 4709 -1185 4731 -1176
rect 4682 -1195 4731 -1185
rect 4682 -1201 4712 -1195
rect 4731 -1200 4736 -1195
rect 4654 -1217 4728 -1201
rect 4746 -1209 4776 -1153
rect 4811 -1163 5019 -1153
rect 5054 -1157 5099 -1153
rect 5102 -1154 5103 -1153
rect 5118 -1154 5131 -1153
rect 4837 -1193 5026 -1163
rect 4852 -1196 5026 -1193
rect 4845 -1199 5026 -1196
rect 4654 -1219 4667 -1217
rect 4682 -1219 4716 -1217
rect 4654 -1235 4728 -1219
rect 4755 -1223 4768 -1209
rect 4783 -1223 4799 -1207
rect 4845 -1212 4856 -1199
rect 0 -1264 33 -1256
rect 0 -1290 7 -1264
rect 14 -1290 33 -1264
rect 97 -1268 159 -1256
rect 171 -1268 246 -1256
rect 304 -1268 379 -1256
rect 391 -1268 422 -1256
rect 428 -1268 463 -1256
rect 97 -1270 259 -1268
rect 0 -1298 33 -1290
rect 115 -1294 128 -1270
rect 143 -1272 158 -1270
rect 14 -1308 27 -1298
rect 42 -1308 72 -1294
rect 115 -1308 158 -1294
rect 182 -1297 189 -1290
rect 192 -1294 259 -1270
rect 291 -1270 463 -1268
rect 261 -1292 289 -1288
rect 291 -1292 371 -1270
rect 392 -1272 407 -1270
rect 261 -1294 371 -1292
rect 192 -1298 371 -1294
rect 165 -1308 195 -1298
rect 197 -1308 350 -1298
rect 358 -1308 388 -1298
rect 392 -1308 422 -1294
rect 450 -1308 463 -1270
rect 535 -1264 570 -1256
rect 535 -1290 536 -1264
rect 543 -1290 570 -1264
rect 478 -1308 508 -1294
rect 535 -1298 570 -1290
rect 572 -1264 613 -1256
rect 572 -1290 587 -1264
rect 594 -1290 613 -1264
rect 677 -1268 739 -1256
rect 751 -1268 826 -1256
rect 884 -1268 959 -1256
rect 971 -1268 1002 -1256
rect 1008 -1268 1043 -1256
rect 677 -1270 839 -1268
rect 572 -1298 613 -1290
rect 695 -1294 708 -1270
rect 723 -1272 738 -1270
rect 535 -1308 536 -1298
rect 551 -1308 564 -1298
rect 578 -1308 579 -1298
rect 594 -1308 607 -1298
rect 622 -1308 652 -1294
rect 695 -1308 738 -1294
rect 762 -1297 769 -1290
rect 772 -1294 839 -1270
rect 871 -1270 1043 -1268
rect 841 -1292 869 -1288
rect 871 -1292 951 -1270
rect 972 -1272 987 -1270
rect 841 -1294 951 -1292
rect 772 -1298 951 -1294
rect 745 -1308 775 -1298
rect 777 -1308 930 -1298
rect 938 -1308 968 -1298
rect 972 -1308 1002 -1294
rect 1030 -1308 1043 -1270
rect 1115 -1264 1150 -1256
rect 1115 -1290 1116 -1264
rect 1123 -1290 1150 -1264
rect 1058 -1308 1088 -1294
rect 1115 -1298 1150 -1290
rect 1152 -1264 1193 -1256
rect 1152 -1290 1167 -1264
rect 1174 -1290 1193 -1264
rect 1257 -1268 1319 -1256
rect 1331 -1268 1406 -1256
rect 1464 -1268 1539 -1256
rect 1551 -1268 1582 -1256
rect 1588 -1268 1623 -1256
rect 1257 -1270 1419 -1268
rect 1152 -1298 1193 -1290
rect 1275 -1294 1288 -1270
rect 1303 -1272 1318 -1270
rect 1115 -1308 1116 -1298
rect 1131 -1308 1144 -1298
rect 1158 -1308 1159 -1298
rect 1174 -1308 1187 -1298
rect 1202 -1308 1232 -1294
rect 1275 -1308 1318 -1294
rect 1342 -1297 1349 -1290
rect 1352 -1294 1419 -1270
rect 1451 -1270 1623 -1268
rect 1421 -1292 1449 -1288
rect 1451 -1292 1531 -1270
rect 1552 -1272 1567 -1270
rect 1421 -1294 1531 -1292
rect 1352 -1298 1531 -1294
rect 1325 -1308 1355 -1298
rect 1357 -1308 1510 -1298
rect 1518 -1308 1548 -1298
rect 1552 -1308 1582 -1294
rect 1610 -1308 1623 -1270
rect 1695 -1264 1730 -1256
rect 1695 -1290 1696 -1264
rect 1703 -1290 1730 -1264
rect 1638 -1308 1668 -1294
rect 1695 -1298 1730 -1290
rect 1732 -1264 1773 -1256
rect 1732 -1290 1747 -1264
rect 1754 -1290 1773 -1264
rect 1837 -1268 1899 -1256
rect 1911 -1268 1986 -1256
rect 2044 -1268 2119 -1256
rect 2131 -1268 2162 -1256
rect 2168 -1268 2203 -1256
rect 1837 -1270 1999 -1268
rect 1732 -1298 1773 -1290
rect 1855 -1294 1868 -1270
rect 1883 -1272 1898 -1270
rect 1695 -1308 1696 -1298
rect 1711 -1308 1724 -1298
rect 1738 -1308 1739 -1298
rect 1754 -1308 1767 -1298
rect 1782 -1308 1812 -1294
rect 1855 -1308 1898 -1294
rect 1922 -1297 1929 -1290
rect 1932 -1294 1999 -1270
rect 2031 -1270 2203 -1268
rect 2001 -1292 2029 -1288
rect 2031 -1292 2111 -1270
rect 2132 -1272 2147 -1270
rect 2001 -1294 2111 -1292
rect 1932 -1298 2111 -1294
rect 1905 -1308 1935 -1298
rect 1937 -1308 2090 -1298
rect 2098 -1308 2128 -1298
rect 2132 -1308 2162 -1294
rect 2190 -1308 2203 -1270
rect 2275 -1264 2310 -1256
rect 2275 -1290 2276 -1264
rect 2283 -1290 2310 -1264
rect 2218 -1308 2248 -1294
rect 2275 -1298 2310 -1290
rect 2312 -1264 2353 -1256
rect 2312 -1290 2327 -1264
rect 2334 -1290 2353 -1264
rect 2417 -1268 2479 -1256
rect 2491 -1268 2566 -1256
rect 2624 -1268 2699 -1256
rect 2711 -1268 2742 -1256
rect 2748 -1268 2783 -1256
rect 2417 -1270 2579 -1268
rect 2312 -1298 2353 -1290
rect 2435 -1294 2448 -1270
rect 2463 -1272 2478 -1270
rect 2275 -1308 2276 -1298
rect 2291 -1308 2304 -1298
rect 2318 -1308 2319 -1298
rect 2334 -1308 2347 -1298
rect 2362 -1308 2392 -1294
rect 2435 -1308 2478 -1294
rect 2502 -1297 2509 -1290
rect 2512 -1294 2579 -1270
rect 2611 -1270 2783 -1268
rect 2581 -1292 2609 -1288
rect 2611 -1292 2691 -1270
rect 2712 -1272 2727 -1270
rect 2581 -1294 2691 -1292
rect 2512 -1298 2691 -1294
rect 2485 -1308 2515 -1298
rect 2517 -1308 2670 -1298
rect 2678 -1308 2708 -1298
rect 2712 -1308 2742 -1294
rect 2770 -1308 2783 -1270
rect 2855 -1264 2890 -1256
rect 2855 -1290 2856 -1264
rect 2863 -1290 2890 -1264
rect 2798 -1308 2828 -1294
rect 2855 -1298 2890 -1290
rect 2892 -1264 2933 -1256
rect 2892 -1290 2907 -1264
rect 2914 -1290 2933 -1264
rect 2997 -1268 3059 -1256
rect 3071 -1268 3146 -1256
rect 3204 -1268 3279 -1256
rect 3291 -1268 3322 -1256
rect 3328 -1268 3363 -1256
rect 2997 -1270 3159 -1268
rect 2892 -1298 2933 -1290
rect 3015 -1294 3028 -1270
rect 3043 -1272 3058 -1270
rect 2855 -1308 2856 -1298
rect 2871 -1308 2884 -1298
rect 2898 -1308 2899 -1298
rect 2914 -1308 2927 -1298
rect 2942 -1308 2972 -1294
rect 3015 -1308 3058 -1294
rect 3082 -1297 3089 -1290
rect 3092 -1294 3159 -1270
rect 3191 -1270 3363 -1268
rect 3161 -1292 3189 -1288
rect 3191 -1292 3271 -1270
rect 3292 -1272 3307 -1270
rect 3161 -1294 3271 -1292
rect 3092 -1298 3271 -1294
rect 3065 -1308 3095 -1298
rect 3097 -1308 3250 -1298
rect 3258 -1308 3288 -1298
rect 3292 -1308 3322 -1294
rect 3350 -1308 3363 -1270
rect 3435 -1264 3470 -1256
rect 3435 -1290 3436 -1264
rect 3443 -1290 3470 -1264
rect 3378 -1308 3408 -1294
rect 3435 -1298 3470 -1290
rect 3472 -1264 3513 -1256
rect 3472 -1290 3487 -1264
rect 3494 -1290 3513 -1264
rect 3577 -1268 3639 -1256
rect 3651 -1268 3726 -1256
rect 3784 -1268 3859 -1256
rect 3871 -1268 3902 -1256
rect 3908 -1268 3943 -1256
rect 3577 -1270 3739 -1268
rect 3472 -1298 3513 -1290
rect 3595 -1294 3608 -1270
rect 3623 -1272 3638 -1270
rect 3435 -1308 3436 -1298
rect 3451 -1308 3464 -1298
rect 3478 -1308 3479 -1298
rect 3494 -1308 3507 -1298
rect 3522 -1308 3552 -1294
rect 3595 -1308 3638 -1294
rect 3662 -1297 3669 -1290
rect 3672 -1294 3739 -1270
rect 3771 -1270 3943 -1268
rect 3741 -1292 3769 -1288
rect 3771 -1292 3851 -1270
rect 3872 -1272 3887 -1270
rect 3741 -1294 3851 -1292
rect 3672 -1298 3851 -1294
rect 3645 -1308 3675 -1298
rect 3677 -1308 3830 -1298
rect 3838 -1308 3868 -1298
rect 3872 -1308 3902 -1294
rect 3930 -1308 3943 -1270
rect 4015 -1264 4050 -1256
rect 4015 -1290 4016 -1264
rect 4023 -1290 4050 -1264
rect 3958 -1308 3988 -1294
rect 4015 -1298 4050 -1290
rect 4052 -1264 4093 -1256
rect 4052 -1290 4067 -1264
rect 4074 -1290 4093 -1264
rect 4157 -1268 4219 -1256
rect 4231 -1268 4306 -1256
rect 4364 -1268 4439 -1256
rect 4451 -1268 4482 -1256
rect 4488 -1268 4523 -1256
rect 4157 -1270 4319 -1268
rect 4052 -1298 4093 -1290
rect 4175 -1294 4188 -1270
rect 4203 -1272 4218 -1270
rect 4015 -1308 4016 -1298
rect 4031 -1308 4044 -1298
rect 4058 -1308 4059 -1298
rect 4074 -1308 4087 -1298
rect 4102 -1308 4132 -1294
rect 4175 -1308 4218 -1294
rect 4242 -1297 4249 -1290
rect 4252 -1294 4319 -1270
rect 4351 -1270 4523 -1268
rect 4321 -1292 4349 -1288
rect 4351 -1292 4431 -1270
rect 4452 -1272 4467 -1270
rect 4321 -1294 4431 -1292
rect 4252 -1298 4431 -1294
rect 4225 -1308 4255 -1298
rect 4257 -1308 4410 -1298
rect 4418 -1308 4448 -1298
rect 4452 -1308 4482 -1294
rect 4510 -1308 4523 -1270
rect 4595 -1264 4630 -1256
rect 4638 -1257 4639 -1241
rect 4654 -1257 4667 -1235
rect 4682 -1257 4712 -1235
rect 4755 -1239 4817 -1223
rect 4845 -1230 4856 -1214
rect 4861 -1219 4871 -1199
rect 4881 -1219 4895 -1199
rect 4898 -1212 4907 -1199
rect 4923 -1212 4932 -1199
rect 4861 -1230 4895 -1219
rect 4898 -1230 4907 -1214
rect 4923 -1230 4932 -1214
rect 4939 -1219 4949 -1199
rect 4959 -1219 4973 -1199
rect 4974 -1212 4985 -1199
rect 4939 -1230 4973 -1219
rect 4974 -1230 4985 -1214
rect 5031 -1223 5047 -1207
rect 5054 -1209 5084 -1157
rect 5118 -1161 5119 -1154
rect 5103 -1169 5119 -1161
rect 5090 -1201 5103 -1182
rect 5118 -1201 5148 -1185
rect 5090 -1217 5164 -1201
rect 5090 -1219 5103 -1217
rect 5118 -1219 5152 -1217
rect 4755 -1241 4768 -1239
rect 4783 -1241 4817 -1239
rect 4755 -1257 4817 -1241
rect 4861 -1246 4877 -1243
rect 4939 -1246 4969 -1235
rect 5017 -1239 5063 -1223
rect 5090 -1235 5164 -1219
rect 5017 -1241 5051 -1239
rect 5016 -1257 5063 -1241
rect 5090 -1257 5103 -1235
rect 5118 -1257 5148 -1235
rect 5175 -1257 5176 -1241
rect 5191 -1257 5204 -1097
rect 5234 -1201 5247 -1097
rect 5292 -1119 5293 -1109
rect 5313 -1111 5321 -1109
rect 5311 -1113 5321 -1111
rect 5309 -1115 5321 -1113
rect 5308 -1119 5321 -1115
rect 5292 -1123 5321 -1119
rect 5326 -1123 5356 -1097
rect 5374 -1111 5390 -1109
rect 5462 -1111 5513 -1097
rect 5463 -1113 5527 -1111
rect 5570 -1113 5585 -1097
rect 5634 -1100 5664 -1097
rect 5634 -1103 5670 -1100
rect 5600 -1111 5616 -1109
rect 5374 -1123 5389 -1119
rect 5292 -1125 5389 -1123
rect 5417 -1125 5585 -1113
rect 5601 -1123 5616 -1119
rect 5634 -1122 5673 -1103
rect 5692 -1109 5699 -1108
rect 5698 -1116 5699 -1109
rect 5682 -1119 5683 -1116
rect 5698 -1119 5711 -1116
rect 5634 -1123 5664 -1122
rect 5673 -1123 5679 -1122
rect 5682 -1123 5711 -1119
rect 5601 -1124 5711 -1123
rect 5601 -1125 5717 -1124
rect 5276 -1133 5327 -1125
rect 5276 -1145 5301 -1133
rect 5308 -1145 5327 -1133
rect 5358 -1133 5408 -1125
rect 5358 -1141 5374 -1133
rect 5381 -1135 5408 -1133
rect 5417 -1135 5638 -1125
rect 5381 -1145 5638 -1135
rect 5667 -1133 5717 -1125
rect 5667 -1142 5683 -1133
rect 5276 -1153 5327 -1145
rect 5374 -1153 5638 -1145
rect 5664 -1145 5683 -1142
rect 5690 -1145 5717 -1133
rect 5664 -1153 5717 -1145
rect 5292 -1161 5293 -1153
rect 5308 -1161 5321 -1153
rect 5292 -1169 5308 -1161
rect 5289 -1176 5308 -1173
rect 5289 -1185 5311 -1176
rect 5262 -1195 5311 -1185
rect 5262 -1201 5292 -1195
rect 5311 -1200 5316 -1195
rect 5234 -1217 5308 -1201
rect 5326 -1209 5356 -1153
rect 5391 -1163 5599 -1153
rect 5634 -1157 5679 -1153
rect 5682 -1154 5683 -1153
rect 5698 -1154 5711 -1153
rect 5417 -1193 5606 -1163
rect 5432 -1196 5606 -1193
rect 5425 -1199 5606 -1196
rect 5234 -1219 5247 -1217
rect 5262 -1219 5296 -1217
rect 5234 -1235 5308 -1219
rect 5335 -1223 5348 -1209
rect 5363 -1223 5379 -1207
rect 5425 -1212 5436 -1199
rect 5218 -1257 5219 -1241
rect 5234 -1257 5247 -1235
rect 5262 -1257 5292 -1235
rect 5335 -1239 5397 -1223
rect 5425 -1230 5436 -1214
rect 5441 -1219 5451 -1199
rect 5461 -1219 5475 -1199
rect 5478 -1212 5487 -1199
rect 5503 -1212 5512 -1199
rect 5441 -1230 5475 -1219
rect 5478 -1230 5487 -1214
rect 5503 -1230 5512 -1214
rect 5519 -1219 5529 -1199
rect 5539 -1219 5553 -1199
rect 5554 -1212 5565 -1199
rect 5519 -1230 5553 -1219
rect 5554 -1230 5565 -1214
rect 5611 -1223 5627 -1207
rect 5634 -1209 5664 -1157
rect 5698 -1161 5699 -1154
rect 5683 -1169 5699 -1161
rect 5670 -1201 5683 -1182
rect 5698 -1201 5728 -1185
rect 5670 -1217 5744 -1201
rect 5670 -1219 5683 -1217
rect 5698 -1219 5732 -1217
rect 5335 -1241 5348 -1239
rect 5363 -1241 5397 -1239
rect 5335 -1257 5397 -1241
rect 5441 -1246 5457 -1243
rect 5519 -1246 5549 -1235
rect 5597 -1239 5643 -1223
rect 5670 -1235 5744 -1219
rect 5597 -1241 5631 -1239
rect 5596 -1257 5643 -1241
rect 5670 -1257 5683 -1235
rect 5698 -1257 5728 -1235
rect 5755 -1257 5756 -1241
rect 5771 -1257 5784 -1097
rect 5814 -1201 5827 -1097
rect 5872 -1119 5873 -1109
rect 5893 -1111 5901 -1109
rect 5891 -1113 5901 -1111
rect 5889 -1115 5901 -1113
rect 5888 -1119 5901 -1115
rect 5872 -1123 5901 -1119
rect 5906 -1123 5936 -1097
rect 5954 -1111 5970 -1109
rect 6042 -1111 6093 -1097
rect 6043 -1113 6107 -1111
rect 6150 -1113 6165 -1097
rect 6214 -1100 6244 -1097
rect 6214 -1103 6250 -1100
rect 6180 -1111 6196 -1109
rect 5954 -1123 5969 -1119
rect 5872 -1125 5969 -1123
rect 5997 -1125 6165 -1113
rect 6181 -1123 6196 -1119
rect 6214 -1122 6253 -1103
rect 6272 -1109 6279 -1108
rect 6278 -1116 6279 -1109
rect 6262 -1119 6263 -1116
rect 6278 -1119 6291 -1116
rect 6214 -1123 6244 -1122
rect 6253 -1123 6259 -1122
rect 6262 -1123 6291 -1119
rect 6181 -1124 6291 -1123
rect 6181 -1125 6297 -1124
rect 5856 -1133 5907 -1125
rect 5856 -1145 5881 -1133
rect 5888 -1145 5907 -1133
rect 5938 -1133 5988 -1125
rect 5938 -1141 5954 -1133
rect 5961 -1135 5988 -1133
rect 5997 -1135 6218 -1125
rect 5961 -1145 6218 -1135
rect 6247 -1133 6297 -1125
rect 6247 -1142 6263 -1133
rect 5856 -1153 5907 -1145
rect 5954 -1153 6218 -1145
rect 6244 -1145 6263 -1142
rect 6270 -1145 6297 -1133
rect 6244 -1153 6297 -1145
rect 5872 -1161 5873 -1153
rect 5888 -1161 5901 -1153
rect 5872 -1169 5888 -1161
rect 5869 -1176 5888 -1173
rect 5869 -1185 5891 -1176
rect 5842 -1195 5891 -1185
rect 5842 -1201 5872 -1195
rect 5891 -1200 5896 -1195
rect 5814 -1217 5888 -1201
rect 5906 -1209 5936 -1153
rect 5971 -1163 6179 -1153
rect 6214 -1157 6259 -1153
rect 6262 -1154 6263 -1153
rect 6278 -1154 6291 -1153
rect 5997 -1193 6186 -1163
rect 6012 -1196 6186 -1193
rect 6005 -1199 6186 -1196
rect 5814 -1219 5827 -1217
rect 5842 -1219 5876 -1217
rect 5814 -1235 5888 -1219
rect 5915 -1223 5928 -1209
rect 5943 -1223 5959 -1207
rect 6005 -1212 6016 -1199
rect 5798 -1257 5799 -1241
rect 5814 -1257 5827 -1235
rect 5842 -1257 5872 -1235
rect 5915 -1239 5977 -1223
rect 6005 -1230 6016 -1214
rect 6021 -1219 6031 -1199
rect 6041 -1219 6055 -1199
rect 6058 -1212 6067 -1199
rect 6083 -1212 6092 -1199
rect 6021 -1230 6055 -1219
rect 6058 -1230 6067 -1214
rect 6083 -1230 6092 -1214
rect 6099 -1219 6109 -1199
rect 6119 -1219 6133 -1199
rect 6134 -1212 6145 -1199
rect 6099 -1230 6133 -1219
rect 6134 -1230 6145 -1214
rect 6191 -1223 6207 -1207
rect 6214 -1209 6244 -1157
rect 6278 -1161 6279 -1154
rect 6263 -1169 6279 -1161
rect 6250 -1201 6263 -1182
rect 6278 -1201 6308 -1185
rect 6250 -1217 6324 -1201
rect 6250 -1219 6263 -1217
rect 6278 -1219 6312 -1217
rect 5915 -1241 5928 -1239
rect 5943 -1241 5977 -1239
rect 5915 -1257 5977 -1241
rect 6021 -1246 6037 -1243
rect 6099 -1246 6129 -1235
rect 6177 -1239 6223 -1223
rect 6250 -1235 6324 -1219
rect 6177 -1241 6211 -1239
rect 6176 -1257 6223 -1241
rect 6250 -1257 6263 -1235
rect 6278 -1257 6308 -1235
rect 6335 -1257 6336 -1241
rect 6351 -1257 6364 -1097
rect 6394 -1201 6407 -1097
rect 6452 -1119 6453 -1109
rect 6473 -1111 6481 -1109
rect 6471 -1113 6481 -1111
rect 6469 -1115 6481 -1113
rect 6468 -1119 6481 -1115
rect 6452 -1123 6481 -1119
rect 6486 -1123 6516 -1097
rect 6534 -1111 6550 -1109
rect 6622 -1111 6673 -1097
rect 6623 -1113 6687 -1111
rect 6730 -1113 6745 -1097
rect 6794 -1100 6824 -1097
rect 6794 -1103 6830 -1100
rect 6760 -1111 6776 -1109
rect 6534 -1123 6549 -1119
rect 6452 -1125 6549 -1123
rect 6577 -1125 6745 -1113
rect 6761 -1123 6776 -1119
rect 6794 -1122 6833 -1103
rect 6852 -1109 6859 -1108
rect 6858 -1116 6859 -1109
rect 6842 -1119 6843 -1116
rect 6858 -1119 6871 -1116
rect 6794 -1123 6824 -1122
rect 6833 -1123 6839 -1122
rect 6842 -1123 6871 -1119
rect 6761 -1124 6871 -1123
rect 6761 -1125 6877 -1124
rect 6436 -1133 6487 -1125
rect 6436 -1145 6461 -1133
rect 6468 -1145 6487 -1133
rect 6518 -1133 6568 -1125
rect 6518 -1141 6534 -1133
rect 6541 -1135 6568 -1133
rect 6577 -1135 6798 -1125
rect 6541 -1145 6798 -1135
rect 6827 -1133 6877 -1125
rect 6827 -1142 6843 -1133
rect 6436 -1153 6487 -1145
rect 6534 -1153 6798 -1145
rect 6824 -1145 6843 -1142
rect 6850 -1145 6877 -1133
rect 6824 -1153 6877 -1145
rect 6452 -1161 6453 -1153
rect 6468 -1161 6481 -1153
rect 6452 -1169 6468 -1161
rect 6449 -1176 6468 -1173
rect 6449 -1185 6471 -1176
rect 6422 -1195 6471 -1185
rect 6422 -1201 6452 -1195
rect 6471 -1200 6476 -1195
rect 6394 -1217 6468 -1201
rect 6486 -1209 6516 -1153
rect 6551 -1163 6759 -1153
rect 6794 -1157 6839 -1153
rect 6842 -1154 6843 -1153
rect 6858 -1154 6871 -1153
rect 6577 -1193 6766 -1163
rect 6592 -1196 6766 -1193
rect 6585 -1199 6766 -1196
rect 6394 -1219 6407 -1217
rect 6422 -1219 6456 -1217
rect 6394 -1235 6468 -1219
rect 6495 -1223 6508 -1209
rect 6523 -1223 6539 -1207
rect 6585 -1212 6596 -1199
rect 6378 -1257 6379 -1241
rect 6394 -1257 6407 -1235
rect 6422 -1257 6452 -1235
rect 6495 -1239 6557 -1223
rect 6585 -1230 6596 -1214
rect 6601 -1219 6611 -1199
rect 6621 -1219 6635 -1199
rect 6638 -1212 6647 -1199
rect 6663 -1212 6672 -1199
rect 6601 -1230 6635 -1219
rect 6638 -1230 6647 -1214
rect 6663 -1230 6672 -1214
rect 6679 -1219 6689 -1199
rect 6699 -1219 6713 -1199
rect 6714 -1212 6725 -1199
rect 6679 -1230 6713 -1219
rect 6714 -1230 6725 -1214
rect 6771 -1223 6787 -1207
rect 6794 -1209 6824 -1157
rect 6858 -1161 6859 -1154
rect 6843 -1169 6859 -1161
rect 6830 -1201 6843 -1182
rect 6858 -1201 6888 -1185
rect 6830 -1217 6904 -1201
rect 6830 -1219 6843 -1217
rect 6858 -1219 6892 -1217
rect 6495 -1241 6508 -1239
rect 6523 -1241 6557 -1239
rect 6495 -1257 6557 -1241
rect 6601 -1246 6617 -1243
rect 6679 -1246 6709 -1235
rect 6757 -1239 6803 -1223
rect 6830 -1235 6904 -1219
rect 6757 -1241 6791 -1239
rect 6756 -1257 6803 -1241
rect 6830 -1257 6843 -1235
rect 6858 -1257 6888 -1235
rect 6915 -1257 6916 -1241
rect 6931 -1257 6944 -1097
rect 4595 -1290 4596 -1264
rect 4603 -1290 4630 -1264
rect 4538 -1308 4568 -1294
rect 4595 -1298 4630 -1290
rect 4632 -1265 4673 -1257
rect 4632 -1291 4647 -1265
rect 4654 -1291 4673 -1265
rect 4737 -1269 4799 -1257
rect 4811 -1269 4886 -1257
rect 4944 -1269 5019 -1257
rect 5031 -1269 5062 -1257
rect 5068 -1269 5103 -1257
rect 4737 -1271 4899 -1269
rect 4595 -1308 4596 -1298
rect 4611 -1308 4624 -1298
rect 4632 -1299 4673 -1291
rect 4755 -1295 4768 -1271
rect 4783 -1273 4798 -1271
rect 4832 -1289 4899 -1271
rect 4931 -1271 5103 -1269
rect 4931 -1289 5011 -1271
rect 5032 -1273 5047 -1271
rect 0 -1309 4624 -1308
rect 4638 -1309 4639 -1299
rect 4654 -1309 4667 -1299
rect 4682 -1309 4712 -1295
rect 4755 -1309 4798 -1295
rect 4822 -1298 4829 -1291
rect 4832 -1299 5011 -1289
rect 4805 -1309 4835 -1299
rect 4837 -1309 4990 -1299
rect 4998 -1309 5028 -1299
rect 5032 -1309 5062 -1295
rect 5090 -1309 5103 -1271
rect 5175 -1265 5210 -1257
rect 5175 -1291 5176 -1265
rect 5183 -1291 5210 -1265
rect 5118 -1309 5148 -1295
rect 5175 -1299 5210 -1291
rect 5212 -1265 5253 -1257
rect 5212 -1291 5227 -1265
rect 5234 -1291 5253 -1265
rect 5317 -1269 5379 -1257
rect 5391 -1269 5466 -1257
rect 5524 -1269 5599 -1257
rect 5611 -1269 5642 -1257
rect 5648 -1269 5683 -1257
rect 5317 -1271 5479 -1269
rect 5212 -1299 5253 -1291
rect 5335 -1295 5348 -1271
rect 5363 -1273 5378 -1271
rect 5412 -1289 5479 -1271
rect 5511 -1271 5683 -1269
rect 5511 -1289 5591 -1271
rect 5612 -1273 5627 -1271
rect 5175 -1309 5176 -1299
rect 5191 -1309 5204 -1299
rect 5218 -1309 5219 -1299
rect 5234 -1309 5247 -1299
rect 5262 -1309 5292 -1295
rect 5335 -1309 5378 -1295
rect 5402 -1298 5409 -1291
rect 5412 -1299 5591 -1289
rect 5385 -1309 5415 -1299
rect 5417 -1309 5570 -1299
rect 5578 -1309 5608 -1299
rect 5612 -1309 5642 -1295
rect 5670 -1309 5683 -1271
rect 5755 -1265 5790 -1257
rect 5755 -1291 5756 -1265
rect 5763 -1291 5790 -1265
rect 5698 -1309 5728 -1295
rect 5755 -1299 5790 -1291
rect 5792 -1265 5833 -1257
rect 5792 -1291 5807 -1265
rect 5814 -1291 5833 -1265
rect 5897 -1269 5959 -1257
rect 5971 -1269 6046 -1257
rect 6104 -1269 6179 -1257
rect 6191 -1269 6222 -1257
rect 6228 -1269 6263 -1257
rect 5897 -1271 6059 -1269
rect 5792 -1299 5833 -1291
rect 5915 -1295 5928 -1271
rect 5943 -1273 5958 -1271
rect 5992 -1289 6059 -1271
rect 6091 -1271 6263 -1269
rect 6091 -1289 6171 -1271
rect 6192 -1273 6207 -1271
rect 5755 -1309 5756 -1299
rect 5771 -1309 5784 -1299
rect 5798 -1309 5799 -1299
rect 5814 -1309 5827 -1299
rect 5842 -1309 5872 -1295
rect 5915 -1309 5958 -1295
rect 5982 -1298 5989 -1291
rect 5992 -1299 6171 -1289
rect 5965 -1309 5995 -1299
rect 5997 -1309 6150 -1299
rect 6158 -1309 6188 -1299
rect 6192 -1309 6222 -1295
rect 6250 -1309 6263 -1271
rect 6335 -1265 6370 -1257
rect 6335 -1291 6336 -1265
rect 6343 -1291 6370 -1265
rect 6278 -1309 6308 -1295
rect 6335 -1299 6370 -1291
rect 6372 -1265 6413 -1257
rect 6372 -1291 6387 -1265
rect 6394 -1291 6413 -1265
rect 6477 -1269 6539 -1257
rect 6551 -1269 6626 -1257
rect 6684 -1269 6759 -1257
rect 6771 -1269 6802 -1257
rect 6808 -1269 6843 -1257
rect 6477 -1271 6639 -1269
rect 6372 -1299 6413 -1291
rect 6495 -1295 6508 -1271
rect 6523 -1273 6538 -1271
rect 6572 -1289 6639 -1271
rect 6671 -1271 6843 -1269
rect 6671 -1289 6751 -1271
rect 6772 -1273 6787 -1271
rect 6335 -1309 6336 -1299
rect 6351 -1309 6364 -1299
rect 6378 -1309 6379 -1299
rect 6394 -1309 6407 -1299
rect 6422 -1309 6452 -1295
rect 6495 -1309 6538 -1295
rect 6562 -1298 6569 -1291
rect 6572 -1299 6751 -1289
rect 6545 -1309 6575 -1299
rect 6577 -1309 6730 -1299
rect 6738 -1309 6768 -1299
rect 6772 -1309 6802 -1295
rect 6830 -1309 6843 -1271
rect 6915 -1265 6950 -1257
rect 6915 -1291 6916 -1265
rect 6923 -1291 6950 -1265
rect 6858 -1309 6888 -1295
rect 6915 -1299 6950 -1291
rect 6915 -1309 6916 -1299
rect 6931 -1309 6944 -1299
rect 0 -1322 6944 -1309
rect 14 -1352 27 -1322
rect 42 -1340 72 -1322
rect 115 -1336 129 -1322
rect 165 -1336 385 -1322
rect 116 -1338 129 -1336
rect 82 -1350 97 -1338
rect 79 -1352 101 -1350
rect 106 -1352 136 -1338
rect 197 -1340 350 -1336
rect 179 -1352 371 -1340
rect 414 -1352 444 -1338
rect 450 -1352 463 -1322
rect 478 -1340 508 -1322
rect 551 -1352 564 -1322
rect 594 -1352 607 -1322
rect 622 -1340 652 -1322
rect 695 -1336 709 -1322
rect 745 -1336 965 -1322
rect 696 -1338 709 -1336
rect 662 -1350 677 -1338
rect 659 -1352 681 -1350
rect 686 -1352 716 -1338
rect 777 -1340 930 -1336
rect 759 -1352 951 -1340
rect 994 -1352 1024 -1338
rect 1030 -1352 1043 -1322
rect 1058 -1340 1088 -1322
rect 1131 -1352 1144 -1322
rect 1174 -1352 1187 -1322
rect 1202 -1340 1232 -1322
rect 1275 -1336 1289 -1322
rect 1325 -1336 1545 -1322
rect 1276 -1338 1289 -1336
rect 1242 -1350 1257 -1338
rect 1239 -1352 1261 -1350
rect 1266 -1352 1296 -1338
rect 1357 -1340 1510 -1336
rect 1339 -1352 1531 -1340
rect 1574 -1352 1604 -1338
rect 1610 -1352 1623 -1322
rect 1638 -1340 1668 -1322
rect 1711 -1352 1724 -1322
rect 1754 -1352 1767 -1322
rect 1782 -1340 1812 -1322
rect 1855 -1336 1869 -1322
rect 1905 -1336 2125 -1322
rect 1856 -1338 1869 -1336
rect 1822 -1350 1837 -1338
rect 1819 -1352 1841 -1350
rect 1846 -1352 1876 -1338
rect 1937 -1340 2090 -1336
rect 1919 -1352 2111 -1340
rect 2154 -1352 2184 -1338
rect 2190 -1352 2203 -1322
rect 2218 -1340 2248 -1322
rect 2291 -1352 2304 -1322
rect 2334 -1352 2347 -1322
rect 2362 -1340 2392 -1322
rect 2435 -1336 2449 -1322
rect 2485 -1336 2705 -1322
rect 2436 -1338 2449 -1336
rect 2402 -1350 2417 -1338
rect 2399 -1352 2421 -1350
rect 2426 -1352 2456 -1338
rect 2517 -1340 2670 -1336
rect 2499 -1352 2691 -1340
rect 2734 -1352 2764 -1338
rect 2770 -1352 2783 -1322
rect 2798 -1340 2828 -1322
rect 2871 -1352 2884 -1322
rect 2914 -1352 2927 -1322
rect 2942 -1340 2972 -1322
rect 3015 -1336 3029 -1322
rect 3065 -1336 3285 -1322
rect 3016 -1338 3029 -1336
rect 2982 -1350 2997 -1338
rect 2979 -1352 3001 -1350
rect 3006 -1352 3036 -1338
rect 3097 -1340 3250 -1336
rect 3079 -1352 3271 -1340
rect 3314 -1352 3344 -1338
rect 3350 -1352 3363 -1322
rect 3378 -1340 3408 -1322
rect 3451 -1352 3464 -1322
rect 3494 -1352 3507 -1322
rect 3522 -1340 3552 -1322
rect 3595 -1336 3609 -1322
rect 3645 -1336 3865 -1322
rect 3596 -1338 3609 -1336
rect 3562 -1350 3577 -1338
rect 3559 -1352 3581 -1350
rect 3586 -1352 3616 -1338
rect 3677 -1340 3830 -1336
rect 3659 -1352 3851 -1340
rect 3894 -1352 3924 -1338
rect 3930 -1352 3943 -1322
rect 3958 -1340 3988 -1322
rect 4031 -1352 4044 -1322
rect 4074 -1352 4087 -1322
rect 4102 -1340 4132 -1322
rect 4175 -1336 4189 -1322
rect 4225 -1336 4445 -1322
rect 4176 -1338 4189 -1336
rect 4142 -1350 4157 -1338
rect 4139 -1352 4161 -1350
rect 4166 -1352 4196 -1338
rect 4257 -1340 4410 -1336
rect 4239 -1352 4431 -1340
rect 4474 -1352 4504 -1338
rect 4510 -1352 4523 -1322
rect 4538 -1340 4568 -1322
rect 4611 -1323 6944 -1322
rect 4611 -1352 4624 -1323
rect 0 -1353 4624 -1352
rect 4654 -1353 4667 -1323
rect 4682 -1341 4712 -1323
rect 4755 -1337 4769 -1323
rect 4805 -1337 5025 -1323
rect 4756 -1339 4769 -1337
rect 4722 -1351 4737 -1339
rect 4719 -1353 4741 -1351
rect 4746 -1353 4776 -1339
rect 4837 -1341 4990 -1337
rect 4819 -1353 5011 -1341
rect 5054 -1353 5084 -1339
rect 5090 -1353 5103 -1323
rect 5118 -1341 5148 -1323
rect 5191 -1353 5204 -1323
rect 5234 -1353 5247 -1323
rect 5262 -1341 5292 -1323
rect 5335 -1337 5349 -1323
rect 5385 -1337 5605 -1323
rect 5336 -1339 5349 -1337
rect 5302 -1351 5317 -1339
rect 5299 -1353 5321 -1351
rect 5326 -1353 5356 -1339
rect 5417 -1341 5570 -1337
rect 5399 -1353 5591 -1341
rect 5634 -1353 5664 -1339
rect 5670 -1353 5683 -1323
rect 5698 -1341 5728 -1323
rect 5771 -1353 5784 -1323
rect 5814 -1353 5827 -1323
rect 5842 -1341 5872 -1323
rect 5915 -1337 5929 -1323
rect 5965 -1337 6185 -1323
rect 5916 -1339 5929 -1337
rect 5882 -1351 5897 -1339
rect 5879 -1353 5901 -1351
rect 5906 -1353 5936 -1339
rect 5997 -1341 6150 -1337
rect 5979 -1353 6171 -1341
rect 6214 -1353 6244 -1339
rect 6250 -1353 6263 -1323
rect 6278 -1341 6308 -1323
rect 6351 -1353 6364 -1323
rect 6394 -1353 6407 -1323
rect 6422 -1341 6452 -1323
rect 6495 -1337 6509 -1323
rect 6545 -1337 6765 -1323
rect 6496 -1339 6509 -1337
rect 6462 -1351 6477 -1339
rect 6459 -1353 6481 -1351
rect 6486 -1353 6516 -1339
rect 6577 -1341 6730 -1337
rect 6559 -1353 6751 -1341
rect 6794 -1353 6824 -1339
rect 6830 -1353 6843 -1323
rect 6858 -1341 6888 -1323
rect 6931 -1353 6944 -1323
rect 0 -1366 6944 -1353
rect 14 -1470 27 -1366
rect 72 -1388 73 -1378
rect 88 -1388 101 -1378
rect 72 -1392 101 -1388
rect 106 -1392 136 -1366
rect 154 -1380 170 -1378
rect 242 -1380 295 -1366
rect 243 -1382 307 -1380
rect 350 -1382 365 -1366
rect 414 -1369 444 -1366
rect 414 -1372 450 -1369
rect 380 -1380 396 -1378
rect 154 -1392 169 -1388
rect 72 -1394 169 -1392
rect 197 -1394 365 -1382
rect 381 -1392 396 -1388
rect 414 -1391 453 -1372
rect 472 -1378 479 -1377
rect 478 -1385 479 -1378
rect 462 -1388 463 -1385
rect 478 -1388 491 -1385
rect 414 -1392 444 -1391
rect 453 -1392 459 -1391
rect 462 -1392 491 -1388
rect 381 -1393 491 -1392
rect 381 -1394 497 -1393
rect 56 -1402 107 -1394
rect 56 -1414 81 -1402
rect 88 -1414 107 -1402
rect 138 -1402 188 -1394
rect 138 -1410 154 -1402
rect 161 -1404 188 -1402
rect 197 -1404 418 -1394
rect 161 -1414 418 -1404
rect 447 -1402 497 -1394
rect 447 -1411 463 -1402
rect 56 -1422 107 -1414
rect 154 -1422 418 -1414
rect 444 -1414 463 -1411
rect 470 -1414 497 -1402
rect 444 -1422 497 -1414
rect 72 -1430 73 -1422
rect 88 -1430 101 -1422
rect 72 -1438 88 -1430
rect 69 -1445 88 -1442
rect 69 -1454 91 -1445
rect 42 -1464 91 -1454
rect 42 -1470 72 -1464
rect 91 -1469 96 -1464
rect 14 -1486 88 -1470
rect 106 -1478 136 -1422
rect 171 -1432 379 -1422
rect 414 -1426 459 -1422
rect 462 -1423 463 -1422
rect 478 -1423 491 -1422
rect 197 -1462 386 -1432
rect 212 -1465 386 -1462
rect 205 -1468 386 -1465
rect 14 -1488 27 -1486
rect 42 -1488 76 -1486
rect 14 -1504 88 -1488
rect 115 -1492 128 -1478
rect 143 -1492 159 -1476
rect 205 -1481 216 -1468
rect 14 -1526 27 -1504
rect 42 -1526 72 -1504
rect 115 -1508 177 -1492
rect 205 -1499 216 -1483
rect 221 -1488 231 -1468
rect 241 -1488 255 -1468
rect 258 -1481 267 -1468
rect 283 -1481 292 -1468
rect 221 -1499 255 -1488
rect 258 -1499 267 -1483
rect 283 -1499 292 -1483
rect 299 -1488 309 -1468
rect 319 -1488 333 -1468
rect 334 -1481 345 -1468
rect 299 -1499 333 -1488
rect 334 -1499 345 -1483
rect 391 -1492 407 -1476
rect 414 -1478 444 -1426
rect 478 -1430 479 -1423
rect 463 -1438 479 -1430
rect 450 -1470 463 -1451
rect 478 -1470 508 -1454
rect 450 -1486 524 -1470
rect 450 -1488 463 -1486
rect 478 -1488 512 -1486
rect 115 -1510 128 -1508
rect 143 -1510 177 -1508
rect 115 -1526 177 -1510
rect 221 -1515 237 -1512
rect 299 -1515 329 -1504
rect 377 -1508 423 -1492
rect 450 -1504 524 -1488
rect 377 -1510 411 -1508
rect 376 -1526 423 -1510
rect 450 -1526 463 -1504
rect 478 -1526 508 -1504
rect 535 -1526 536 -1510
rect 551 -1526 564 -1366
rect 594 -1470 607 -1366
rect 652 -1388 653 -1378
rect 668 -1388 681 -1378
rect 652 -1392 681 -1388
rect 686 -1392 716 -1366
rect 734 -1380 750 -1378
rect 822 -1380 875 -1366
rect 823 -1382 887 -1380
rect 930 -1382 945 -1366
rect 994 -1369 1024 -1366
rect 994 -1372 1030 -1369
rect 960 -1380 976 -1378
rect 734 -1392 749 -1388
rect 652 -1394 749 -1392
rect 777 -1394 945 -1382
rect 961 -1392 976 -1388
rect 994 -1391 1033 -1372
rect 1052 -1378 1059 -1377
rect 1058 -1385 1059 -1378
rect 1042 -1388 1043 -1385
rect 1058 -1388 1071 -1385
rect 994 -1392 1024 -1391
rect 1033 -1392 1039 -1391
rect 1042 -1392 1071 -1388
rect 961 -1393 1071 -1392
rect 961 -1394 1077 -1393
rect 636 -1402 687 -1394
rect 636 -1414 661 -1402
rect 668 -1414 687 -1402
rect 718 -1402 768 -1394
rect 718 -1410 734 -1402
rect 741 -1404 768 -1402
rect 777 -1404 998 -1394
rect 741 -1414 998 -1404
rect 1027 -1402 1077 -1394
rect 1027 -1411 1043 -1402
rect 636 -1422 687 -1414
rect 734 -1422 998 -1414
rect 1024 -1414 1043 -1411
rect 1050 -1414 1077 -1402
rect 1024 -1422 1077 -1414
rect 652 -1430 653 -1422
rect 668 -1430 681 -1422
rect 652 -1438 668 -1430
rect 649 -1445 668 -1442
rect 649 -1454 671 -1445
rect 622 -1464 671 -1454
rect 622 -1470 652 -1464
rect 671 -1469 676 -1464
rect 594 -1486 668 -1470
rect 686 -1478 716 -1422
rect 751 -1432 959 -1422
rect 994 -1426 1039 -1422
rect 1042 -1423 1043 -1422
rect 1058 -1423 1071 -1422
rect 777 -1462 966 -1432
rect 792 -1465 966 -1462
rect 785 -1468 966 -1465
rect 594 -1488 607 -1486
rect 622 -1488 656 -1486
rect 594 -1504 668 -1488
rect 695 -1492 708 -1478
rect 723 -1492 739 -1476
rect 785 -1481 796 -1468
rect 578 -1526 579 -1510
rect 594 -1526 607 -1504
rect 622 -1526 652 -1504
rect 695 -1508 757 -1492
rect 785 -1499 796 -1483
rect 801 -1488 811 -1468
rect 821 -1488 835 -1468
rect 838 -1481 847 -1468
rect 863 -1481 872 -1468
rect 801 -1499 835 -1488
rect 838 -1499 847 -1483
rect 863 -1499 872 -1483
rect 879 -1488 889 -1468
rect 899 -1488 913 -1468
rect 914 -1481 925 -1468
rect 879 -1499 913 -1488
rect 914 -1499 925 -1483
rect 971 -1492 987 -1476
rect 994 -1478 1024 -1426
rect 1058 -1430 1059 -1423
rect 1043 -1438 1059 -1430
rect 1030 -1470 1043 -1451
rect 1058 -1470 1088 -1454
rect 1030 -1486 1104 -1470
rect 1030 -1488 1043 -1486
rect 1058 -1488 1092 -1486
rect 695 -1510 708 -1508
rect 723 -1510 757 -1508
rect 695 -1526 757 -1510
rect 801 -1515 817 -1512
rect 879 -1515 909 -1504
rect 957 -1508 1003 -1492
rect 1030 -1504 1104 -1488
rect 957 -1510 991 -1508
rect 956 -1526 1003 -1510
rect 1030 -1526 1043 -1504
rect 1058 -1526 1088 -1504
rect 1115 -1526 1116 -1510
rect 1131 -1526 1144 -1366
rect 1174 -1470 1187 -1366
rect 1232 -1388 1233 -1378
rect 1248 -1388 1261 -1378
rect 1232 -1392 1261 -1388
rect 1266 -1392 1296 -1366
rect 1314 -1380 1330 -1378
rect 1402 -1380 1455 -1366
rect 1403 -1382 1467 -1380
rect 1510 -1382 1525 -1366
rect 1574 -1369 1604 -1366
rect 1574 -1372 1610 -1369
rect 1540 -1380 1556 -1378
rect 1314 -1392 1329 -1388
rect 1232 -1394 1329 -1392
rect 1357 -1394 1525 -1382
rect 1541 -1392 1556 -1388
rect 1574 -1391 1613 -1372
rect 1632 -1378 1639 -1377
rect 1638 -1385 1639 -1378
rect 1622 -1388 1623 -1385
rect 1638 -1388 1651 -1385
rect 1574 -1392 1604 -1391
rect 1613 -1392 1619 -1391
rect 1622 -1392 1651 -1388
rect 1541 -1393 1651 -1392
rect 1541 -1394 1657 -1393
rect 1216 -1402 1267 -1394
rect 1216 -1414 1241 -1402
rect 1248 -1414 1267 -1402
rect 1298 -1402 1348 -1394
rect 1298 -1410 1314 -1402
rect 1321 -1404 1348 -1402
rect 1357 -1404 1578 -1394
rect 1321 -1414 1578 -1404
rect 1607 -1402 1657 -1394
rect 1607 -1411 1623 -1402
rect 1216 -1422 1267 -1414
rect 1314 -1422 1578 -1414
rect 1604 -1414 1623 -1411
rect 1630 -1414 1657 -1402
rect 1604 -1422 1657 -1414
rect 1232 -1430 1233 -1422
rect 1248 -1430 1261 -1422
rect 1232 -1438 1248 -1430
rect 1229 -1445 1248 -1442
rect 1229 -1454 1251 -1445
rect 1202 -1464 1251 -1454
rect 1202 -1470 1232 -1464
rect 1251 -1469 1256 -1464
rect 1174 -1486 1248 -1470
rect 1266 -1478 1296 -1422
rect 1331 -1432 1539 -1422
rect 1574 -1426 1619 -1422
rect 1622 -1423 1623 -1422
rect 1638 -1423 1651 -1422
rect 1357 -1462 1546 -1432
rect 1372 -1465 1546 -1462
rect 1365 -1468 1546 -1465
rect 1174 -1488 1187 -1486
rect 1202 -1488 1236 -1486
rect 1174 -1504 1248 -1488
rect 1275 -1492 1288 -1478
rect 1303 -1492 1319 -1476
rect 1365 -1481 1376 -1468
rect 1158 -1526 1159 -1510
rect 1174 -1526 1187 -1504
rect 1202 -1526 1232 -1504
rect 1275 -1508 1337 -1492
rect 1365 -1499 1376 -1483
rect 1381 -1488 1391 -1468
rect 1401 -1488 1415 -1468
rect 1418 -1481 1427 -1468
rect 1443 -1481 1452 -1468
rect 1381 -1499 1415 -1488
rect 1418 -1499 1427 -1483
rect 1443 -1499 1452 -1483
rect 1459 -1488 1469 -1468
rect 1479 -1488 1493 -1468
rect 1494 -1481 1505 -1468
rect 1459 -1499 1493 -1488
rect 1494 -1499 1505 -1483
rect 1551 -1492 1567 -1476
rect 1574 -1478 1604 -1426
rect 1638 -1430 1639 -1423
rect 1623 -1438 1639 -1430
rect 1610 -1470 1623 -1451
rect 1638 -1470 1668 -1454
rect 1610 -1486 1684 -1470
rect 1610 -1488 1623 -1486
rect 1638 -1488 1672 -1486
rect 1275 -1510 1288 -1508
rect 1303 -1510 1337 -1508
rect 1275 -1526 1337 -1510
rect 1381 -1515 1397 -1512
rect 1459 -1515 1489 -1504
rect 1537 -1508 1583 -1492
rect 1610 -1504 1684 -1488
rect 1537 -1510 1571 -1508
rect 1536 -1526 1583 -1510
rect 1610 -1526 1623 -1504
rect 1638 -1526 1668 -1504
rect 1695 -1526 1696 -1510
rect 1711 -1526 1724 -1366
rect 1754 -1470 1767 -1366
rect 1812 -1388 1813 -1378
rect 1828 -1388 1841 -1378
rect 1812 -1392 1841 -1388
rect 1846 -1392 1876 -1366
rect 1894 -1380 1910 -1378
rect 1982 -1380 2035 -1366
rect 1983 -1382 2047 -1380
rect 2090 -1382 2105 -1366
rect 2154 -1369 2184 -1366
rect 2154 -1372 2190 -1369
rect 2120 -1380 2136 -1378
rect 1894 -1392 1909 -1388
rect 1812 -1394 1909 -1392
rect 1937 -1394 2105 -1382
rect 2121 -1392 2136 -1388
rect 2154 -1391 2193 -1372
rect 2212 -1378 2219 -1377
rect 2218 -1385 2219 -1378
rect 2202 -1388 2203 -1385
rect 2218 -1388 2231 -1385
rect 2154 -1392 2184 -1391
rect 2193 -1392 2199 -1391
rect 2202 -1392 2231 -1388
rect 2121 -1393 2231 -1392
rect 2121 -1394 2237 -1393
rect 1796 -1402 1847 -1394
rect 1796 -1414 1821 -1402
rect 1828 -1414 1847 -1402
rect 1878 -1402 1928 -1394
rect 1878 -1410 1894 -1402
rect 1901 -1404 1928 -1402
rect 1937 -1404 2158 -1394
rect 1901 -1414 2158 -1404
rect 2187 -1402 2237 -1394
rect 2187 -1411 2203 -1402
rect 1796 -1422 1847 -1414
rect 1894 -1422 2158 -1414
rect 2184 -1414 2203 -1411
rect 2210 -1414 2237 -1402
rect 2184 -1422 2237 -1414
rect 1812 -1430 1813 -1422
rect 1828 -1430 1841 -1422
rect 1812 -1438 1828 -1430
rect 1809 -1445 1828 -1442
rect 1809 -1454 1831 -1445
rect 1782 -1464 1831 -1454
rect 1782 -1470 1812 -1464
rect 1831 -1469 1836 -1464
rect 1754 -1486 1828 -1470
rect 1846 -1478 1876 -1422
rect 1911 -1432 2119 -1422
rect 2154 -1426 2199 -1422
rect 2202 -1423 2203 -1422
rect 2218 -1423 2231 -1422
rect 1937 -1462 2126 -1432
rect 1952 -1465 2126 -1462
rect 1945 -1468 2126 -1465
rect 1754 -1488 1767 -1486
rect 1782 -1488 1816 -1486
rect 1754 -1504 1828 -1488
rect 1855 -1492 1868 -1478
rect 1883 -1492 1899 -1476
rect 1945 -1481 1956 -1468
rect 1738 -1526 1739 -1510
rect 1754 -1526 1767 -1504
rect 1782 -1526 1812 -1504
rect 1855 -1508 1917 -1492
rect 1945 -1499 1956 -1483
rect 1961 -1488 1971 -1468
rect 1981 -1488 1995 -1468
rect 1998 -1481 2007 -1468
rect 2023 -1481 2032 -1468
rect 1961 -1499 1995 -1488
rect 1998 -1499 2007 -1483
rect 2023 -1499 2032 -1483
rect 2039 -1488 2049 -1468
rect 2059 -1488 2073 -1468
rect 2074 -1481 2085 -1468
rect 2039 -1499 2073 -1488
rect 2074 -1499 2085 -1483
rect 2131 -1492 2147 -1476
rect 2154 -1478 2184 -1426
rect 2218 -1430 2219 -1423
rect 2203 -1438 2219 -1430
rect 2190 -1470 2203 -1451
rect 2218 -1470 2248 -1454
rect 2190 -1486 2264 -1470
rect 2190 -1488 2203 -1486
rect 2218 -1488 2252 -1486
rect 1855 -1510 1868 -1508
rect 1883 -1510 1917 -1508
rect 1855 -1526 1917 -1510
rect 1961 -1515 1977 -1512
rect 2039 -1515 2069 -1504
rect 2117 -1508 2163 -1492
rect 2190 -1504 2264 -1488
rect 2117 -1510 2151 -1508
rect 2116 -1526 2163 -1510
rect 2190 -1526 2203 -1504
rect 2218 -1526 2248 -1504
rect 2275 -1526 2276 -1510
rect 2291 -1526 2304 -1366
rect 2334 -1470 2347 -1366
rect 2392 -1388 2393 -1378
rect 2408 -1388 2421 -1378
rect 2392 -1392 2421 -1388
rect 2426 -1392 2456 -1366
rect 2474 -1380 2490 -1378
rect 2562 -1380 2615 -1366
rect 2563 -1382 2627 -1380
rect 2670 -1382 2685 -1366
rect 2734 -1369 2764 -1366
rect 2734 -1372 2770 -1369
rect 2700 -1380 2716 -1378
rect 2474 -1392 2489 -1388
rect 2392 -1394 2489 -1392
rect 2517 -1394 2685 -1382
rect 2701 -1392 2716 -1388
rect 2734 -1391 2773 -1372
rect 2792 -1378 2799 -1377
rect 2798 -1385 2799 -1378
rect 2782 -1388 2783 -1385
rect 2798 -1388 2811 -1385
rect 2734 -1392 2764 -1391
rect 2773 -1392 2779 -1391
rect 2782 -1392 2811 -1388
rect 2701 -1393 2811 -1392
rect 2701 -1394 2817 -1393
rect 2376 -1402 2427 -1394
rect 2376 -1414 2401 -1402
rect 2408 -1414 2427 -1402
rect 2458 -1402 2508 -1394
rect 2458 -1410 2474 -1402
rect 2481 -1404 2508 -1402
rect 2517 -1404 2738 -1394
rect 2481 -1414 2738 -1404
rect 2767 -1402 2817 -1394
rect 2767 -1411 2783 -1402
rect 2376 -1422 2427 -1414
rect 2474 -1422 2738 -1414
rect 2764 -1414 2783 -1411
rect 2790 -1414 2817 -1402
rect 2764 -1422 2817 -1414
rect 2392 -1430 2393 -1422
rect 2408 -1430 2421 -1422
rect 2392 -1438 2408 -1430
rect 2389 -1445 2408 -1442
rect 2389 -1454 2411 -1445
rect 2362 -1464 2411 -1454
rect 2362 -1470 2392 -1464
rect 2411 -1469 2416 -1464
rect 2334 -1486 2408 -1470
rect 2426 -1478 2456 -1422
rect 2491 -1432 2699 -1422
rect 2734 -1426 2779 -1422
rect 2782 -1423 2783 -1422
rect 2798 -1423 2811 -1422
rect 2517 -1462 2706 -1432
rect 2532 -1465 2706 -1462
rect 2525 -1468 2706 -1465
rect 2334 -1488 2347 -1486
rect 2362 -1488 2396 -1486
rect 2334 -1504 2408 -1488
rect 2435 -1492 2448 -1478
rect 2463 -1492 2479 -1476
rect 2525 -1481 2536 -1468
rect 2318 -1526 2319 -1510
rect 2334 -1526 2347 -1504
rect 2362 -1526 2392 -1504
rect 2435 -1508 2497 -1492
rect 2525 -1499 2536 -1483
rect 2541 -1488 2551 -1468
rect 2561 -1488 2575 -1468
rect 2578 -1481 2587 -1468
rect 2603 -1481 2612 -1468
rect 2541 -1499 2575 -1488
rect 2578 -1499 2587 -1483
rect 2603 -1499 2612 -1483
rect 2619 -1488 2629 -1468
rect 2639 -1488 2653 -1468
rect 2654 -1481 2665 -1468
rect 2619 -1499 2653 -1488
rect 2654 -1499 2665 -1483
rect 2711 -1492 2727 -1476
rect 2734 -1478 2764 -1426
rect 2798 -1430 2799 -1423
rect 2783 -1438 2799 -1430
rect 2770 -1470 2783 -1451
rect 2798 -1470 2828 -1454
rect 2770 -1486 2844 -1470
rect 2770 -1488 2783 -1486
rect 2798 -1488 2832 -1486
rect 2435 -1510 2448 -1508
rect 2463 -1510 2497 -1508
rect 2435 -1526 2497 -1510
rect 2541 -1515 2557 -1512
rect 2619 -1515 2649 -1504
rect 2697 -1508 2743 -1492
rect 2770 -1504 2844 -1488
rect 2697 -1510 2731 -1508
rect 2696 -1526 2743 -1510
rect 2770 -1526 2783 -1504
rect 2798 -1526 2828 -1504
rect 2855 -1526 2856 -1510
rect 2871 -1526 2884 -1366
rect 2914 -1470 2927 -1366
rect 2972 -1388 2973 -1378
rect 2988 -1388 3001 -1378
rect 2972 -1392 3001 -1388
rect 3006 -1392 3036 -1366
rect 3054 -1380 3070 -1378
rect 3142 -1380 3195 -1366
rect 3143 -1382 3205 -1380
rect 3250 -1382 3265 -1366
rect 3314 -1369 3344 -1366
rect 3314 -1372 3350 -1369
rect 3280 -1380 3296 -1378
rect 3054 -1392 3069 -1388
rect 2972 -1394 3069 -1392
rect 3097 -1394 3265 -1382
rect 3281 -1392 3296 -1388
rect 3314 -1391 3353 -1372
rect 3372 -1378 3379 -1377
rect 3378 -1385 3379 -1378
rect 3362 -1388 3363 -1385
rect 3378 -1388 3391 -1385
rect 3314 -1392 3344 -1391
rect 3353 -1392 3359 -1391
rect 3362 -1392 3391 -1388
rect 3281 -1393 3391 -1392
rect 3281 -1394 3397 -1393
rect 2956 -1402 3007 -1394
rect 2956 -1414 2981 -1402
rect 2988 -1414 3007 -1402
rect 3038 -1402 3088 -1394
rect 3038 -1410 3054 -1402
rect 3061 -1404 3088 -1402
rect 3097 -1404 3318 -1394
rect 3061 -1414 3318 -1404
rect 3347 -1402 3397 -1394
rect 3347 -1411 3363 -1402
rect 2956 -1422 3007 -1414
rect 3054 -1422 3318 -1414
rect 3344 -1414 3363 -1411
rect 3370 -1414 3397 -1402
rect 3344 -1422 3397 -1414
rect 2972 -1430 2973 -1422
rect 2988 -1430 3001 -1422
rect 2972 -1438 2988 -1430
rect 2969 -1445 2988 -1442
rect 2969 -1454 2991 -1445
rect 2942 -1464 2991 -1454
rect 2942 -1470 2972 -1464
rect 2991 -1469 2996 -1464
rect 2914 -1486 2988 -1470
rect 3006 -1478 3036 -1422
rect 3071 -1432 3279 -1422
rect 3314 -1426 3359 -1422
rect 3362 -1423 3363 -1422
rect 3378 -1423 3391 -1422
rect 3097 -1462 3286 -1432
rect 3112 -1465 3286 -1462
rect 3105 -1468 3286 -1465
rect 2914 -1488 2927 -1486
rect 2942 -1488 2976 -1486
rect 2914 -1504 2988 -1488
rect 3015 -1492 3028 -1478
rect 3043 -1492 3059 -1476
rect 3105 -1481 3116 -1468
rect 2898 -1526 2899 -1510
rect 2914 -1526 2927 -1504
rect 2942 -1526 2972 -1504
rect 3015 -1508 3077 -1492
rect 3105 -1499 3116 -1483
rect 3121 -1488 3131 -1468
rect 3141 -1488 3155 -1468
rect 3158 -1481 3167 -1468
rect 3183 -1481 3192 -1468
rect 3121 -1499 3155 -1488
rect 3158 -1499 3167 -1483
rect 3183 -1499 3192 -1483
rect 3199 -1488 3209 -1468
rect 3219 -1488 3233 -1468
rect 3234 -1481 3245 -1468
rect 3199 -1499 3233 -1488
rect 3234 -1499 3245 -1483
rect 3291 -1492 3307 -1476
rect 3314 -1478 3344 -1426
rect 3378 -1430 3379 -1423
rect 3363 -1438 3379 -1430
rect 3350 -1470 3363 -1451
rect 3378 -1470 3408 -1454
rect 3350 -1486 3424 -1470
rect 3350 -1488 3363 -1486
rect 3378 -1488 3412 -1486
rect 3015 -1510 3028 -1508
rect 3043 -1510 3077 -1508
rect 3015 -1526 3077 -1510
rect 3121 -1515 3137 -1512
rect 3199 -1515 3229 -1504
rect 3277 -1508 3323 -1492
rect 3350 -1504 3424 -1488
rect 3277 -1510 3311 -1508
rect 3276 -1526 3323 -1510
rect 3350 -1526 3363 -1504
rect 3378 -1526 3408 -1504
rect 3435 -1526 3436 -1510
rect 3451 -1526 3464 -1366
rect 3494 -1470 3507 -1366
rect 3552 -1388 3553 -1378
rect 3568 -1388 3581 -1378
rect 3552 -1392 3581 -1388
rect 3586 -1392 3616 -1366
rect 3634 -1380 3650 -1378
rect 3722 -1380 3775 -1366
rect 3723 -1382 3787 -1380
rect 3830 -1382 3845 -1366
rect 3894 -1369 3924 -1366
rect 3894 -1372 3930 -1369
rect 3860 -1380 3876 -1378
rect 3634 -1392 3649 -1388
rect 3552 -1394 3649 -1392
rect 3677 -1394 3845 -1382
rect 3861 -1392 3876 -1388
rect 3894 -1391 3933 -1372
rect 3952 -1378 3959 -1377
rect 3958 -1385 3959 -1378
rect 3942 -1388 3943 -1385
rect 3958 -1388 3971 -1385
rect 3894 -1392 3924 -1391
rect 3933 -1392 3939 -1391
rect 3942 -1392 3971 -1388
rect 3861 -1393 3971 -1392
rect 3861 -1394 3977 -1393
rect 3536 -1402 3587 -1394
rect 3536 -1414 3561 -1402
rect 3568 -1414 3587 -1402
rect 3618 -1402 3668 -1394
rect 3618 -1410 3634 -1402
rect 3641 -1404 3668 -1402
rect 3677 -1404 3898 -1394
rect 3641 -1414 3898 -1404
rect 3927 -1402 3977 -1394
rect 3927 -1411 3943 -1402
rect 3536 -1422 3587 -1414
rect 3634 -1422 3898 -1414
rect 3924 -1414 3943 -1411
rect 3950 -1414 3977 -1402
rect 3924 -1422 3977 -1414
rect 3552 -1430 3553 -1422
rect 3568 -1430 3581 -1422
rect 3552 -1438 3568 -1430
rect 3549 -1445 3568 -1442
rect 3549 -1454 3571 -1445
rect 3522 -1464 3571 -1454
rect 3522 -1470 3552 -1464
rect 3571 -1469 3576 -1464
rect 3494 -1486 3568 -1470
rect 3586 -1478 3616 -1422
rect 3651 -1432 3859 -1422
rect 3894 -1426 3939 -1422
rect 3942 -1423 3943 -1422
rect 3958 -1423 3971 -1422
rect 3677 -1462 3866 -1432
rect 3692 -1465 3866 -1462
rect 3685 -1468 3866 -1465
rect 3494 -1488 3507 -1486
rect 3522 -1488 3556 -1486
rect 3494 -1504 3568 -1488
rect 3595 -1492 3608 -1478
rect 3623 -1492 3639 -1476
rect 3685 -1481 3696 -1468
rect 3478 -1526 3479 -1510
rect 3494 -1526 3507 -1504
rect 3522 -1526 3552 -1504
rect 3595 -1508 3657 -1492
rect 3685 -1499 3696 -1483
rect 3701 -1488 3711 -1468
rect 3721 -1488 3735 -1468
rect 3738 -1481 3747 -1468
rect 3763 -1481 3772 -1468
rect 3701 -1499 3735 -1488
rect 3738 -1499 3747 -1483
rect 3763 -1499 3772 -1483
rect 3779 -1488 3789 -1468
rect 3799 -1488 3813 -1468
rect 3814 -1481 3825 -1468
rect 3779 -1499 3813 -1488
rect 3814 -1499 3825 -1483
rect 3871 -1492 3887 -1476
rect 3894 -1478 3924 -1426
rect 3958 -1430 3959 -1423
rect 3943 -1438 3959 -1430
rect 3930 -1470 3943 -1451
rect 3958 -1470 3988 -1454
rect 3930 -1486 4004 -1470
rect 3930 -1488 3943 -1486
rect 3958 -1488 3992 -1486
rect 3595 -1510 3608 -1508
rect 3623 -1510 3657 -1508
rect 3595 -1526 3657 -1510
rect 3701 -1515 3717 -1512
rect 3779 -1515 3809 -1504
rect 3857 -1508 3903 -1492
rect 3930 -1504 4004 -1488
rect 3857 -1510 3891 -1508
rect 3856 -1526 3903 -1510
rect 3930 -1526 3943 -1504
rect 3958 -1526 3988 -1504
rect 4015 -1526 4016 -1510
rect 4031 -1526 4044 -1366
rect 4074 -1470 4087 -1366
rect 4132 -1388 4133 -1378
rect 4148 -1388 4161 -1378
rect 4132 -1392 4161 -1388
rect 4166 -1392 4196 -1366
rect 4214 -1380 4230 -1378
rect 4302 -1380 4355 -1366
rect 4303 -1382 4367 -1380
rect 4410 -1382 4425 -1366
rect 4474 -1369 4504 -1366
rect 4611 -1367 6944 -1366
rect 4474 -1372 4510 -1369
rect 4440 -1380 4456 -1378
rect 4214 -1392 4229 -1388
rect 4132 -1394 4229 -1392
rect 4257 -1394 4425 -1382
rect 4441 -1392 4456 -1388
rect 4474 -1391 4513 -1372
rect 4532 -1378 4539 -1377
rect 4538 -1385 4539 -1378
rect 4522 -1388 4523 -1385
rect 4538 -1388 4551 -1385
rect 4474 -1392 4504 -1391
rect 4513 -1392 4519 -1391
rect 4522 -1392 4551 -1388
rect 4441 -1393 4551 -1392
rect 4441 -1394 4557 -1393
rect 4116 -1402 4167 -1394
rect 4116 -1414 4141 -1402
rect 4148 -1414 4167 -1402
rect 4198 -1402 4248 -1394
rect 4198 -1410 4214 -1402
rect 4221 -1404 4248 -1402
rect 4257 -1404 4478 -1394
rect 4221 -1414 4478 -1404
rect 4507 -1402 4557 -1394
rect 4507 -1411 4523 -1402
rect 4116 -1422 4167 -1414
rect 4214 -1422 4478 -1414
rect 4504 -1414 4523 -1411
rect 4530 -1414 4557 -1402
rect 4504 -1422 4557 -1414
rect 4132 -1430 4133 -1422
rect 4148 -1430 4161 -1422
rect 4132 -1438 4148 -1430
rect 4129 -1445 4148 -1442
rect 4129 -1454 4151 -1445
rect 4102 -1464 4151 -1454
rect 4102 -1470 4132 -1464
rect 4151 -1469 4156 -1464
rect 4074 -1486 4148 -1470
rect 4166 -1478 4196 -1422
rect 4231 -1432 4439 -1422
rect 4474 -1426 4519 -1422
rect 4522 -1423 4523 -1422
rect 4538 -1423 4551 -1422
rect 4257 -1462 4446 -1432
rect 4272 -1465 4446 -1462
rect 4265 -1468 4446 -1465
rect 4074 -1488 4087 -1486
rect 4102 -1488 4136 -1486
rect 4074 -1504 4148 -1488
rect 4175 -1492 4188 -1478
rect 4203 -1492 4219 -1476
rect 4265 -1481 4276 -1468
rect 4058 -1526 4059 -1510
rect 4074 -1526 4087 -1504
rect 4102 -1526 4132 -1504
rect 4175 -1508 4237 -1492
rect 4265 -1499 4276 -1483
rect 4281 -1488 4291 -1468
rect 4301 -1488 4315 -1468
rect 4318 -1481 4327 -1468
rect 4343 -1481 4352 -1468
rect 4281 -1499 4315 -1488
rect 4318 -1499 4327 -1483
rect 4343 -1499 4352 -1483
rect 4359 -1488 4369 -1468
rect 4379 -1488 4393 -1468
rect 4394 -1481 4405 -1468
rect 4359 -1499 4393 -1488
rect 4394 -1499 4405 -1483
rect 4451 -1492 4467 -1476
rect 4474 -1478 4504 -1426
rect 4538 -1430 4539 -1423
rect 4523 -1438 4539 -1430
rect 4510 -1470 4523 -1451
rect 4538 -1470 4568 -1454
rect 4510 -1486 4584 -1470
rect 4510 -1488 4523 -1486
rect 4538 -1488 4572 -1486
rect 4175 -1510 4188 -1508
rect 4203 -1510 4237 -1508
rect 4175 -1526 4237 -1510
rect 4281 -1515 4297 -1512
rect 4359 -1515 4389 -1504
rect 4437 -1508 4483 -1492
rect 4510 -1504 4584 -1488
rect 4437 -1510 4471 -1508
rect 4436 -1526 4483 -1510
rect 4510 -1526 4523 -1504
rect 4538 -1526 4568 -1504
rect 4595 -1526 4596 -1510
rect 4611 -1526 4624 -1367
rect 4654 -1471 4667 -1367
rect 4712 -1389 4713 -1379
rect 4733 -1381 4741 -1379
rect 4731 -1383 4741 -1381
rect 4728 -1389 4741 -1383
rect 4712 -1393 4741 -1389
rect 4746 -1393 4776 -1367
rect 4794 -1381 4810 -1379
rect 4882 -1381 4933 -1367
rect 4883 -1383 4947 -1381
rect 4990 -1383 5005 -1367
rect 5054 -1370 5084 -1367
rect 5054 -1373 5090 -1370
rect 5020 -1381 5036 -1379
rect 4794 -1393 4809 -1389
rect 4712 -1395 4809 -1393
rect 4837 -1395 5005 -1383
rect 5021 -1393 5036 -1389
rect 5054 -1392 5093 -1373
rect 5112 -1379 5119 -1378
rect 5118 -1386 5119 -1379
rect 5102 -1389 5103 -1386
rect 5118 -1389 5131 -1386
rect 5054 -1393 5084 -1392
rect 5093 -1393 5099 -1392
rect 5102 -1393 5131 -1389
rect 5021 -1394 5131 -1393
rect 5021 -1395 5137 -1394
rect 4696 -1403 4747 -1395
rect 4696 -1415 4721 -1403
rect 4728 -1415 4747 -1403
rect 4778 -1403 4828 -1395
rect 4778 -1411 4794 -1403
rect 4801 -1405 4828 -1403
rect 4837 -1405 5058 -1395
rect 4801 -1415 5058 -1405
rect 5087 -1403 5137 -1395
rect 5087 -1412 5103 -1403
rect 4696 -1423 4747 -1415
rect 4794 -1423 5058 -1415
rect 5084 -1415 5103 -1412
rect 5110 -1415 5137 -1403
rect 5084 -1423 5137 -1415
rect 4712 -1431 4713 -1423
rect 4728 -1431 4741 -1423
rect 4712 -1439 4728 -1431
rect 4709 -1446 4728 -1443
rect 4709 -1455 4731 -1446
rect 4682 -1465 4731 -1455
rect 4682 -1471 4712 -1465
rect 4731 -1470 4736 -1465
rect 4654 -1487 4728 -1471
rect 4746 -1479 4776 -1423
rect 4811 -1433 5019 -1423
rect 5054 -1427 5099 -1423
rect 5102 -1424 5103 -1423
rect 5118 -1424 5131 -1423
rect 4837 -1463 5026 -1433
rect 4852 -1466 5026 -1463
rect 4845 -1469 5026 -1466
rect 4654 -1489 4667 -1487
rect 4682 -1489 4716 -1487
rect 4654 -1505 4728 -1489
rect 4755 -1493 4768 -1479
rect 4783 -1493 4799 -1477
rect 4845 -1482 4856 -1469
rect 0 -1534 33 -1526
rect 0 -1560 7 -1534
rect 14 -1560 33 -1534
rect 97 -1538 159 -1526
rect 171 -1538 246 -1526
rect 304 -1538 379 -1526
rect 391 -1538 422 -1526
rect 428 -1538 463 -1526
rect 97 -1540 259 -1538
rect 0 -1568 33 -1560
rect 115 -1564 128 -1540
rect 143 -1542 158 -1540
rect 14 -1578 27 -1568
rect 42 -1578 72 -1564
rect 115 -1578 158 -1564
rect 182 -1567 189 -1560
rect 192 -1564 259 -1540
rect 291 -1540 463 -1538
rect 261 -1562 289 -1558
rect 291 -1562 371 -1540
rect 392 -1542 407 -1540
rect 261 -1564 371 -1562
rect 192 -1568 371 -1564
rect 165 -1578 195 -1568
rect 197 -1578 350 -1568
rect 358 -1578 388 -1568
rect 392 -1578 422 -1564
rect 450 -1578 463 -1540
rect 535 -1534 570 -1526
rect 535 -1560 536 -1534
rect 543 -1560 570 -1534
rect 478 -1578 508 -1564
rect 535 -1568 570 -1560
rect 572 -1534 613 -1526
rect 572 -1560 587 -1534
rect 594 -1560 613 -1534
rect 677 -1538 739 -1526
rect 751 -1538 826 -1526
rect 884 -1538 959 -1526
rect 971 -1538 1002 -1526
rect 1008 -1538 1043 -1526
rect 677 -1540 839 -1538
rect 572 -1568 613 -1560
rect 695 -1564 708 -1540
rect 723 -1542 738 -1540
rect 535 -1578 536 -1568
rect 551 -1578 564 -1568
rect 578 -1578 579 -1568
rect 594 -1578 607 -1568
rect 622 -1578 652 -1564
rect 695 -1578 738 -1564
rect 762 -1567 769 -1560
rect 772 -1564 839 -1540
rect 871 -1540 1043 -1538
rect 841 -1562 869 -1558
rect 871 -1562 951 -1540
rect 972 -1542 987 -1540
rect 841 -1564 951 -1562
rect 772 -1568 951 -1564
rect 745 -1578 775 -1568
rect 777 -1578 930 -1568
rect 938 -1578 968 -1568
rect 972 -1578 1002 -1564
rect 1030 -1578 1043 -1540
rect 1115 -1534 1150 -1526
rect 1115 -1560 1116 -1534
rect 1123 -1560 1150 -1534
rect 1058 -1578 1088 -1564
rect 1115 -1568 1150 -1560
rect 1152 -1534 1193 -1526
rect 1152 -1560 1167 -1534
rect 1174 -1560 1193 -1534
rect 1257 -1538 1319 -1526
rect 1331 -1538 1406 -1526
rect 1464 -1538 1539 -1526
rect 1551 -1538 1582 -1526
rect 1588 -1538 1623 -1526
rect 1257 -1540 1419 -1538
rect 1152 -1568 1193 -1560
rect 1275 -1564 1288 -1540
rect 1303 -1542 1318 -1540
rect 1115 -1578 1116 -1568
rect 1131 -1578 1144 -1568
rect 1158 -1578 1159 -1568
rect 1174 -1578 1187 -1568
rect 1202 -1578 1232 -1564
rect 1275 -1578 1318 -1564
rect 1342 -1567 1349 -1560
rect 1352 -1564 1419 -1540
rect 1451 -1540 1623 -1538
rect 1421 -1562 1449 -1558
rect 1451 -1562 1531 -1540
rect 1552 -1542 1567 -1540
rect 1421 -1564 1531 -1562
rect 1352 -1568 1531 -1564
rect 1325 -1578 1355 -1568
rect 1357 -1578 1510 -1568
rect 1518 -1578 1548 -1568
rect 1552 -1578 1582 -1564
rect 1610 -1578 1623 -1540
rect 1695 -1534 1730 -1526
rect 1695 -1560 1696 -1534
rect 1703 -1560 1730 -1534
rect 1638 -1578 1668 -1564
rect 1695 -1568 1730 -1560
rect 1732 -1534 1773 -1526
rect 1732 -1560 1747 -1534
rect 1754 -1560 1773 -1534
rect 1837 -1538 1899 -1526
rect 1911 -1538 1986 -1526
rect 2044 -1538 2119 -1526
rect 2131 -1538 2162 -1526
rect 2168 -1538 2203 -1526
rect 1837 -1540 1999 -1538
rect 1732 -1568 1773 -1560
rect 1855 -1564 1868 -1540
rect 1883 -1542 1898 -1540
rect 1695 -1578 1696 -1568
rect 1711 -1578 1724 -1568
rect 1738 -1578 1739 -1568
rect 1754 -1578 1767 -1568
rect 1782 -1578 1812 -1564
rect 1855 -1578 1898 -1564
rect 1922 -1567 1929 -1560
rect 1932 -1564 1999 -1540
rect 2031 -1540 2203 -1538
rect 2001 -1562 2029 -1558
rect 2031 -1562 2111 -1540
rect 2132 -1542 2147 -1540
rect 2001 -1564 2111 -1562
rect 1932 -1568 2111 -1564
rect 1905 -1578 1935 -1568
rect 1937 -1578 2090 -1568
rect 2098 -1578 2128 -1568
rect 2132 -1578 2162 -1564
rect 2190 -1578 2203 -1540
rect 2275 -1534 2310 -1526
rect 2275 -1560 2276 -1534
rect 2283 -1560 2310 -1534
rect 2218 -1578 2248 -1564
rect 2275 -1568 2310 -1560
rect 2312 -1534 2353 -1526
rect 2312 -1560 2327 -1534
rect 2334 -1560 2353 -1534
rect 2417 -1538 2479 -1526
rect 2491 -1538 2566 -1526
rect 2624 -1538 2699 -1526
rect 2711 -1538 2742 -1526
rect 2748 -1538 2783 -1526
rect 2417 -1540 2579 -1538
rect 2312 -1568 2353 -1560
rect 2435 -1564 2448 -1540
rect 2463 -1542 2478 -1540
rect 2275 -1578 2276 -1568
rect 2291 -1578 2304 -1568
rect 2318 -1578 2319 -1568
rect 2334 -1578 2347 -1568
rect 2362 -1578 2392 -1564
rect 2435 -1578 2478 -1564
rect 2502 -1567 2509 -1560
rect 2512 -1564 2579 -1540
rect 2611 -1540 2783 -1538
rect 2581 -1562 2609 -1558
rect 2611 -1562 2691 -1540
rect 2712 -1542 2727 -1540
rect 2581 -1564 2691 -1562
rect 2512 -1568 2691 -1564
rect 2485 -1578 2515 -1568
rect 2517 -1578 2670 -1568
rect 2678 -1578 2708 -1568
rect 2712 -1578 2742 -1564
rect 2770 -1578 2783 -1540
rect 2855 -1534 2890 -1526
rect 2855 -1560 2856 -1534
rect 2863 -1560 2890 -1534
rect 2798 -1578 2828 -1564
rect 2855 -1568 2890 -1560
rect 2892 -1534 2933 -1526
rect 2892 -1560 2907 -1534
rect 2914 -1560 2933 -1534
rect 2997 -1538 3059 -1526
rect 3071 -1538 3146 -1526
rect 3204 -1538 3279 -1526
rect 3291 -1538 3322 -1526
rect 3328 -1538 3363 -1526
rect 2997 -1540 3159 -1538
rect 2892 -1568 2933 -1560
rect 3015 -1564 3028 -1540
rect 3043 -1542 3058 -1540
rect 2855 -1578 2856 -1568
rect 2871 -1578 2884 -1568
rect 2898 -1578 2899 -1568
rect 2914 -1578 2927 -1568
rect 2942 -1578 2972 -1564
rect 3015 -1578 3058 -1564
rect 3082 -1567 3089 -1560
rect 3092 -1564 3159 -1540
rect 3191 -1540 3363 -1538
rect 3161 -1562 3189 -1558
rect 3191 -1562 3271 -1540
rect 3292 -1542 3307 -1540
rect 3161 -1564 3271 -1562
rect 3092 -1568 3271 -1564
rect 3065 -1578 3095 -1568
rect 3097 -1578 3250 -1568
rect 3258 -1578 3288 -1568
rect 3292 -1578 3322 -1564
rect 3350 -1578 3363 -1540
rect 3435 -1534 3470 -1526
rect 3435 -1560 3436 -1534
rect 3443 -1560 3470 -1534
rect 3378 -1578 3408 -1564
rect 3435 -1568 3470 -1560
rect 3472 -1534 3513 -1526
rect 3472 -1560 3487 -1534
rect 3494 -1560 3513 -1534
rect 3577 -1538 3639 -1526
rect 3651 -1538 3726 -1526
rect 3784 -1538 3859 -1526
rect 3871 -1538 3902 -1526
rect 3908 -1538 3943 -1526
rect 3577 -1540 3739 -1538
rect 3472 -1568 3513 -1560
rect 3595 -1564 3608 -1540
rect 3623 -1542 3638 -1540
rect 3435 -1578 3436 -1568
rect 3451 -1578 3464 -1568
rect 3478 -1578 3479 -1568
rect 3494 -1578 3507 -1568
rect 3522 -1578 3552 -1564
rect 3595 -1578 3638 -1564
rect 3662 -1567 3669 -1560
rect 3672 -1564 3739 -1540
rect 3771 -1540 3943 -1538
rect 3741 -1562 3769 -1558
rect 3771 -1562 3851 -1540
rect 3872 -1542 3887 -1540
rect 3741 -1564 3851 -1562
rect 3672 -1568 3851 -1564
rect 3645 -1578 3675 -1568
rect 3677 -1578 3830 -1568
rect 3838 -1578 3868 -1568
rect 3872 -1578 3902 -1564
rect 3930 -1578 3943 -1540
rect 4015 -1534 4050 -1526
rect 4015 -1560 4016 -1534
rect 4023 -1560 4050 -1534
rect 3958 -1578 3988 -1564
rect 4015 -1568 4050 -1560
rect 4052 -1534 4093 -1526
rect 4052 -1560 4067 -1534
rect 4074 -1560 4093 -1534
rect 4157 -1538 4219 -1526
rect 4231 -1538 4306 -1526
rect 4364 -1538 4439 -1526
rect 4451 -1538 4482 -1526
rect 4488 -1538 4523 -1526
rect 4157 -1540 4319 -1538
rect 4052 -1568 4093 -1560
rect 4175 -1564 4188 -1540
rect 4203 -1542 4218 -1540
rect 4015 -1578 4016 -1568
rect 4031 -1578 4044 -1568
rect 4058 -1578 4059 -1568
rect 4074 -1578 4087 -1568
rect 4102 -1578 4132 -1564
rect 4175 -1578 4218 -1564
rect 4242 -1567 4249 -1560
rect 4252 -1564 4319 -1540
rect 4351 -1540 4523 -1538
rect 4321 -1562 4349 -1558
rect 4351 -1562 4431 -1540
rect 4452 -1542 4467 -1540
rect 4321 -1564 4431 -1562
rect 4252 -1568 4431 -1564
rect 4225 -1578 4255 -1568
rect 4257 -1578 4410 -1568
rect 4418 -1578 4448 -1568
rect 4452 -1578 4482 -1564
rect 4510 -1578 4523 -1540
rect 4595 -1534 4630 -1526
rect 4638 -1527 4639 -1511
rect 4654 -1527 4667 -1505
rect 4682 -1527 4712 -1505
rect 4755 -1509 4817 -1493
rect 4845 -1500 4856 -1484
rect 4861 -1489 4871 -1469
rect 4881 -1489 4895 -1469
rect 4898 -1482 4907 -1469
rect 4923 -1482 4932 -1469
rect 4861 -1500 4895 -1489
rect 4898 -1500 4907 -1484
rect 4923 -1500 4932 -1484
rect 4939 -1489 4949 -1469
rect 4959 -1489 4973 -1469
rect 4974 -1482 4985 -1469
rect 4939 -1500 4973 -1489
rect 4974 -1500 4985 -1484
rect 5031 -1493 5047 -1477
rect 5054 -1479 5084 -1427
rect 5118 -1431 5119 -1424
rect 5103 -1439 5119 -1431
rect 5090 -1471 5103 -1452
rect 5118 -1471 5148 -1455
rect 5090 -1487 5164 -1471
rect 5090 -1489 5103 -1487
rect 5118 -1489 5152 -1487
rect 4755 -1511 4768 -1509
rect 4783 -1511 4817 -1509
rect 4755 -1527 4817 -1511
rect 4861 -1516 4877 -1513
rect 4939 -1516 4969 -1505
rect 5017 -1509 5063 -1493
rect 5090 -1505 5164 -1489
rect 5017 -1511 5051 -1509
rect 5016 -1527 5063 -1511
rect 5090 -1527 5103 -1505
rect 5118 -1527 5148 -1505
rect 5175 -1527 5176 -1511
rect 5191 -1527 5204 -1367
rect 5234 -1471 5247 -1367
rect 5292 -1389 5293 -1379
rect 5313 -1381 5321 -1379
rect 5311 -1383 5321 -1381
rect 5308 -1389 5321 -1383
rect 5292 -1393 5321 -1389
rect 5326 -1393 5356 -1367
rect 5374 -1381 5390 -1379
rect 5462 -1381 5513 -1367
rect 5463 -1383 5527 -1381
rect 5570 -1383 5585 -1367
rect 5634 -1370 5664 -1367
rect 5634 -1373 5670 -1370
rect 5600 -1381 5616 -1379
rect 5374 -1393 5389 -1389
rect 5292 -1395 5389 -1393
rect 5417 -1395 5585 -1383
rect 5601 -1393 5616 -1389
rect 5634 -1392 5673 -1373
rect 5692 -1379 5699 -1378
rect 5698 -1386 5699 -1379
rect 5682 -1389 5683 -1386
rect 5698 -1389 5711 -1386
rect 5634 -1393 5664 -1392
rect 5673 -1393 5679 -1392
rect 5682 -1393 5711 -1389
rect 5601 -1394 5711 -1393
rect 5601 -1395 5717 -1394
rect 5276 -1403 5327 -1395
rect 5276 -1415 5301 -1403
rect 5308 -1415 5327 -1403
rect 5358 -1403 5408 -1395
rect 5358 -1411 5374 -1403
rect 5381 -1405 5408 -1403
rect 5417 -1405 5638 -1395
rect 5381 -1415 5638 -1405
rect 5667 -1403 5717 -1395
rect 5667 -1412 5683 -1403
rect 5276 -1423 5327 -1415
rect 5374 -1423 5638 -1415
rect 5664 -1415 5683 -1412
rect 5690 -1415 5717 -1403
rect 5664 -1423 5717 -1415
rect 5292 -1431 5293 -1423
rect 5308 -1431 5321 -1423
rect 5292 -1439 5308 -1431
rect 5289 -1446 5308 -1443
rect 5289 -1455 5311 -1446
rect 5262 -1465 5311 -1455
rect 5262 -1471 5292 -1465
rect 5311 -1470 5316 -1465
rect 5234 -1487 5308 -1471
rect 5326 -1479 5356 -1423
rect 5391 -1433 5599 -1423
rect 5634 -1427 5679 -1423
rect 5682 -1424 5683 -1423
rect 5698 -1424 5711 -1423
rect 5417 -1463 5606 -1433
rect 5432 -1466 5606 -1463
rect 5425 -1469 5606 -1466
rect 5234 -1489 5247 -1487
rect 5262 -1489 5296 -1487
rect 5234 -1505 5308 -1489
rect 5335 -1493 5348 -1479
rect 5363 -1493 5379 -1477
rect 5425 -1482 5436 -1469
rect 5218 -1527 5219 -1511
rect 5234 -1527 5247 -1505
rect 5262 -1527 5292 -1505
rect 5335 -1509 5397 -1493
rect 5425 -1500 5436 -1484
rect 5441 -1489 5451 -1469
rect 5461 -1489 5475 -1469
rect 5478 -1482 5487 -1469
rect 5503 -1482 5512 -1469
rect 5441 -1500 5475 -1489
rect 5478 -1500 5487 -1484
rect 5503 -1500 5512 -1484
rect 5519 -1489 5529 -1469
rect 5539 -1489 5553 -1469
rect 5554 -1482 5565 -1469
rect 5519 -1500 5553 -1489
rect 5554 -1500 5565 -1484
rect 5611 -1493 5627 -1477
rect 5634 -1479 5664 -1427
rect 5698 -1431 5699 -1424
rect 5683 -1439 5699 -1431
rect 5670 -1471 5683 -1452
rect 5698 -1471 5728 -1455
rect 5670 -1487 5744 -1471
rect 5670 -1489 5683 -1487
rect 5698 -1489 5732 -1487
rect 5335 -1511 5348 -1509
rect 5363 -1511 5397 -1509
rect 5335 -1527 5397 -1511
rect 5441 -1516 5457 -1513
rect 5519 -1516 5549 -1505
rect 5597 -1509 5643 -1493
rect 5670 -1505 5744 -1489
rect 5597 -1511 5631 -1509
rect 5596 -1527 5643 -1511
rect 5670 -1527 5683 -1505
rect 5698 -1527 5728 -1505
rect 5755 -1527 5756 -1511
rect 5771 -1527 5784 -1367
rect 5814 -1471 5827 -1367
rect 5872 -1389 5873 -1379
rect 5893 -1381 5901 -1379
rect 5891 -1383 5901 -1381
rect 5888 -1389 5901 -1383
rect 5872 -1393 5901 -1389
rect 5906 -1393 5936 -1367
rect 5954 -1381 5970 -1379
rect 6042 -1381 6093 -1367
rect 6043 -1383 6107 -1381
rect 6150 -1383 6165 -1367
rect 6214 -1370 6244 -1367
rect 6214 -1373 6250 -1370
rect 6180 -1381 6196 -1379
rect 5954 -1393 5969 -1389
rect 5872 -1395 5969 -1393
rect 5997 -1395 6165 -1383
rect 6181 -1393 6196 -1389
rect 6214 -1392 6253 -1373
rect 6272 -1379 6279 -1378
rect 6278 -1386 6279 -1379
rect 6262 -1389 6263 -1386
rect 6278 -1389 6291 -1386
rect 6214 -1393 6244 -1392
rect 6253 -1393 6259 -1392
rect 6262 -1393 6291 -1389
rect 6181 -1394 6291 -1393
rect 6181 -1395 6297 -1394
rect 5856 -1403 5907 -1395
rect 5856 -1415 5881 -1403
rect 5888 -1415 5907 -1403
rect 5938 -1403 5988 -1395
rect 5938 -1411 5954 -1403
rect 5961 -1405 5988 -1403
rect 5997 -1405 6218 -1395
rect 5961 -1415 6218 -1405
rect 6247 -1403 6297 -1395
rect 6247 -1412 6263 -1403
rect 5856 -1423 5907 -1415
rect 5954 -1423 6218 -1415
rect 6244 -1415 6263 -1412
rect 6270 -1415 6297 -1403
rect 6244 -1423 6297 -1415
rect 5872 -1431 5873 -1423
rect 5888 -1431 5901 -1423
rect 5872 -1439 5888 -1431
rect 5869 -1446 5888 -1443
rect 5869 -1455 5891 -1446
rect 5842 -1465 5891 -1455
rect 5842 -1471 5872 -1465
rect 5891 -1470 5896 -1465
rect 5814 -1487 5888 -1471
rect 5906 -1479 5936 -1423
rect 5971 -1433 6179 -1423
rect 6214 -1427 6259 -1423
rect 6262 -1424 6263 -1423
rect 6278 -1424 6291 -1423
rect 5997 -1463 6186 -1433
rect 6012 -1466 6186 -1463
rect 6005 -1469 6186 -1466
rect 5814 -1489 5827 -1487
rect 5842 -1489 5876 -1487
rect 5814 -1505 5888 -1489
rect 5915 -1493 5928 -1479
rect 5943 -1493 5959 -1477
rect 6005 -1482 6016 -1469
rect 5798 -1527 5799 -1511
rect 5814 -1527 5827 -1505
rect 5842 -1527 5872 -1505
rect 5915 -1509 5977 -1493
rect 6005 -1500 6016 -1484
rect 6021 -1489 6031 -1469
rect 6041 -1489 6055 -1469
rect 6058 -1482 6067 -1469
rect 6083 -1482 6092 -1469
rect 6021 -1500 6055 -1489
rect 6058 -1500 6067 -1484
rect 6083 -1500 6092 -1484
rect 6099 -1489 6109 -1469
rect 6119 -1489 6133 -1469
rect 6134 -1482 6145 -1469
rect 6099 -1500 6133 -1489
rect 6134 -1500 6145 -1484
rect 6191 -1493 6207 -1477
rect 6214 -1479 6244 -1427
rect 6278 -1431 6279 -1424
rect 6263 -1439 6279 -1431
rect 6250 -1471 6263 -1452
rect 6278 -1471 6308 -1455
rect 6250 -1487 6324 -1471
rect 6250 -1489 6263 -1487
rect 6278 -1489 6312 -1487
rect 5915 -1511 5928 -1509
rect 5943 -1511 5977 -1509
rect 5915 -1527 5977 -1511
rect 6021 -1516 6037 -1513
rect 6099 -1516 6129 -1505
rect 6177 -1509 6223 -1493
rect 6250 -1505 6324 -1489
rect 6177 -1511 6211 -1509
rect 6176 -1527 6223 -1511
rect 6250 -1527 6263 -1505
rect 6278 -1527 6308 -1505
rect 6335 -1527 6336 -1511
rect 6351 -1527 6364 -1367
rect 6394 -1471 6407 -1367
rect 6452 -1389 6453 -1379
rect 6473 -1381 6481 -1379
rect 6471 -1383 6481 -1381
rect 6468 -1389 6481 -1383
rect 6452 -1393 6481 -1389
rect 6486 -1393 6516 -1367
rect 6534 -1381 6550 -1379
rect 6622 -1381 6673 -1367
rect 6623 -1383 6687 -1381
rect 6730 -1383 6745 -1367
rect 6794 -1370 6824 -1367
rect 6794 -1373 6830 -1370
rect 6760 -1381 6776 -1379
rect 6534 -1393 6549 -1389
rect 6452 -1395 6549 -1393
rect 6577 -1395 6745 -1383
rect 6761 -1393 6776 -1389
rect 6794 -1392 6833 -1373
rect 6852 -1379 6859 -1378
rect 6858 -1386 6859 -1379
rect 6842 -1389 6843 -1386
rect 6858 -1389 6871 -1386
rect 6794 -1393 6824 -1392
rect 6833 -1393 6839 -1392
rect 6842 -1393 6871 -1389
rect 6761 -1394 6871 -1393
rect 6761 -1395 6877 -1394
rect 6436 -1403 6487 -1395
rect 6436 -1415 6461 -1403
rect 6468 -1415 6487 -1403
rect 6518 -1403 6568 -1395
rect 6518 -1411 6534 -1403
rect 6541 -1405 6568 -1403
rect 6577 -1405 6798 -1395
rect 6541 -1415 6798 -1405
rect 6827 -1403 6877 -1395
rect 6827 -1412 6843 -1403
rect 6436 -1423 6487 -1415
rect 6534 -1423 6798 -1415
rect 6824 -1415 6843 -1412
rect 6850 -1415 6877 -1403
rect 6824 -1423 6877 -1415
rect 6452 -1431 6453 -1423
rect 6468 -1431 6481 -1423
rect 6452 -1439 6468 -1431
rect 6449 -1446 6468 -1443
rect 6449 -1455 6471 -1446
rect 6422 -1465 6471 -1455
rect 6422 -1471 6452 -1465
rect 6471 -1470 6476 -1465
rect 6394 -1487 6468 -1471
rect 6486 -1479 6516 -1423
rect 6551 -1433 6759 -1423
rect 6794 -1427 6839 -1423
rect 6842 -1424 6843 -1423
rect 6858 -1424 6871 -1423
rect 6577 -1463 6766 -1433
rect 6592 -1466 6766 -1463
rect 6585 -1469 6766 -1466
rect 6394 -1489 6407 -1487
rect 6422 -1489 6456 -1487
rect 6394 -1505 6468 -1489
rect 6495 -1493 6508 -1479
rect 6523 -1493 6539 -1477
rect 6585 -1482 6596 -1469
rect 6378 -1527 6379 -1511
rect 6394 -1527 6407 -1505
rect 6422 -1527 6452 -1505
rect 6495 -1509 6557 -1493
rect 6585 -1500 6596 -1484
rect 6601 -1489 6611 -1469
rect 6621 -1489 6635 -1469
rect 6638 -1482 6647 -1469
rect 6663 -1482 6672 -1469
rect 6601 -1500 6635 -1489
rect 6638 -1500 6647 -1484
rect 6663 -1500 6672 -1484
rect 6679 -1489 6689 -1469
rect 6699 -1489 6713 -1469
rect 6714 -1482 6725 -1469
rect 6679 -1500 6713 -1489
rect 6714 -1500 6725 -1484
rect 6771 -1493 6787 -1477
rect 6794 -1479 6824 -1427
rect 6858 -1431 6859 -1424
rect 6843 -1439 6859 -1431
rect 6830 -1471 6843 -1452
rect 6858 -1471 6888 -1455
rect 6830 -1487 6904 -1471
rect 6830 -1489 6843 -1487
rect 6858 -1489 6892 -1487
rect 6495 -1511 6508 -1509
rect 6523 -1511 6557 -1509
rect 6495 -1527 6557 -1511
rect 6601 -1516 6617 -1513
rect 6679 -1516 6709 -1505
rect 6757 -1509 6803 -1493
rect 6830 -1505 6904 -1489
rect 6757 -1511 6791 -1509
rect 6756 -1527 6803 -1511
rect 6830 -1527 6843 -1505
rect 6858 -1527 6888 -1505
rect 6915 -1527 6916 -1511
rect 6931 -1527 6944 -1367
rect 4595 -1560 4596 -1534
rect 4603 -1560 4630 -1534
rect 4538 -1578 4568 -1564
rect 4595 -1568 4630 -1560
rect 4632 -1535 4673 -1527
rect 4632 -1561 4647 -1535
rect 4654 -1561 4673 -1535
rect 4737 -1539 4799 -1527
rect 4811 -1539 4886 -1527
rect 4944 -1539 5019 -1527
rect 5031 -1539 5062 -1527
rect 5068 -1539 5103 -1527
rect 4737 -1541 4899 -1539
rect 4755 -1559 4768 -1541
rect 4783 -1543 4798 -1541
rect 4595 -1578 4596 -1568
rect 4611 -1578 4624 -1568
rect 4632 -1569 4673 -1561
rect 4756 -1565 4768 -1559
rect 4832 -1559 4899 -1541
rect 4931 -1541 5103 -1539
rect 4931 -1559 5011 -1541
rect 5032 -1543 5047 -1541
rect 0 -1579 4624 -1578
rect 4638 -1579 4639 -1569
rect 4654 -1579 4667 -1569
rect 4682 -1579 4712 -1565
rect 4756 -1579 4798 -1565
rect 4822 -1568 4829 -1561
rect 4832 -1569 5011 -1559
rect 4805 -1579 4835 -1569
rect 4837 -1579 4990 -1569
rect 4998 -1579 5028 -1569
rect 5032 -1579 5062 -1565
rect 5090 -1579 5103 -1541
rect 5175 -1535 5210 -1527
rect 5175 -1561 5176 -1535
rect 5183 -1561 5210 -1535
rect 5118 -1579 5148 -1565
rect 5175 -1569 5210 -1561
rect 5212 -1535 5253 -1527
rect 5212 -1561 5227 -1535
rect 5234 -1561 5253 -1535
rect 5317 -1539 5379 -1527
rect 5391 -1539 5466 -1527
rect 5524 -1539 5599 -1527
rect 5611 -1539 5642 -1527
rect 5648 -1539 5683 -1527
rect 5317 -1541 5479 -1539
rect 5335 -1559 5348 -1541
rect 5363 -1543 5378 -1541
rect 5212 -1569 5253 -1561
rect 5336 -1565 5348 -1559
rect 5412 -1559 5479 -1541
rect 5511 -1541 5683 -1539
rect 5511 -1559 5591 -1541
rect 5612 -1543 5627 -1541
rect 5175 -1579 5176 -1569
rect 5191 -1579 5204 -1569
rect 5218 -1579 5219 -1569
rect 5234 -1579 5247 -1569
rect 5262 -1579 5292 -1565
rect 5336 -1579 5378 -1565
rect 5402 -1568 5409 -1561
rect 5412 -1569 5591 -1559
rect 5385 -1579 5415 -1569
rect 5417 -1579 5570 -1569
rect 5578 -1579 5608 -1569
rect 5612 -1579 5642 -1565
rect 5670 -1579 5683 -1541
rect 5755 -1535 5790 -1527
rect 5755 -1561 5756 -1535
rect 5763 -1561 5790 -1535
rect 5698 -1579 5728 -1565
rect 5755 -1569 5790 -1561
rect 5792 -1535 5833 -1527
rect 5792 -1561 5807 -1535
rect 5814 -1561 5833 -1535
rect 5897 -1539 5959 -1527
rect 5971 -1539 6046 -1527
rect 6104 -1539 6179 -1527
rect 6191 -1539 6222 -1527
rect 6228 -1539 6263 -1527
rect 5897 -1541 6059 -1539
rect 5915 -1559 5928 -1541
rect 5943 -1543 5958 -1541
rect 5792 -1569 5833 -1561
rect 5916 -1565 5928 -1559
rect 5992 -1559 6059 -1541
rect 6091 -1541 6263 -1539
rect 6091 -1559 6171 -1541
rect 6192 -1543 6207 -1541
rect 5755 -1579 5756 -1569
rect 5771 -1579 5784 -1569
rect 5798 -1579 5799 -1569
rect 5814 -1579 5827 -1569
rect 5842 -1579 5872 -1565
rect 5916 -1579 5958 -1565
rect 5982 -1568 5989 -1561
rect 5992 -1569 6171 -1559
rect 5965 -1579 5995 -1569
rect 5997 -1579 6150 -1569
rect 6158 -1579 6188 -1569
rect 6192 -1579 6222 -1565
rect 6250 -1579 6263 -1541
rect 6335 -1535 6370 -1527
rect 6335 -1561 6336 -1535
rect 6343 -1561 6370 -1535
rect 6278 -1579 6308 -1565
rect 6335 -1569 6370 -1561
rect 6372 -1535 6413 -1527
rect 6372 -1561 6387 -1535
rect 6394 -1561 6413 -1535
rect 6477 -1539 6539 -1527
rect 6551 -1539 6626 -1527
rect 6684 -1539 6759 -1527
rect 6771 -1539 6802 -1527
rect 6808 -1539 6843 -1527
rect 6477 -1541 6639 -1539
rect 6495 -1559 6508 -1541
rect 6523 -1543 6538 -1541
rect 6372 -1569 6413 -1561
rect 6496 -1565 6508 -1559
rect 6572 -1559 6639 -1541
rect 6671 -1541 6843 -1539
rect 6671 -1559 6751 -1541
rect 6772 -1543 6787 -1541
rect 6335 -1579 6336 -1569
rect 6351 -1579 6364 -1569
rect 6378 -1579 6379 -1569
rect 6394 -1579 6407 -1569
rect 6422 -1579 6452 -1565
rect 6496 -1579 6538 -1565
rect 6562 -1568 6569 -1561
rect 6572 -1569 6751 -1559
rect 6545 -1579 6575 -1569
rect 6577 -1579 6730 -1569
rect 6738 -1579 6768 -1569
rect 6772 -1579 6802 -1565
rect 6830 -1579 6843 -1541
rect 6915 -1535 6950 -1527
rect 6915 -1561 6916 -1535
rect 6923 -1561 6950 -1535
rect 6858 -1579 6888 -1565
rect 6915 -1569 6950 -1561
rect 6915 -1579 6916 -1569
rect 6931 -1579 6944 -1569
rect 0 -1592 6944 -1579
rect 14 -1622 27 -1592
rect 42 -1610 72 -1592
rect 115 -1606 129 -1592
rect 165 -1606 385 -1592
rect 116 -1608 129 -1606
rect 82 -1620 97 -1608
rect 79 -1622 101 -1620
rect 106 -1622 136 -1608
rect 197 -1610 350 -1606
rect 179 -1622 371 -1610
rect 414 -1622 444 -1608
rect 450 -1622 463 -1592
rect 478 -1610 508 -1592
rect 551 -1622 564 -1592
rect 594 -1622 607 -1592
rect 622 -1610 652 -1592
rect 695 -1606 709 -1592
rect 745 -1606 965 -1592
rect 696 -1608 709 -1606
rect 662 -1620 677 -1608
rect 659 -1622 681 -1620
rect 686 -1622 716 -1608
rect 777 -1610 930 -1606
rect 759 -1622 951 -1610
rect 994 -1622 1024 -1608
rect 1030 -1622 1043 -1592
rect 1058 -1610 1088 -1592
rect 1131 -1622 1144 -1592
rect 1174 -1622 1187 -1592
rect 1202 -1610 1232 -1592
rect 1275 -1606 1289 -1592
rect 1325 -1606 1545 -1592
rect 1276 -1608 1289 -1606
rect 1242 -1620 1257 -1608
rect 1239 -1622 1261 -1620
rect 1266 -1622 1296 -1608
rect 1357 -1610 1510 -1606
rect 1339 -1622 1531 -1610
rect 1574 -1622 1604 -1608
rect 1610 -1622 1623 -1592
rect 1638 -1610 1668 -1592
rect 1711 -1622 1724 -1592
rect 1754 -1622 1767 -1592
rect 1782 -1610 1812 -1592
rect 1855 -1606 1869 -1592
rect 1905 -1606 2125 -1592
rect 1856 -1608 1869 -1606
rect 1822 -1620 1837 -1608
rect 1819 -1622 1841 -1620
rect 1846 -1622 1876 -1608
rect 1937 -1610 2090 -1606
rect 1919 -1622 2111 -1610
rect 2154 -1622 2184 -1608
rect 2190 -1622 2203 -1592
rect 2218 -1610 2248 -1592
rect 2291 -1622 2304 -1592
rect 2334 -1622 2347 -1592
rect 2362 -1610 2392 -1592
rect 2435 -1606 2449 -1592
rect 2485 -1606 2705 -1592
rect 2436 -1608 2449 -1606
rect 2402 -1620 2417 -1608
rect 2399 -1622 2421 -1620
rect 2426 -1622 2456 -1608
rect 2517 -1610 2670 -1606
rect 2499 -1622 2691 -1610
rect 2734 -1622 2764 -1608
rect 2770 -1622 2783 -1592
rect 2798 -1610 2828 -1592
rect 2871 -1622 2884 -1592
rect 2914 -1622 2927 -1592
rect 2942 -1610 2972 -1592
rect 3015 -1606 3029 -1592
rect 3065 -1606 3285 -1592
rect 3016 -1608 3029 -1606
rect 2982 -1620 2997 -1608
rect 2979 -1622 3001 -1620
rect 3006 -1622 3036 -1608
rect 3097 -1610 3250 -1606
rect 3079 -1622 3271 -1610
rect 3314 -1622 3344 -1608
rect 3350 -1622 3363 -1592
rect 3378 -1610 3408 -1592
rect 3451 -1622 3464 -1592
rect 3494 -1622 3507 -1592
rect 3522 -1610 3552 -1592
rect 3595 -1606 3609 -1592
rect 3645 -1606 3865 -1592
rect 3596 -1608 3609 -1606
rect 3562 -1620 3577 -1608
rect 3559 -1622 3581 -1620
rect 3586 -1622 3616 -1608
rect 3677 -1610 3830 -1606
rect 3659 -1622 3851 -1610
rect 3894 -1622 3924 -1608
rect 3930 -1622 3943 -1592
rect 3958 -1610 3988 -1592
rect 4031 -1622 4044 -1592
rect 4074 -1622 4087 -1592
rect 4102 -1610 4132 -1592
rect 4175 -1606 4189 -1592
rect 4225 -1606 4445 -1592
rect 4176 -1608 4189 -1606
rect 4142 -1620 4157 -1608
rect 4139 -1622 4161 -1620
rect 4166 -1622 4196 -1608
rect 4257 -1610 4410 -1606
rect 4239 -1622 4431 -1610
rect 4474 -1622 4504 -1608
rect 4510 -1622 4523 -1592
rect 4538 -1610 4568 -1592
rect 4611 -1593 6944 -1592
rect 4611 -1622 4624 -1593
rect 0 -1623 4624 -1622
rect 4654 -1623 4667 -1593
rect 4682 -1611 4712 -1593
rect 4756 -1609 4769 -1593
rect 4805 -1607 5025 -1593
rect 4722 -1621 4737 -1609
rect 4719 -1623 4741 -1621
rect 4746 -1623 4776 -1609
rect 4837 -1611 4990 -1607
rect 4819 -1623 5011 -1611
rect 5054 -1623 5084 -1609
rect 5090 -1623 5103 -1593
rect 5118 -1611 5148 -1593
rect 5191 -1623 5204 -1593
rect 5234 -1623 5247 -1593
rect 5262 -1611 5292 -1593
rect 5336 -1609 5349 -1593
rect 5385 -1607 5605 -1593
rect 5302 -1621 5317 -1609
rect 5299 -1623 5321 -1621
rect 5326 -1623 5356 -1609
rect 5417 -1611 5570 -1607
rect 5399 -1623 5591 -1611
rect 5634 -1623 5664 -1609
rect 5670 -1623 5683 -1593
rect 5698 -1611 5728 -1593
rect 5771 -1623 5784 -1593
rect 5814 -1623 5827 -1593
rect 5842 -1611 5872 -1593
rect 5916 -1609 5929 -1593
rect 5965 -1607 6185 -1593
rect 5882 -1621 5897 -1609
rect 5879 -1623 5901 -1621
rect 5906 -1623 5936 -1609
rect 5997 -1611 6150 -1607
rect 5979 -1623 6171 -1611
rect 6214 -1623 6244 -1609
rect 6250 -1623 6263 -1593
rect 6278 -1611 6308 -1593
rect 6351 -1623 6364 -1593
rect 6394 -1623 6407 -1593
rect 6422 -1611 6452 -1593
rect 6496 -1609 6509 -1593
rect 6545 -1607 6765 -1593
rect 6462 -1621 6477 -1609
rect 6459 -1623 6481 -1621
rect 6486 -1623 6516 -1609
rect 6577 -1611 6730 -1607
rect 6559 -1623 6751 -1611
rect 6794 -1623 6824 -1609
rect 6830 -1623 6843 -1593
rect 6858 -1611 6888 -1593
rect 6931 -1623 6944 -1593
rect 0 -1636 6944 -1623
rect 14 -1740 27 -1636
rect 72 -1658 73 -1648
rect 88 -1658 101 -1648
rect 72 -1662 101 -1658
rect 106 -1662 136 -1636
rect 154 -1650 170 -1648
rect 242 -1650 295 -1636
rect 243 -1652 307 -1650
rect 350 -1652 365 -1636
rect 414 -1639 444 -1636
rect 414 -1642 450 -1639
rect 380 -1650 396 -1648
rect 154 -1662 169 -1658
rect 72 -1664 169 -1662
rect 197 -1664 365 -1652
rect 381 -1662 396 -1658
rect 414 -1661 453 -1642
rect 472 -1648 479 -1647
rect 478 -1655 479 -1648
rect 462 -1658 463 -1655
rect 478 -1658 491 -1655
rect 414 -1662 444 -1661
rect 453 -1662 459 -1661
rect 462 -1662 491 -1658
rect 381 -1663 491 -1662
rect 381 -1664 497 -1663
rect 56 -1672 107 -1664
rect 56 -1684 81 -1672
rect 88 -1684 107 -1672
rect 138 -1672 188 -1664
rect 138 -1680 154 -1672
rect 161 -1674 188 -1672
rect 197 -1674 418 -1664
rect 161 -1684 418 -1674
rect 447 -1672 497 -1664
rect 447 -1681 463 -1672
rect 56 -1692 107 -1684
rect 154 -1692 418 -1684
rect 444 -1684 463 -1681
rect 470 -1684 497 -1672
rect 444 -1692 497 -1684
rect 72 -1700 73 -1692
rect 88 -1700 101 -1692
rect 72 -1708 88 -1700
rect 69 -1715 88 -1712
rect 69 -1724 91 -1715
rect 42 -1734 91 -1724
rect 42 -1740 72 -1734
rect 91 -1739 96 -1734
rect 14 -1756 88 -1740
rect 106 -1748 136 -1692
rect 171 -1702 379 -1692
rect 414 -1696 459 -1692
rect 462 -1693 463 -1692
rect 478 -1693 491 -1692
rect 197 -1732 386 -1702
rect 212 -1735 386 -1732
rect 205 -1738 386 -1735
rect 14 -1758 27 -1756
rect 42 -1758 76 -1756
rect 14 -1774 88 -1758
rect 115 -1762 128 -1748
rect 143 -1762 159 -1746
rect 205 -1751 216 -1738
rect 14 -1796 27 -1774
rect 42 -1796 72 -1774
rect 115 -1778 177 -1762
rect 205 -1769 216 -1753
rect 221 -1758 231 -1738
rect 241 -1758 255 -1738
rect 258 -1751 267 -1738
rect 283 -1751 292 -1738
rect 221 -1769 255 -1758
rect 258 -1769 267 -1753
rect 283 -1769 292 -1753
rect 299 -1758 309 -1738
rect 319 -1758 333 -1738
rect 334 -1751 345 -1738
rect 299 -1769 333 -1758
rect 334 -1769 345 -1753
rect 391 -1762 407 -1746
rect 414 -1748 444 -1696
rect 478 -1700 479 -1693
rect 463 -1708 479 -1700
rect 450 -1740 463 -1721
rect 478 -1740 508 -1724
rect 450 -1756 524 -1740
rect 450 -1758 463 -1756
rect 478 -1758 512 -1756
rect 115 -1780 128 -1778
rect 143 -1780 177 -1778
rect 115 -1796 177 -1780
rect 221 -1785 237 -1782
rect 299 -1785 329 -1774
rect 377 -1778 423 -1762
rect 450 -1774 524 -1758
rect 377 -1780 411 -1778
rect 376 -1796 423 -1780
rect 450 -1796 463 -1774
rect 478 -1796 508 -1774
rect 535 -1796 536 -1780
rect 551 -1796 564 -1636
rect 594 -1740 607 -1636
rect 652 -1658 653 -1648
rect 668 -1658 681 -1648
rect 652 -1662 681 -1658
rect 686 -1662 716 -1636
rect 734 -1650 750 -1648
rect 822 -1650 875 -1636
rect 823 -1652 887 -1650
rect 930 -1652 945 -1636
rect 994 -1639 1024 -1636
rect 994 -1642 1030 -1639
rect 960 -1650 976 -1648
rect 734 -1662 749 -1658
rect 652 -1664 749 -1662
rect 777 -1664 945 -1652
rect 961 -1662 976 -1658
rect 994 -1661 1033 -1642
rect 1052 -1648 1059 -1647
rect 1058 -1655 1059 -1648
rect 1042 -1658 1043 -1655
rect 1058 -1658 1071 -1655
rect 994 -1662 1024 -1661
rect 1033 -1662 1039 -1661
rect 1042 -1662 1071 -1658
rect 961 -1663 1071 -1662
rect 961 -1664 1077 -1663
rect 636 -1672 687 -1664
rect 636 -1684 661 -1672
rect 668 -1684 687 -1672
rect 718 -1672 768 -1664
rect 718 -1680 734 -1672
rect 741 -1674 768 -1672
rect 777 -1674 998 -1664
rect 741 -1684 998 -1674
rect 1027 -1672 1077 -1664
rect 1027 -1681 1043 -1672
rect 636 -1692 687 -1684
rect 734 -1692 998 -1684
rect 1024 -1684 1043 -1681
rect 1050 -1684 1077 -1672
rect 1024 -1692 1077 -1684
rect 652 -1700 653 -1692
rect 668 -1700 681 -1692
rect 652 -1708 668 -1700
rect 649 -1715 668 -1712
rect 649 -1724 671 -1715
rect 622 -1734 671 -1724
rect 622 -1740 652 -1734
rect 671 -1739 676 -1734
rect 594 -1756 668 -1740
rect 686 -1748 716 -1692
rect 751 -1702 959 -1692
rect 994 -1696 1039 -1692
rect 1042 -1693 1043 -1692
rect 1058 -1693 1071 -1692
rect 777 -1732 966 -1702
rect 792 -1735 966 -1732
rect 785 -1738 966 -1735
rect 594 -1758 607 -1756
rect 622 -1758 656 -1756
rect 594 -1774 668 -1758
rect 695 -1762 708 -1748
rect 723 -1762 739 -1746
rect 785 -1751 796 -1738
rect 578 -1796 579 -1780
rect 594 -1796 607 -1774
rect 622 -1796 652 -1774
rect 695 -1778 757 -1762
rect 785 -1769 796 -1753
rect 801 -1758 811 -1738
rect 821 -1758 835 -1738
rect 838 -1751 847 -1738
rect 863 -1751 872 -1738
rect 801 -1769 835 -1758
rect 838 -1769 847 -1753
rect 863 -1769 872 -1753
rect 879 -1758 889 -1738
rect 899 -1758 913 -1738
rect 914 -1751 925 -1738
rect 879 -1769 913 -1758
rect 914 -1769 925 -1753
rect 971 -1762 987 -1746
rect 994 -1748 1024 -1696
rect 1058 -1700 1059 -1693
rect 1043 -1708 1059 -1700
rect 1030 -1740 1043 -1721
rect 1058 -1740 1088 -1724
rect 1030 -1756 1104 -1740
rect 1030 -1758 1043 -1756
rect 1058 -1758 1092 -1756
rect 695 -1780 708 -1778
rect 723 -1780 757 -1778
rect 695 -1796 757 -1780
rect 801 -1785 817 -1782
rect 879 -1785 909 -1774
rect 957 -1778 1003 -1762
rect 1030 -1774 1104 -1758
rect 957 -1780 991 -1778
rect 956 -1796 1003 -1780
rect 1030 -1796 1043 -1774
rect 1058 -1796 1088 -1774
rect 1115 -1796 1116 -1780
rect 1131 -1796 1144 -1636
rect 1174 -1740 1187 -1636
rect 1232 -1658 1233 -1648
rect 1248 -1658 1261 -1648
rect 1232 -1662 1261 -1658
rect 1266 -1662 1296 -1636
rect 1314 -1650 1330 -1648
rect 1402 -1650 1455 -1636
rect 1403 -1652 1467 -1650
rect 1510 -1652 1525 -1636
rect 1574 -1639 1604 -1636
rect 1574 -1642 1610 -1639
rect 1540 -1650 1556 -1648
rect 1314 -1662 1329 -1658
rect 1232 -1664 1329 -1662
rect 1357 -1664 1525 -1652
rect 1541 -1662 1556 -1658
rect 1574 -1661 1613 -1642
rect 1632 -1648 1639 -1647
rect 1638 -1655 1639 -1648
rect 1622 -1658 1623 -1655
rect 1638 -1658 1651 -1655
rect 1574 -1662 1604 -1661
rect 1613 -1662 1619 -1661
rect 1622 -1662 1651 -1658
rect 1541 -1663 1651 -1662
rect 1541 -1664 1657 -1663
rect 1216 -1672 1267 -1664
rect 1216 -1684 1241 -1672
rect 1248 -1684 1267 -1672
rect 1298 -1672 1348 -1664
rect 1298 -1680 1314 -1672
rect 1321 -1674 1348 -1672
rect 1357 -1674 1578 -1664
rect 1321 -1684 1578 -1674
rect 1607 -1672 1657 -1664
rect 1607 -1681 1623 -1672
rect 1216 -1692 1267 -1684
rect 1314 -1692 1578 -1684
rect 1604 -1684 1623 -1681
rect 1630 -1684 1657 -1672
rect 1604 -1692 1657 -1684
rect 1232 -1700 1233 -1692
rect 1248 -1700 1261 -1692
rect 1232 -1708 1248 -1700
rect 1229 -1715 1248 -1712
rect 1229 -1724 1251 -1715
rect 1202 -1734 1251 -1724
rect 1202 -1740 1232 -1734
rect 1251 -1739 1256 -1734
rect 1174 -1756 1248 -1740
rect 1266 -1748 1296 -1692
rect 1331 -1702 1539 -1692
rect 1574 -1696 1619 -1692
rect 1622 -1693 1623 -1692
rect 1638 -1693 1651 -1692
rect 1357 -1732 1546 -1702
rect 1372 -1735 1546 -1732
rect 1365 -1738 1546 -1735
rect 1174 -1758 1187 -1756
rect 1202 -1758 1236 -1756
rect 1174 -1774 1248 -1758
rect 1275 -1762 1288 -1748
rect 1303 -1762 1319 -1746
rect 1365 -1751 1376 -1738
rect 1158 -1796 1159 -1780
rect 1174 -1796 1187 -1774
rect 1202 -1796 1232 -1774
rect 1275 -1778 1337 -1762
rect 1365 -1769 1376 -1753
rect 1381 -1758 1391 -1738
rect 1401 -1758 1415 -1738
rect 1418 -1751 1427 -1738
rect 1443 -1751 1452 -1738
rect 1381 -1769 1415 -1758
rect 1418 -1769 1427 -1753
rect 1443 -1769 1452 -1753
rect 1459 -1758 1469 -1738
rect 1479 -1758 1493 -1738
rect 1494 -1751 1505 -1738
rect 1459 -1769 1493 -1758
rect 1494 -1769 1505 -1753
rect 1551 -1762 1567 -1746
rect 1574 -1748 1604 -1696
rect 1638 -1700 1639 -1693
rect 1623 -1708 1639 -1700
rect 1610 -1740 1623 -1721
rect 1638 -1740 1668 -1724
rect 1610 -1756 1684 -1740
rect 1610 -1758 1623 -1756
rect 1638 -1758 1672 -1756
rect 1275 -1780 1288 -1778
rect 1303 -1780 1337 -1778
rect 1275 -1796 1337 -1780
rect 1381 -1785 1397 -1782
rect 1459 -1785 1489 -1774
rect 1537 -1778 1583 -1762
rect 1610 -1774 1684 -1758
rect 1537 -1780 1571 -1778
rect 1536 -1796 1583 -1780
rect 1610 -1796 1623 -1774
rect 1638 -1796 1668 -1774
rect 1695 -1796 1696 -1780
rect 1711 -1796 1724 -1636
rect 1754 -1740 1767 -1636
rect 1812 -1658 1813 -1648
rect 1828 -1658 1841 -1648
rect 1812 -1662 1841 -1658
rect 1846 -1662 1876 -1636
rect 1894 -1650 1910 -1648
rect 1982 -1650 2035 -1636
rect 1983 -1652 2047 -1650
rect 2090 -1652 2105 -1636
rect 2154 -1639 2184 -1636
rect 2154 -1642 2190 -1639
rect 2120 -1650 2136 -1648
rect 1894 -1662 1909 -1658
rect 1812 -1664 1909 -1662
rect 1937 -1664 2105 -1652
rect 2121 -1662 2136 -1658
rect 2154 -1661 2193 -1642
rect 2212 -1648 2219 -1647
rect 2218 -1655 2219 -1648
rect 2202 -1658 2203 -1655
rect 2218 -1658 2231 -1655
rect 2154 -1662 2184 -1661
rect 2193 -1662 2199 -1661
rect 2202 -1662 2231 -1658
rect 2121 -1663 2231 -1662
rect 2121 -1664 2237 -1663
rect 1796 -1672 1847 -1664
rect 1796 -1684 1821 -1672
rect 1828 -1684 1847 -1672
rect 1878 -1672 1928 -1664
rect 1878 -1680 1894 -1672
rect 1901 -1674 1928 -1672
rect 1937 -1674 2158 -1664
rect 1901 -1684 2158 -1674
rect 2187 -1672 2237 -1664
rect 2187 -1681 2203 -1672
rect 1796 -1692 1847 -1684
rect 1894 -1692 2158 -1684
rect 2184 -1684 2203 -1681
rect 2210 -1684 2237 -1672
rect 2184 -1692 2237 -1684
rect 1812 -1700 1813 -1692
rect 1828 -1700 1841 -1692
rect 1812 -1708 1828 -1700
rect 1809 -1715 1828 -1712
rect 1809 -1724 1831 -1715
rect 1782 -1734 1831 -1724
rect 1782 -1740 1812 -1734
rect 1831 -1739 1836 -1734
rect 1754 -1756 1828 -1740
rect 1846 -1748 1876 -1692
rect 1911 -1702 2119 -1692
rect 2154 -1696 2199 -1692
rect 2202 -1693 2203 -1692
rect 2218 -1693 2231 -1692
rect 1937 -1732 2126 -1702
rect 1952 -1735 2126 -1732
rect 1945 -1738 2126 -1735
rect 1754 -1758 1767 -1756
rect 1782 -1758 1816 -1756
rect 1754 -1774 1828 -1758
rect 1855 -1762 1868 -1748
rect 1883 -1762 1899 -1746
rect 1945 -1751 1956 -1738
rect 1738 -1796 1739 -1780
rect 1754 -1796 1767 -1774
rect 1782 -1796 1812 -1774
rect 1855 -1778 1917 -1762
rect 1945 -1769 1956 -1753
rect 1961 -1758 1971 -1738
rect 1981 -1758 1995 -1738
rect 1998 -1751 2007 -1738
rect 2023 -1751 2032 -1738
rect 1961 -1769 1995 -1758
rect 1998 -1769 2007 -1753
rect 2023 -1769 2032 -1753
rect 2039 -1758 2049 -1738
rect 2059 -1758 2073 -1738
rect 2074 -1751 2085 -1738
rect 2039 -1769 2073 -1758
rect 2074 -1769 2085 -1753
rect 2131 -1762 2147 -1746
rect 2154 -1748 2184 -1696
rect 2218 -1700 2219 -1693
rect 2203 -1708 2219 -1700
rect 2190 -1740 2203 -1721
rect 2218 -1740 2248 -1724
rect 2190 -1756 2264 -1740
rect 2190 -1758 2203 -1756
rect 2218 -1758 2252 -1756
rect 1855 -1780 1868 -1778
rect 1883 -1780 1917 -1778
rect 1855 -1796 1917 -1780
rect 1961 -1785 1977 -1782
rect 2039 -1785 2069 -1774
rect 2117 -1778 2163 -1762
rect 2190 -1774 2264 -1758
rect 2117 -1780 2151 -1778
rect 2116 -1796 2163 -1780
rect 2190 -1796 2203 -1774
rect 2218 -1796 2248 -1774
rect 2275 -1796 2276 -1780
rect 2291 -1796 2304 -1636
rect 2334 -1740 2347 -1636
rect 2392 -1658 2393 -1648
rect 2408 -1658 2421 -1648
rect 2392 -1662 2421 -1658
rect 2426 -1662 2456 -1636
rect 2474 -1650 2490 -1648
rect 2562 -1650 2615 -1636
rect 2563 -1652 2627 -1650
rect 2670 -1652 2685 -1636
rect 2734 -1639 2764 -1636
rect 2734 -1642 2770 -1639
rect 2700 -1650 2716 -1648
rect 2474 -1662 2489 -1658
rect 2392 -1664 2489 -1662
rect 2517 -1664 2685 -1652
rect 2701 -1662 2716 -1658
rect 2734 -1661 2773 -1642
rect 2792 -1648 2799 -1647
rect 2798 -1655 2799 -1648
rect 2782 -1658 2783 -1655
rect 2798 -1658 2811 -1655
rect 2734 -1662 2764 -1661
rect 2773 -1662 2779 -1661
rect 2782 -1662 2811 -1658
rect 2701 -1663 2811 -1662
rect 2701 -1664 2817 -1663
rect 2376 -1672 2427 -1664
rect 2376 -1684 2401 -1672
rect 2408 -1684 2427 -1672
rect 2458 -1672 2508 -1664
rect 2458 -1680 2474 -1672
rect 2481 -1674 2508 -1672
rect 2517 -1674 2738 -1664
rect 2481 -1684 2738 -1674
rect 2767 -1672 2817 -1664
rect 2767 -1681 2783 -1672
rect 2376 -1692 2427 -1684
rect 2474 -1692 2738 -1684
rect 2764 -1684 2783 -1681
rect 2790 -1684 2817 -1672
rect 2764 -1692 2817 -1684
rect 2392 -1700 2393 -1692
rect 2408 -1700 2421 -1692
rect 2392 -1708 2408 -1700
rect 2389 -1715 2408 -1712
rect 2389 -1724 2411 -1715
rect 2362 -1734 2411 -1724
rect 2362 -1740 2392 -1734
rect 2411 -1739 2416 -1734
rect 2334 -1756 2408 -1740
rect 2426 -1748 2456 -1692
rect 2491 -1702 2699 -1692
rect 2734 -1696 2779 -1692
rect 2782 -1693 2783 -1692
rect 2798 -1693 2811 -1692
rect 2517 -1732 2706 -1702
rect 2532 -1735 2706 -1732
rect 2525 -1738 2706 -1735
rect 2334 -1758 2347 -1756
rect 2362 -1758 2396 -1756
rect 2334 -1774 2408 -1758
rect 2435 -1762 2448 -1748
rect 2463 -1762 2479 -1746
rect 2525 -1751 2536 -1738
rect 2318 -1796 2319 -1780
rect 2334 -1796 2347 -1774
rect 2362 -1796 2392 -1774
rect 2435 -1778 2497 -1762
rect 2525 -1769 2536 -1753
rect 2541 -1758 2551 -1738
rect 2561 -1758 2575 -1738
rect 2578 -1751 2587 -1738
rect 2603 -1751 2612 -1738
rect 2541 -1769 2575 -1758
rect 2578 -1769 2587 -1753
rect 2603 -1769 2612 -1753
rect 2619 -1758 2629 -1738
rect 2639 -1758 2653 -1738
rect 2654 -1751 2665 -1738
rect 2619 -1769 2653 -1758
rect 2654 -1769 2665 -1753
rect 2711 -1762 2727 -1746
rect 2734 -1748 2764 -1696
rect 2798 -1700 2799 -1693
rect 2783 -1708 2799 -1700
rect 2770 -1740 2783 -1721
rect 2798 -1740 2828 -1724
rect 2770 -1756 2844 -1740
rect 2770 -1758 2783 -1756
rect 2798 -1758 2832 -1756
rect 2435 -1780 2448 -1778
rect 2463 -1780 2497 -1778
rect 2435 -1796 2497 -1780
rect 2541 -1785 2557 -1782
rect 2619 -1785 2649 -1774
rect 2697 -1778 2743 -1762
rect 2770 -1774 2844 -1758
rect 2697 -1780 2731 -1778
rect 2696 -1796 2743 -1780
rect 2770 -1796 2783 -1774
rect 2798 -1796 2828 -1774
rect 2855 -1796 2856 -1780
rect 2871 -1796 2884 -1636
rect 2914 -1740 2927 -1636
rect 2972 -1658 2973 -1648
rect 2988 -1658 3001 -1648
rect 2972 -1662 3001 -1658
rect 3006 -1662 3036 -1636
rect 3054 -1650 3070 -1648
rect 3142 -1650 3195 -1636
rect 3143 -1652 3205 -1650
rect 3250 -1652 3265 -1636
rect 3314 -1639 3344 -1636
rect 3314 -1642 3350 -1639
rect 3280 -1650 3296 -1648
rect 3054 -1662 3069 -1658
rect 2972 -1664 3069 -1662
rect 3097 -1664 3265 -1652
rect 3281 -1662 3296 -1658
rect 3314 -1661 3353 -1642
rect 3372 -1648 3379 -1647
rect 3378 -1655 3379 -1648
rect 3362 -1658 3363 -1655
rect 3378 -1658 3391 -1655
rect 3314 -1662 3344 -1661
rect 3353 -1662 3359 -1661
rect 3362 -1662 3391 -1658
rect 3281 -1663 3391 -1662
rect 3281 -1664 3397 -1663
rect 2956 -1672 3007 -1664
rect 2956 -1684 2981 -1672
rect 2988 -1684 3007 -1672
rect 3038 -1672 3088 -1664
rect 3038 -1680 3054 -1672
rect 3061 -1674 3088 -1672
rect 3097 -1674 3318 -1664
rect 3061 -1684 3318 -1674
rect 3347 -1672 3397 -1664
rect 3347 -1681 3363 -1672
rect 2956 -1692 3007 -1684
rect 3054 -1692 3318 -1684
rect 3344 -1684 3363 -1681
rect 3370 -1684 3397 -1672
rect 3344 -1692 3397 -1684
rect 2972 -1700 2973 -1692
rect 2988 -1700 3001 -1692
rect 2972 -1708 2988 -1700
rect 2969 -1715 2988 -1712
rect 2969 -1724 2991 -1715
rect 2942 -1734 2991 -1724
rect 2942 -1740 2972 -1734
rect 2991 -1739 2996 -1734
rect 2914 -1756 2988 -1740
rect 3006 -1748 3036 -1692
rect 3071 -1702 3279 -1692
rect 3314 -1696 3359 -1692
rect 3362 -1693 3363 -1692
rect 3378 -1693 3391 -1692
rect 3097 -1732 3286 -1702
rect 3112 -1735 3286 -1732
rect 3105 -1738 3286 -1735
rect 2914 -1758 2927 -1756
rect 2942 -1758 2976 -1756
rect 2914 -1774 2988 -1758
rect 3015 -1762 3028 -1748
rect 3043 -1762 3059 -1746
rect 3105 -1751 3116 -1738
rect 2898 -1796 2899 -1780
rect 2914 -1796 2927 -1774
rect 2942 -1796 2972 -1774
rect 3015 -1778 3077 -1762
rect 3105 -1769 3116 -1753
rect 3121 -1758 3131 -1738
rect 3141 -1758 3155 -1738
rect 3158 -1751 3167 -1738
rect 3183 -1751 3192 -1738
rect 3121 -1769 3155 -1758
rect 3158 -1769 3167 -1753
rect 3183 -1769 3192 -1753
rect 3199 -1758 3209 -1738
rect 3219 -1758 3233 -1738
rect 3234 -1751 3245 -1738
rect 3199 -1769 3233 -1758
rect 3234 -1769 3245 -1753
rect 3291 -1762 3307 -1746
rect 3314 -1748 3344 -1696
rect 3378 -1700 3379 -1693
rect 3363 -1708 3379 -1700
rect 3350 -1740 3363 -1721
rect 3378 -1740 3408 -1724
rect 3350 -1756 3424 -1740
rect 3350 -1758 3363 -1756
rect 3378 -1758 3412 -1756
rect 3015 -1780 3028 -1778
rect 3043 -1780 3077 -1778
rect 3015 -1796 3077 -1780
rect 3121 -1785 3137 -1782
rect 3199 -1785 3229 -1774
rect 3277 -1778 3323 -1762
rect 3350 -1774 3424 -1758
rect 3277 -1780 3311 -1778
rect 3276 -1796 3323 -1780
rect 3350 -1796 3363 -1774
rect 3378 -1796 3408 -1774
rect 3435 -1796 3436 -1780
rect 3451 -1796 3464 -1636
rect 3494 -1740 3507 -1636
rect 3552 -1658 3553 -1648
rect 3568 -1658 3581 -1648
rect 3552 -1662 3581 -1658
rect 3586 -1662 3616 -1636
rect 3634 -1650 3650 -1648
rect 3722 -1650 3775 -1636
rect 3723 -1652 3787 -1650
rect 3830 -1652 3845 -1636
rect 3894 -1639 3924 -1636
rect 3894 -1642 3930 -1639
rect 3860 -1650 3876 -1648
rect 3634 -1662 3649 -1658
rect 3552 -1664 3649 -1662
rect 3677 -1664 3845 -1652
rect 3861 -1662 3876 -1658
rect 3894 -1661 3933 -1642
rect 3952 -1648 3959 -1647
rect 3958 -1655 3959 -1648
rect 3942 -1658 3943 -1655
rect 3958 -1658 3971 -1655
rect 3894 -1662 3924 -1661
rect 3933 -1662 3939 -1661
rect 3942 -1662 3971 -1658
rect 3861 -1663 3971 -1662
rect 3861 -1664 3977 -1663
rect 3536 -1672 3587 -1664
rect 3536 -1684 3561 -1672
rect 3568 -1684 3587 -1672
rect 3618 -1672 3668 -1664
rect 3618 -1680 3634 -1672
rect 3641 -1674 3668 -1672
rect 3677 -1674 3898 -1664
rect 3641 -1684 3898 -1674
rect 3927 -1672 3977 -1664
rect 3927 -1681 3943 -1672
rect 3536 -1692 3587 -1684
rect 3634 -1692 3898 -1684
rect 3924 -1684 3943 -1681
rect 3950 -1684 3977 -1672
rect 3924 -1692 3977 -1684
rect 3552 -1700 3553 -1692
rect 3568 -1700 3581 -1692
rect 3552 -1708 3568 -1700
rect 3549 -1715 3568 -1712
rect 3549 -1724 3571 -1715
rect 3522 -1734 3571 -1724
rect 3522 -1740 3552 -1734
rect 3571 -1739 3576 -1734
rect 3494 -1756 3568 -1740
rect 3586 -1748 3616 -1692
rect 3651 -1702 3859 -1692
rect 3894 -1696 3939 -1692
rect 3942 -1693 3943 -1692
rect 3958 -1693 3971 -1692
rect 3677 -1732 3866 -1702
rect 3692 -1735 3866 -1732
rect 3685 -1738 3866 -1735
rect 3494 -1758 3507 -1756
rect 3522 -1758 3556 -1756
rect 3494 -1774 3568 -1758
rect 3595 -1762 3608 -1748
rect 3623 -1762 3639 -1746
rect 3685 -1751 3696 -1738
rect 3478 -1796 3479 -1780
rect 3494 -1796 3507 -1774
rect 3522 -1796 3552 -1774
rect 3595 -1778 3657 -1762
rect 3685 -1769 3696 -1753
rect 3701 -1758 3711 -1738
rect 3721 -1758 3735 -1738
rect 3738 -1751 3747 -1738
rect 3763 -1751 3772 -1738
rect 3701 -1769 3735 -1758
rect 3738 -1769 3747 -1753
rect 3763 -1769 3772 -1753
rect 3779 -1758 3789 -1738
rect 3799 -1758 3813 -1738
rect 3814 -1751 3825 -1738
rect 3779 -1769 3813 -1758
rect 3814 -1769 3825 -1753
rect 3871 -1762 3887 -1746
rect 3894 -1748 3924 -1696
rect 3958 -1700 3959 -1693
rect 3943 -1708 3959 -1700
rect 3930 -1740 3943 -1721
rect 3958 -1740 3988 -1724
rect 3930 -1756 4004 -1740
rect 3930 -1758 3943 -1756
rect 3958 -1758 3992 -1756
rect 3595 -1780 3608 -1778
rect 3623 -1780 3657 -1778
rect 3595 -1796 3657 -1780
rect 3701 -1785 3717 -1782
rect 3779 -1785 3809 -1774
rect 3857 -1778 3903 -1762
rect 3930 -1774 4004 -1758
rect 3857 -1780 3891 -1778
rect 3856 -1796 3903 -1780
rect 3930 -1796 3943 -1774
rect 3958 -1796 3988 -1774
rect 4015 -1796 4016 -1780
rect 4031 -1796 4044 -1636
rect 4074 -1740 4087 -1636
rect 4132 -1658 4133 -1648
rect 4148 -1658 4161 -1648
rect 4132 -1662 4161 -1658
rect 4166 -1662 4196 -1636
rect 4214 -1650 4230 -1648
rect 4302 -1650 4355 -1636
rect 4303 -1652 4367 -1650
rect 4410 -1652 4425 -1636
rect 4474 -1639 4504 -1636
rect 4611 -1637 6944 -1636
rect 4474 -1642 4510 -1639
rect 4440 -1650 4456 -1648
rect 4214 -1662 4229 -1658
rect 4132 -1664 4229 -1662
rect 4257 -1664 4425 -1652
rect 4441 -1662 4456 -1658
rect 4474 -1661 4513 -1642
rect 4532 -1648 4539 -1647
rect 4538 -1655 4539 -1648
rect 4522 -1658 4523 -1655
rect 4538 -1658 4551 -1655
rect 4474 -1662 4504 -1661
rect 4513 -1662 4519 -1661
rect 4522 -1662 4551 -1658
rect 4441 -1663 4551 -1662
rect 4441 -1664 4557 -1663
rect 4116 -1672 4167 -1664
rect 4116 -1684 4141 -1672
rect 4148 -1684 4167 -1672
rect 4198 -1672 4248 -1664
rect 4198 -1680 4214 -1672
rect 4221 -1674 4248 -1672
rect 4257 -1674 4478 -1664
rect 4221 -1684 4478 -1674
rect 4507 -1672 4557 -1664
rect 4507 -1681 4523 -1672
rect 4116 -1692 4167 -1684
rect 4214 -1692 4478 -1684
rect 4504 -1684 4523 -1681
rect 4530 -1684 4557 -1672
rect 4504 -1692 4557 -1684
rect 4132 -1700 4133 -1692
rect 4148 -1700 4161 -1692
rect 4132 -1708 4148 -1700
rect 4129 -1715 4148 -1712
rect 4129 -1724 4151 -1715
rect 4102 -1734 4151 -1724
rect 4102 -1740 4132 -1734
rect 4151 -1739 4156 -1734
rect 4074 -1756 4148 -1740
rect 4166 -1748 4196 -1692
rect 4231 -1702 4439 -1692
rect 4474 -1696 4519 -1692
rect 4522 -1693 4523 -1692
rect 4538 -1693 4551 -1692
rect 4257 -1732 4446 -1702
rect 4272 -1735 4446 -1732
rect 4265 -1738 4446 -1735
rect 4074 -1758 4087 -1756
rect 4102 -1758 4136 -1756
rect 4074 -1774 4148 -1758
rect 4175 -1762 4188 -1748
rect 4203 -1762 4219 -1746
rect 4265 -1751 4276 -1738
rect 4058 -1796 4059 -1780
rect 4074 -1796 4087 -1774
rect 4102 -1796 4132 -1774
rect 4175 -1778 4237 -1762
rect 4265 -1769 4276 -1753
rect 4281 -1758 4291 -1738
rect 4301 -1758 4315 -1738
rect 4318 -1751 4327 -1738
rect 4343 -1751 4352 -1738
rect 4281 -1769 4315 -1758
rect 4318 -1769 4327 -1753
rect 4343 -1769 4352 -1753
rect 4359 -1758 4369 -1738
rect 4379 -1758 4393 -1738
rect 4394 -1751 4405 -1738
rect 4359 -1769 4393 -1758
rect 4394 -1769 4405 -1753
rect 4451 -1762 4467 -1746
rect 4474 -1748 4504 -1696
rect 4538 -1700 4539 -1693
rect 4523 -1708 4539 -1700
rect 4510 -1740 4523 -1721
rect 4538 -1740 4568 -1724
rect 4510 -1756 4584 -1740
rect 4510 -1758 4523 -1756
rect 4538 -1758 4572 -1756
rect 4175 -1780 4188 -1778
rect 4203 -1780 4237 -1778
rect 4175 -1796 4237 -1780
rect 4281 -1785 4297 -1782
rect 4359 -1785 4389 -1774
rect 4437 -1778 4483 -1762
rect 4510 -1774 4584 -1758
rect 4437 -1780 4471 -1778
rect 4436 -1796 4483 -1780
rect 4510 -1796 4523 -1774
rect 4538 -1796 4568 -1774
rect 4595 -1796 4596 -1780
rect 4611 -1796 4624 -1637
rect 4654 -1741 4667 -1637
rect 4712 -1659 4713 -1649
rect 4733 -1651 4741 -1649
rect 4731 -1653 4741 -1651
rect 4729 -1655 4741 -1653
rect 4728 -1659 4741 -1655
rect 4712 -1663 4741 -1659
rect 4746 -1663 4776 -1637
rect 4794 -1651 4810 -1649
rect 4882 -1651 4933 -1637
rect 4883 -1653 4947 -1651
rect 4990 -1653 5005 -1637
rect 5054 -1640 5084 -1637
rect 5054 -1643 5090 -1640
rect 5020 -1651 5036 -1649
rect 4794 -1663 4809 -1659
rect 4712 -1665 4809 -1663
rect 4837 -1665 5005 -1653
rect 5021 -1663 5036 -1659
rect 5054 -1662 5093 -1643
rect 5112 -1649 5119 -1648
rect 5118 -1656 5119 -1649
rect 5102 -1659 5103 -1656
rect 5118 -1659 5131 -1656
rect 5054 -1663 5084 -1662
rect 5093 -1663 5099 -1662
rect 5102 -1663 5131 -1659
rect 5021 -1664 5131 -1663
rect 5021 -1665 5137 -1664
rect 4696 -1673 4747 -1665
rect 4696 -1685 4721 -1673
rect 4728 -1685 4747 -1673
rect 4778 -1673 4828 -1665
rect 4778 -1681 4794 -1673
rect 4801 -1675 4828 -1673
rect 4837 -1675 5058 -1665
rect 4801 -1685 5058 -1675
rect 5087 -1673 5137 -1665
rect 5087 -1682 5103 -1673
rect 4696 -1693 4747 -1685
rect 4794 -1693 5058 -1685
rect 5084 -1685 5103 -1682
rect 5110 -1685 5137 -1673
rect 5084 -1693 5137 -1685
rect 4712 -1701 4713 -1693
rect 4728 -1701 4741 -1693
rect 4712 -1709 4728 -1701
rect 4709 -1716 4728 -1713
rect 4709 -1725 4731 -1716
rect 4682 -1735 4731 -1725
rect 4682 -1741 4712 -1735
rect 4731 -1740 4736 -1735
rect 4654 -1757 4728 -1741
rect 4746 -1749 4776 -1693
rect 4811 -1703 5019 -1693
rect 5054 -1697 5099 -1693
rect 5102 -1694 5103 -1693
rect 5118 -1694 5131 -1693
rect 4837 -1733 5026 -1703
rect 4852 -1736 5026 -1733
rect 4845 -1739 5026 -1736
rect 4654 -1759 4667 -1757
rect 4682 -1759 4716 -1757
rect 4654 -1775 4728 -1759
rect 4755 -1763 4768 -1749
rect 4783 -1763 4799 -1747
rect 4845 -1752 4856 -1739
rect 0 -1804 33 -1796
rect 0 -1830 7 -1804
rect 14 -1830 33 -1804
rect 97 -1808 159 -1796
rect 171 -1808 246 -1796
rect 304 -1808 379 -1796
rect 391 -1808 422 -1796
rect 428 -1808 463 -1796
rect 97 -1810 259 -1808
rect 0 -1838 33 -1830
rect 115 -1834 128 -1810
rect 143 -1812 158 -1810
rect 14 -1848 27 -1838
rect 42 -1848 72 -1834
rect 115 -1848 158 -1834
rect 182 -1837 189 -1830
rect 192 -1834 259 -1810
rect 291 -1810 463 -1808
rect 261 -1832 289 -1828
rect 291 -1832 371 -1810
rect 392 -1812 407 -1810
rect 261 -1834 371 -1832
rect 192 -1838 371 -1834
rect 165 -1848 195 -1838
rect 197 -1848 350 -1838
rect 358 -1848 388 -1838
rect 392 -1848 422 -1834
rect 450 -1848 463 -1810
rect 535 -1804 570 -1796
rect 535 -1830 536 -1804
rect 543 -1830 570 -1804
rect 478 -1848 508 -1834
rect 535 -1838 570 -1830
rect 572 -1804 613 -1796
rect 572 -1830 587 -1804
rect 594 -1830 613 -1804
rect 677 -1808 739 -1796
rect 751 -1808 826 -1796
rect 884 -1808 959 -1796
rect 971 -1808 1002 -1796
rect 1008 -1808 1043 -1796
rect 677 -1810 839 -1808
rect 572 -1838 613 -1830
rect 695 -1834 708 -1810
rect 723 -1812 738 -1810
rect 535 -1848 536 -1838
rect 551 -1848 564 -1838
rect 578 -1848 579 -1838
rect 594 -1848 607 -1838
rect 622 -1848 652 -1834
rect 695 -1848 738 -1834
rect 762 -1837 769 -1830
rect 772 -1834 839 -1810
rect 871 -1810 1043 -1808
rect 841 -1832 869 -1828
rect 871 -1832 951 -1810
rect 972 -1812 987 -1810
rect 841 -1834 951 -1832
rect 772 -1838 951 -1834
rect 745 -1848 775 -1838
rect 777 -1848 930 -1838
rect 938 -1848 968 -1838
rect 972 -1848 1002 -1834
rect 1030 -1848 1043 -1810
rect 1115 -1804 1150 -1796
rect 1115 -1830 1116 -1804
rect 1123 -1830 1150 -1804
rect 1058 -1848 1088 -1834
rect 1115 -1838 1150 -1830
rect 1152 -1804 1193 -1796
rect 1152 -1830 1167 -1804
rect 1174 -1830 1193 -1804
rect 1257 -1808 1319 -1796
rect 1331 -1808 1406 -1796
rect 1464 -1808 1539 -1796
rect 1551 -1808 1582 -1796
rect 1588 -1808 1623 -1796
rect 1257 -1810 1419 -1808
rect 1152 -1838 1193 -1830
rect 1275 -1834 1288 -1810
rect 1303 -1812 1318 -1810
rect 1115 -1848 1116 -1838
rect 1131 -1848 1144 -1838
rect 1158 -1848 1159 -1838
rect 1174 -1848 1187 -1838
rect 1202 -1848 1232 -1834
rect 1275 -1848 1318 -1834
rect 1342 -1837 1349 -1830
rect 1352 -1834 1419 -1810
rect 1451 -1810 1623 -1808
rect 1421 -1832 1449 -1828
rect 1451 -1832 1531 -1810
rect 1552 -1812 1567 -1810
rect 1421 -1834 1531 -1832
rect 1352 -1838 1531 -1834
rect 1325 -1848 1355 -1838
rect 1357 -1848 1510 -1838
rect 1518 -1848 1548 -1838
rect 1552 -1848 1582 -1834
rect 1610 -1848 1623 -1810
rect 1695 -1804 1730 -1796
rect 1695 -1830 1696 -1804
rect 1703 -1830 1730 -1804
rect 1638 -1848 1668 -1834
rect 1695 -1838 1730 -1830
rect 1732 -1804 1773 -1796
rect 1732 -1830 1747 -1804
rect 1754 -1830 1773 -1804
rect 1837 -1808 1899 -1796
rect 1911 -1808 1986 -1796
rect 2044 -1808 2119 -1796
rect 2131 -1808 2162 -1796
rect 2168 -1808 2203 -1796
rect 1837 -1810 1999 -1808
rect 1732 -1838 1773 -1830
rect 1855 -1834 1868 -1810
rect 1883 -1812 1898 -1810
rect 1695 -1848 1696 -1838
rect 1711 -1848 1724 -1838
rect 1738 -1848 1739 -1838
rect 1754 -1848 1767 -1838
rect 1782 -1848 1812 -1834
rect 1855 -1848 1898 -1834
rect 1922 -1837 1929 -1830
rect 1932 -1834 1999 -1810
rect 2031 -1810 2203 -1808
rect 2001 -1832 2029 -1828
rect 2031 -1832 2111 -1810
rect 2132 -1812 2147 -1810
rect 2001 -1834 2111 -1832
rect 1932 -1838 2111 -1834
rect 1905 -1848 1935 -1838
rect 1937 -1848 2090 -1838
rect 2098 -1848 2128 -1838
rect 2132 -1848 2162 -1834
rect 2190 -1848 2203 -1810
rect 2275 -1804 2310 -1796
rect 2275 -1830 2276 -1804
rect 2283 -1830 2310 -1804
rect 2218 -1848 2248 -1834
rect 2275 -1838 2310 -1830
rect 2312 -1804 2353 -1796
rect 2312 -1830 2327 -1804
rect 2334 -1830 2353 -1804
rect 2417 -1808 2479 -1796
rect 2491 -1808 2566 -1796
rect 2624 -1808 2699 -1796
rect 2711 -1808 2742 -1796
rect 2748 -1808 2783 -1796
rect 2417 -1810 2579 -1808
rect 2312 -1838 2353 -1830
rect 2435 -1834 2448 -1810
rect 2463 -1812 2478 -1810
rect 2275 -1848 2276 -1838
rect 2291 -1848 2304 -1838
rect 2318 -1848 2319 -1838
rect 2334 -1848 2347 -1838
rect 2362 -1848 2392 -1834
rect 2435 -1848 2478 -1834
rect 2502 -1837 2509 -1830
rect 2512 -1834 2579 -1810
rect 2611 -1810 2783 -1808
rect 2581 -1832 2609 -1828
rect 2611 -1832 2691 -1810
rect 2712 -1812 2727 -1810
rect 2581 -1834 2691 -1832
rect 2512 -1838 2691 -1834
rect 2485 -1848 2515 -1838
rect 2517 -1848 2670 -1838
rect 2678 -1848 2708 -1838
rect 2712 -1848 2742 -1834
rect 2770 -1848 2783 -1810
rect 2855 -1804 2890 -1796
rect 2855 -1830 2856 -1804
rect 2863 -1830 2890 -1804
rect 2798 -1848 2828 -1834
rect 2855 -1838 2890 -1830
rect 2892 -1804 2933 -1796
rect 2892 -1830 2907 -1804
rect 2914 -1830 2933 -1804
rect 2997 -1808 3059 -1796
rect 3071 -1808 3146 -1796
rect 3204 -1808 3279 -1796
rect 3291 -1808 3322 -1796
rect 3328 -1808 3363 -1796
rect 2997 -1810 3159 -1808
rect 2892 -1838 2933 -1830
rect 3015 -1834 3028 -1810
rect 3043 -1812 3058 -1810
rect 2855 -1848 2856 -1838
rect 2871 -1848 2884 -1838
rect 2898 -1848 2899 -1838
rect 2914 -1848 2927 -1838
rect 2942 -1848 2972 -1834
rect 3015 -1848 3058 -1834
rect 3082 -1837 3089 -1830
rect 3092 -1834 3159 -1810
rect 3191 -1810 3363 -1808
rect 3161 -1832 3189 -1828
rect 3191 -1832 3271 -1810
rect 3292 -1812 3307 -1810
rect 3161 -1834 3271 -1832
rect 3092 -1838 3271 -1834
rect 3065 -1848 3095 -1838
rect 3097 -1848 3250 -1838
rect 3258 -1848 3288 -1838
rect 3292 -1848 3322 -1834
rect 3350 -1848 3363 -1810
rect 3435 -1804 3470 -1796
rect 3435 -1830 3436 -1804
rect 3443 -1830 3470 -1804
rect 3378 -1848 3408 -1834
rect 3435 -1838 3470 -1830
rect 3472 -1804 3513 -1796
rect 3472 -1830 3487 -1804
rect 3494 -1830 3513 -1804
rect 3577 -1808 3639 -1796
rect 3651 -1808 3726 -1796
rect 3784 -1808 3859 -1796
rect 3871 -1808 3902 -1796
rect 3908 -1808 3943 -1796
rect 3577 -1810 3739 -1808
rect 3472 -1838 3513 -1830
rect 3595 -1834 3608 -1810
rect 3623 -1812 3638 -1810
rect 3435 -1848 3436 -1838
rect 3451 -1848 3464 -1838
rect 3478 -1848 3479 -1838
rect 3494 -1848 3507 -1838
rect 3522 -1848 3552 -1834
rect 3595 -1848 3638 -1834
rect 3662 -1837 3669 -1830
rect 3672 -1834 3739 -1810
rect 3771 -1810 3943 -1808
rect 3741 -1832 3769 -1828
rect 3771 -1832 3851 -1810
rect 3872 -1812 3887 -1810
rect 3741 -1834 3851 -1832
rect 3672 -1838 3851 -1834
rect 3645 -1848 3675 -1838
rect 3677 -1848 3830 -1838
rect 3838 -1848 3868 -1838
rect 3872 -1848 3902 -1834
rect 3930 -1848 3943 -1810
rect 4015 -1804 4050 -1796
rect 4015 -1830 4016 -1804
rect 4023 -1830 4050 -1804
rect 3958 -1848 3988 -1834
rect 4015 -1838 4050 -1830
rect 4052 -1804 4093 -1796
rect 4052 -1830 4067 -1804
rect 4074 -1830 4093 -1804
rect 4157 -1808 4219 -1796
rect 4231 -1808 4306 -1796
rect 4364 -1808 4439 -1796
rect 4451 -1808 4482 -1796
rect 4488 -1808 4523 -1796
rect 4157 -1810 4319 -1808
rect 4052 -1838 4093 -1830
rect 4175 -1834 4188 -1810
rect 4203 -1812 4218 -1810
rect 4015 -1848 4016 -1838
rect 4031 -1848 4044 -1838
rect 4058 -1848 4059 -1838
rect 4074 -1848 4087 -1838
rect 4102 -1848 4132 -1834
rect 4175 -1848 4218 -1834
rect 4242 -1837 4249 -1830
rect 4252 -1834 4319 -1810
rect 4351 -1810 4523 -1808
rect 4321 -1832 4349 -1828
rect 4351 -1832 4431 -1810
rect 4452 -1812 4467 -1810
rect 4321 -1834 4431 -1832
rect 4252 -1838 4431 -1834
rect 4225 -1848 4255 -1838
rect 4257 -1848 4410 -1838
rect 4418 -1848 4448 -1838
rect 4452 -1848 4482 -1834
rect 4510 -1848 4523 -1810
rect 4595 -1804 4630 -1796
rect 4638 -1797 4639 -1781
rect 4654 -1797 4667 -1775
rect 4682 -1797 4712 -1775
rect 4755 -1779 4817 -1763
rect 4845 -1770 4856 -1754
rect 4861 -1759 4871 -1739
rect 4881 -1759 4895 -1739
rect 4898 -1752 4907 -1739
rect 4923 -1752 4932 -1739
rect 4861 -1770 4895 -1759
rect 4898 -1770 4907 -1754
rect 4923 -1770 4932 -1754
rect 4939 -1759 4949 -1739
rect 4959 -1759 4973 -1739
rect 4974 -1752 4985 -1739
rect 4939 -1770 4973 -1759
rect 4974 -1770 4985 -1754
rect 5031 -1763 5047 -1747
rect 5054 -1749 5084 -1697
rect 5118 -1701 5119 -1694
rect 5103 -1709 5119 -1701
rect 5090 -1741 5103 -1722
rect 5118 -1741 5148 -1725
rect 5090 -1757 5164 -1741
rect 5090 -1759 5103 -1757
rect 5118 -1759 5152 -1757
rect 4755 -1781 4768 -1779
rect 4783 -1781 4817 -1779
rect 4755 -1797 4817 -1781
rect 4861 -1786 4877 -1783
rect 4939 -1786 4969 -1775
rect 5017 -1779 5063 -1763
rect 5090 -1775 5164 -1759
rect 5017 -1781 5051 -1779
rect 5016 -1797 5063 -1781
rect 5090 -1797 5103 -1775
rect 5118 -1797 5148 -1775
rect 5175 -1797 5176 -1781
rect 5191 -1797 5204 -1637
rect 5234 -1741 5247 -1637
rect 5292 -1659 5293 -1649
rect 5313 -1651 5321 -1649
rect 5311 -1653 5321 -1651
rect 5309 -1655 5321 -1653
rect 5308 -1659 5321 -1655
rect 5292 -1663 5321 -1659
rect 5326 -1663 5356 -1637
rect 5374 -1651 5390 -1649
rect 5462 -1651 5513 -1637
rect 5463 -1653 5527 -1651
rect 5570 -1653 5585 -1637
rect 5634 -1640 5664 -1637
rect 5634 -1643 5670 -1640
rect 5600 -1651 5616 -1649
rect 5374 -1663 5389 -1659
rect 5292 -1665 5389 -1663
rect 5417 -1665 5585 -1653
rect 5601 -1663 5616 -1659
rect 5634 -1662 5673 -1643
rect 5692 -1649 5699 -1648
rect 5698 -1656 5699 -1649
rect 5682 -1659 5683 -1656
rect 5698 -1659 5711 -1656
rect 5634 -1663 5664 -1662
rect 5673 -1663 5679 -1662
rect 5682 -1663 5711 -1659
rect 5601 -1664 5711 -1663
rect 5601 -1665 5717 -1664
rect 5276 -1673 5327 -1665
rect 5276 -1685 5301 -1673
rect 5308 -1685 5327 -1673
rect 5358 -1673 5408 -1665
rect 5358 -1681 5374 -1673
rect 5381 -1675 5408 -1673
rect 5417 -1675 5638 -1665
rect 5381 -1685 5638 -1675
rect 5667 -1673 5717 -1665
rect 5667 -1682 5683 -1673
rect 5276 -1693 5327 -1685
rect 5374 -1693 5638 -1685
rect 5664 -1685 5683 -1682
rect 5690 -1685 5717 -1673
rect 5664 -1693 5717 -1685
rect 5292 -1701 5293 -1693
rect 5308 -1701 5321 -1693
rect 5292 -1709 5308 -1701
rect 5289 -1716 5308 -1713
rect 5289 -1725 5311 -1716
rect 5262 -1735 5311 -1725
rect 5262 -1741 5292 -1735
rect 5311 -1740 5316 -1735
rect 5234 -1757 5308 -1741
rect 5326 -1749 5356 -1693
rect 5391 -1703 5599 -1693
rect 5634 -1697 5679 -1693
rect 5682 -1694 5683 -1693
rect 5698 -1694 5711 -1693
rect 5417 -1733 5606 -1703
rect 5432 -1736 5606 -1733
rect 5425 -1739 5606 -1736
rect 5234 -1759 5247 -1757
rect 5262 -1759 5296 -1757
rect 5234 -1775 5308 -1759
rect 5335 -1763 5348 -1749
rect 5363 -1763 5379 -1747
rect 5425 -1752 5436 -1739
rect 5218 -1797 5219 -1781
rect 5234 -1797 5247 -1775
rect 5262 -1797 5292 -1775
rect 5335 -1779 5397 -1763
rect 5425 -1770 5436 -1754
rect 5441 -1759 5451 -1739
rect 5461 -1759 5475 -1739
rect 5478 -1752 5487 -1739
rect 5503 -1752 5512 -1739
rect 5441 -1770 5475 -1759
rect 5478 -1770 5487 -1754
rect 5503 -1770 5512 -1754
rect 5519 -1759 5529 -1739
rect 5539 -1759 5553 -1739
rect 5554 -1752 5565 -1739
rect 5519 -1770 5553 -1759
rect 5554 -1770 5565 -1754
rect 5611 -1763 5627 -1747
rect 5634 -1749 5664 -1697
rect 5698 -1701 5699 -1694
rect 5683 -1709 5699 -1701
rect 5670 -1741 5683 -1722
rect 5698 -1741 5728 -1725
rect 5670 -1757 5744 -1741
rect 5670 -1759 5683 -1757
rect 5698 -1759 5732 -1757
rect 5335 -1781 5348 -1779
rect 5363 -1781 5397 -1779
rect 5335 -1797 5397 -1781
rect 5441 -1786 5457 -1783
rect 5519 -1786 5549 -1775
rect 5597 -1779 5643 -1763
rect 5670 -1775 5744 -1759
rect 5597 -1781 5631 -1779
rect 5596 -1797 5643 -1781
rect 5670 -1797 5683 -1775
rect 5698 -1797 5728 -1775
rect 5755 -1797 5756 -1781
rect 5771 -1797 5784 -1637
rect 5814 -1741 5827 -1637
rect 5872 -1659 5873 -1649
rect 5893 -1651 5901 -1649
rect 5891 -1653 5901 -1651
rect 5889 -1655 5901 -1653
rect 5888 -1659 5901 -1655
rect 5872 -1663 5901 -1659
rect 5906 -1663 5936 -1637
rect 5954 -1651 5970 -1649
rect 6042 -1651 6093 -1637
rect 6043 -1653 6107 -1651
rect 6150 -1653 6165 -1637
rect 6214 -1640 6244 -1637
rect 6214 -1643 6250 -1640
rect 6180 -1651 6196 -1649
rect 5954 -1663 5969 -1659
rect 5872 -1665 5969 -1663
rect 5997 -1665 6165 -1653
rect 6181 -1663 6196 -1659
rect 6214 -1662 6253 -1643
rect 6272 -1649 6279 -1648
rect 6278 -1656 6279 -1649
rect 6262 -1659 6263 -1656
rect 6278 -1659 6291 -1656
rect 6214 -1663 6244 -1662
rect 6253 -1663 6259 -1662
rect 6262 -1663 6291 -1659
rect 6181 -1664 6291 -1663
rect 6181 -1665 6297 -1664
rect 5856 -1673 5907 -1665
rect 5856 -1685 5881 -1673
rect 5888 -1685 5907 -1673
rect 5938 -1673 5988 -1665
rect 5938 -1681 5954 -1673
rect 5961 -1675 5988 -1673
rect 5997 -1675 6218 -1665
rect 5961 -1685 6218 -1675
rect 6247 -1673 6297 -1665
rect 6247 -1682 6263 -1673
rect 5856 -1693 5907 -1685
rect 5954 -1693 6218 -1685
rect 6244 -1685 6263 -1682
rect 6270 -1685 6297 -1673
rect 6244 -1693 6297 -1685
rect 5872 -1701 5873 -1693
rect 5888 -1701 5901 -1693
rect 5872 -1709 5888 -1701
rect 5869 -1716 5888 -1713
rect 5869 -1725 5891 -1716
rect 5842 -1735 5891 -1725
rect 5842 -1741 5872 -1735
rect 5891 -1740 5896 -1735
rect 5814 -1757 5888 -1741
rect 5906 -1749 5936 -1693
rect 5971 -1703 6179 -1693
rect 6214 -1697 6259 -1693
rect 6262 -1694 6263 -1693
rect 6278 -1694 6291 -1693
rect 5997 -1733 6186 -1703
rect 6012 -1736 6186 -1733
rect 6005 -1739 6186 -1736
rect 5814 -1759 5827 -1757
rect 5842 -1759 5876 -1757
rect 5814 -1775 5888 -1759
rect 5915 -1763 5928 -1749
rect 5943 -1763 5959 -1747
rect 6005 -1752 6016 -1739
rect 5798 -1797 5799 -1781
rect 5814 -1797 5827 -1775
rect 5842 -1797 5872 -1775
rect 5915 -1779 5977 -1763
rect 6005 -1770 6016 -1754
rect 6021 -1759 6031 -1739
rect 6041 -1759 6055 -1739
rect 6058 -1752 6067 -1739
rect 6083 -1752 6092 -1739
rect 6021 -1770 6055 -1759
rect 6058 -1770 6067 -1754
rect 6083 -1770 6092 -1754
rect 6099 -1759 6109 -1739
rect 6119 -1759 6133 -1739
rect 6134 -1752 6145 -1739
rect 6099 -1770 6133 -1759
rect 6134 -1770 6145 -1754
rect 6191 -1763 6207 -1747
rect 6214 -1749 6244 -1697
rect 6278 -1701 6279 -1694
rect 6263 -1709 6279 -1701
rect 6250 -1741 6263 -1722
rect 6278 -1741 6308 -1725
rect 6250 -1757 6324 -1741
rect 6250 -1759 6263 -1757
rect 6278 -1759 6312 -1757
rect 5915 -1781 5928 -1779
rect 5943 -1781 5977 -1779
rect 5915 -1797 5977 -1781
rect 6021 -1786 6037 -1783
rect 6099 -1786 6129 -1775
rect 6177 -1779 6223 -1763
rect 6250 -1775 6324 -1759
rect 6177 -1781 6211 -1779
rect 6176 -1797 6223 -1781
rect 6250 -1797 6263 -1775
rect 6278 -1797 6308 -1775
rect 6335 -1797 6336 -1781
rect 6351 -1797 6364 -1637
rect 6394 -1741 6407 -1637
rect 6452 -1659 6453 -1649
rect 6473 -1651 6481 -1649
rect 6471 -1653 6481 -1651
rect 6469 -1655 6481 -1653
rect 6468 -1659 6481 -1655
rect 6452 -1663 6481 -1659
rect 6486 -1663 6516 -1637
rect 6534 -1651 6550 -1649
rect 6622 -1651 6673 -1637
rect 6623 -1653 6687 -1651
rect 6730 -1653 6745 -1637
rect 6794 -1640 6824 -1637
rect 6794 -1643 6830 -1640
rect 6760 -1651 6776 -1649
rect 6534 -1663 6549 -1659
rect 6452 -1665 6549 -1663
rect 6577 -1665 6745 -1653
rect 6761 -1663 6776 -1659
rect 6794 -1662 6833 -1643
rect 6852 -1649 6859 -1648
rect 6858 -1656 6859 -1649
rect 6842 -1659 6843 -1656
rect 6858 -1659 6871 -1656
rect 6794 -1663 6824 -1662
rect 6833 -1663 6839 -1662
rect 6842 -1663 6871 -1659
rect 6761 -1664 6871 -1663
rect 6761 -1665 6877 -1664
rect 6436 -1673 6487 -1665
rect 6436 -1685 6461 -1673
rect 6468 -1685 6487 -1673
rect 6518 -1673 6568 -1665
rect 6518 -1681 6534 -1673
rect 6541 -1675 6568 -1673
rect 6577 -1675 6798 -1665
rect 6541 -1685 6798 -1675
rect 6827 -1673 6877 -1665
rect 6827 -1682 6843 -1673
rect 6436 -1693 6487 -1685
rect 6534 -1693 6798 -1685
rect 6824 -1685 6843 -1682
rect 6850 -1685 6877 -1673
rect 6824 -1693 6877 -1685
rect 6452 -1701 6453 -1693
rect 6468 -1701 6481 -1693
rect 6452 -1709 6468 -1701
rect 6449 -1716 6468 -1713
rect 6449 -1725 6471 -1716
rect 6422 -1735 6471 -1725
rect 6422 -1741 6452 -1735
rect 6471 -1740 6476 -1735
rect 6394 -1757 6468 -1741
rect 6486 -1749 6516 -1693
rect 6551 -1703 6759 -1693
rect 6794 -1697 6839 -1693
rect 6842 -1694 6843 -1693
rect 6858 -1694 6871 -1693
rect 6577 -1733 6766 -1703
rect 6592 -1736 6766 -1733
rect 6585 -1739 6766 -1736
rect 6394 -1759 6407 -1757
rect 6422 -1759 6456 -1757
rect 6394 -1775 6468 -1759
rect 6495 -1763 6508 -1749
rect 6523 -1763 6539 -1747
rect 6585 -1752 6596 -1739
rect 6378 -1797 6379 -1781
rect 6394 -1797 6407 -1775
rect 6422 -1797 6452 -1775
rect 6495 -1779 6557 -1763
rect 6585 -1770 6596 -1754
rect 6601 -1759 6611 -1739
rect 6621 -1759 6635 -1739
rect 6638 -1752 6647 -1739
rect 6663 -1752 6672 -1739
rect 6601 -1770 6635 -1759
rect 6638 -1770 6647 -1754
rect 6663 -1770 6672 -1754
rect 6679 -1759 6689 -1739
rect 6699 -1759 6713 -1739
rect 6714 -1752 6725 -1739
rect 6679 -1770 6713 -1759
rect 6714 -1770 6725 -1754
rect 6771 -1763 6787 -1747
rect 6794 -1749 6824 -1697
rect 6858 -1701 6859 -1694
rect 6843 -1709 6859 -1701
rect 6830 -1741 6843 -1722
rect 6858 -1741 6888 -1725
rect 6830 -1757 6904 -1741
rect 6830 -1759 6843 -1757
rect 6858 -1759 6892 -1757
rect 6495 -1781 6508 -1779
rect 6523 -1781 6557 -1779
rect 6495 -1797 6557 -1781
rect 6601 -1786 6617 -1783
rect 6679 -1786 6709 -1775
rect 6757 -1779 6803 -1763
rect 6830 -1775 6904 -1759
rect 6757 -1781 6791 -1779
rect 6756 -1797 6803 -1781
rect 6830 -1797 6843 -1775
rect 6858 -1797 6888 -1775
rect 6915 -1797 6916 -1781
rect 6931 -1797 6944 -1637
rect 4595 -1830 4596 -1804
rect 4603 -1830 4630 -1804
rect 4538 -1848 4568 -1834
rect 4595 -1838 4630 -1830
rect 4632 -1805 4673 -1797
rect 4632 -1831 4647 -1805
rect 4654 -1831 4673 -1805
rect 4737 -1809 4799 -1797
rect 4811 -1809 4886 -1797
rect 4944 -1809 5019 -1797
rect 5031 -1809 5062 -1797
rect 5068 -1809 5103 -1797
rect 4737 -1811 4899 -1809
rect 4595 -1848 4596 -1838
rect 4611 -1848 4624 -1838
rect 4632 -1839 4673 -1831
rect 4755 -1835 4768 -1811
rect 4783 -1813 4798 -1811
rect 4832 -1829 4899 -1811
rect 4931 -1811 5103 -1809
rect 4931 -1829 5011 -1811
rect 5032 -1813 5047 -1811
rect 0 -1849 4624 -1848
rect 4638 -1849 4639 -1839
rect 4654 -1849 4667 -1839
rect 4682 -1849 4712 -1835
rect 4755 -1849 4798 -1835
rect 4822 -1838 4829 -1831
rect 4832 -1839 5011 -1829
rect 4805 -1849 4835 -1839
rect 4837 -1849 4990 -1839
rect 4998 -1849 5028 -1839
rect 5032 -1849 5062 -1835
rect 5090 -1849 5103 -1811
rect 5175 -1805 5210 -1797
rect 5175 -1831 5176 -1805
rect 5183 -1831 5210 -1805
rect 5118 -1849 5148 -1835
rect 5175 -1839 5210 -1831
rect 5212 -1805 5253 -1797
rect 5212 -1831 5227 -1805
rect 5234 -1831 5253 -1805
rect 5317 -1809 5379 -1797
rect 5391 -1809 5466 -1797
rect 5524 -1809 5599 -1797
rect 5611 -1809 5642 -1797
rect 5648 -1809 5683 -1797
rect 5317 -1811 5479 -1809
rect 5212 -1839 5253 -1831
rect 5335 -1835 5348 -1811
rect 5363 -1813 5378 -1811
rect 5412 -1829 5479 -1811
rect 5511 -1811 5683 -1809
rect 5511 -1829 5591 -1811
rect 5612 -1813 5627 -1811
rect 5175 -1849 5176 -1839
rect 5191 -1849 5204 -1839
rect 5218 -1849 5219 -1839
rect 5234 -1849 5247 -1839
rect 5262 -1849 5292 -1835
rect 5335 -1849 5378 -1835
rect 5402 -1838 5409 -1831
rect 5412 -1839 5591 -1829
rect 5385 -1849 5415 -1839
rect 5417 -1849 5570 -1839
rect 5578 -1849 5608 -1839
rect 5612 -1849 5642 -1835
rect 5670 -1849 5683 -1811
rect 5755 -1805 5790 -1797
rect 5755 -1831 5756 -1805
rect 5763 -1831 5790 -1805
rect 5698 -1849 5728 -1835
rect 5755 -1839 5790 -1831
rect 5792 -1805 5833 -1797
rect 5792 -1831 5807 -1805
rect 5814 -1831 5833 -1805
rect 5897 -1809 5959 -1797
rect 5971 -1809 6046 -1797
rect 6104 -1809 6179 -1797
rect 6191 -1809 6222 -1797
rect 6228 -1809 6263 -1797
rect 5897 -1811 6059 -1809
rect 5792 -1839 5833 -1831
rect 5915 -1835 5928 -1811
rect 5943 -1813 5958 -1811
rect 5992 -1829 6059 -1811
rect 6091 -1811 6263 -1809
rect 6091 -1829 6171 -1811
rect 6192 -1813 6207 -1811
rect 5755 -1849 5756 -1839
rect 5771 -1849 5784 -1839
rect 5798 -1849 5799 -1839
rect 5814 -1849 5827 -1839
rect 5842 -1849 5872 -1835
rect 5915 -1849 5958 -1835
rect 5982 -1838 5989 -1831
rect 5992 -1839 6171 -1829
rect 5965 -1849 5995 -1839
rect 5997 -1849 6150 -1839
rect 6158 -1849 6188 -1839
rect 6192 -1849 6222 -1835
rect 6250 -1849 6263 -1811
rect 6335 -1805 6370 -1797
rect 6335 -1831 6336 -1805
rect 6343 -1831 6370 -1805
rect 6278 -1849 6308 -1835
rect 6335 -1839 6370 -1831
rect 6372 -1805 6413 -1797
rect 6372 -1831 6387 -1805
rect 6394 -1831 6413 -1805
rect 6477 -1809 6539 -1797
rect 6551 -1809 6626 -1797
rect 6684 -1809 6759 -1797
rect 6771 -1809 6802 -1797
rect 6808 -1809 6843 -1797
rect 6477 -1811 6639 -1809
rect 6372 -1839 6413 -1831
rect 6495 -1835 6508 -1811
rect 6523 -1813 6538 -1811
rect 6572 -1829 6639 -1811
rect 6671 -1811 6843 -1809
rect 6671 -1829 6751 -1811
rect 6772 -1813 6787 -1811
rect 6335 -1849 6336 -1839
rect 6351 -1849 6364 -1839
rect 6378 -1849 6379 -1839
rect 6394 -1849 6407 -1839
rect 6422 -1849 6452 -1835
rect 6495 -1849 6538 -1835
rect 6562 -1838 6569 -1831
rect 6572 -1839 6751 -1829
rect 6545 -1849 6575 -1839
rect 6577 -1849 6730 -1839
rect 6738 -1849 6768 -1839
rect 6772 -1849 6802 -1835
rect 6830 -1849 6843 -1811
rect 6915 -1805 6950 -1797
rect 6915 -1831 6916 -1805
rect 6923 -1831 6950 -1805
rect 6858 -1849 6888 -1835
rect 6915 -1839 6950 -1831
rect 6915 -1849 6916 -1839
rect 6931 -1849 6944 -1839
rect 0 -1862 6944 -1849
rect 14 -1892 27 -1862
rect 42 -1880 72 -1862
rect 115 -1876 129 -1862
rect 165 -1876 385 -1862
rect 116 -1878 129 -1876
rect 82 -1890 97 -1878
rect 79 -1892 101 -1890
rect 106 -1892 136 -1878
rect 197 -1880 350 -1876
rect 179 -1892 371 -1880
rect 414 -1892 444 -1878
rect 450 -1892 463 -1862
rect 478 -1880 508 -1862
rect 551 -1892 564 -1862
rect 594 -1892 607 -1862
rect 622 -1880 652 -1862
rect 695 -1876 709 -1862
rect 745 -1876 965 -1862
rect 696 -1878 709 -1876
rect 662 -1890 677 -1878
rect 659 -1892 681 -1890
rect 686 -1892 716 -1878
rect 777 -1880 930 -1876
rect 759 -1892 951 -1880
rect 994 -1892 1024 -1878
rect 1030 -1892 1043 -1862
rect 1058 -1880 1088 -1862
rect 1131 -1892 1144 -1862
rect 1174 -1892 1187 -1862
rect 1202 -1880 1232 -1862
rect 1275 -1876 1289 -1862
rect 1325 -1876 1545 -1862
rect 1276 -1878 1289 -1876
rect 1242 -1890 1257 -1878
rect 1239 -1892 1261 -1890
rect 1266 -1892 1296 -1878
rect 1357 -1880 1510 -1876
rect 1339 -1892 1531 -1880
rect 1574 -1892 1604 -1878
rect 1610 -1892 1623 -1862
rect 1638 -1880 1668 -1862
rect 1711 -1892 1724 -1862
rect 1754 -1892 1767 -1862
rect 1782 -1880 1812 -1862
rect 1855 -1876 1869 -1862
rect 1905 -1876 2125 -1862
rect 1856 -1878 1869 -1876
rect 1822 -1890 1837 -1878
rect 1819 -1892 1841 -1890
rect 1846 -1892 1876 -1878
rect 1937 -1880 2090 -1876
rect 1919 -1892 2111 -1880
rect 2154 -1892 2184 -1878
rect 2190 -1892 2203 -1862
rect 2218 -1880 2248 -1862
rect 2291 -1892 2304 -1862
rect 2334 -1892 2347 -1862
rect 2362 -1880 2392 -1862
rect 2435 -1876 2449 -1862
rect 2485 -1876 2705 -1862
rect 2436 -1878 2449 -1876
rect 2402 -1890 2417 -1878
rect 2399 -1892 2421 -1890
rect 2426 -1892 2456 -1878
rect 2517 -1880 2670 -1876
rect 2499 -1892 2691 -1880
rect 2734 -1892 2764 -1878
rect 2770 -1892 2783 -1862
rect 2798 -1880 2828 -1862
rect 2871 -1892 2884 -1862
rect 2914 -1892 2927 -1862
rect 2942 -1880 2972 -1862
rect 3015 -1876 3029 -1862
rect 3065 -1876 3285 -1862
rect 3016 -1878 3029 -1876
rect 2982 -1890 2997 -1878
rect 2979 -1892 3001 -1890
rect 3006 -1892 3036 -1878
rect 3097 -1880 3250 -1876
rect 3079 -1892 3271 -1880
rect 3314 -1892 3344 -1878
rect 3350 -1892 3363 -1862
rect 3378 -1880 3408 -1862
rect 3451 -1892 3464 -1862
rect 3494 -1892 3507 -1862
rect 3522 -1880 3552 -1862
rect 3595 -1876 3609 -1862
rect 3645 -1876 3865 -1862
rect 3596 -1878 3609 -1876
rect 3562 -1890 3577 -1878
rect 3559 -1892 3581 -1890
rect 3586 -1892 3616 -1878
rect 3677 -1880 3830 -1876
rect 3659 -1892 3851 -1880
rect 3894 -1892 3924 -1878
rect 3930 -1892 3943 -1862
rect 3958 -1880 3988 -1862
rect 4031 -1892 4044 -1862
rect 4074 -1892 4087 -1862
rect 4102 -1880 4132 -1862
rect 4175 -1876 4189 -1862
rect 4225 -1876 4445 -1862
rect 4176 -1878 4189 -1876
rect 4142 -1890 4157 -1878
rect 4139 -1892 4161 -1890
rect 4166 -1892 4196 -1878
rect 4257 -1880 4410 -1876
rect 4239 -1892 4431 -1880
rect 4474 -1892 4504 -1878
rect 4510 -1892 4523 -1862
rect 4538 -1880 4568 -1862
rect 4611 -1863 6944 -1862
rect 4611 -1892 4624 -1863
rect 0 -1893 4624 -1892
rect 4654 -1893 4667 -1863
rect 4682 -1881 4712 -1863
rect 4755 -1877 4769 -1863
rect 4805 -1877 5025 -1863
rect 4756 -1879 4769 -1877
rect 4722 -1891 4737 -1879
rect 4719 -1893 4741 -1891
rect 4746 -1893 4776 -1879
rect 4837 -1881 4990 -1877
rect 4819 -1893 5011 -1881
rect 5054 -1893 5084 -1879
rect 5090 -1893 5103 -1863
rect 5118 -1881 5148 -1863
rect 5191 -1893 5204 -1863
rect 5234 -1893 5247 -1863
rect 5262 -1881 5292 -1863
rect 5335 -1877 5349 -1863
rect 5385 -1877 5605 -1863
rect 5336 -1879 5349 -1877
rect 5302 -1891 5317 -1879
rect 5299 -1893 5321 -1891
rect 5326 -1893 5356 -1879
rect 5417 -1881 5570 -1877
rect 5399 -1893 5591 -1881
rect 5634 -1893 5664 -1879
rect 5670 -1893 5683 -1863
rect 5698 -1881 5728 -1863
rect 5771 -1893 5784 -1863
rect 5814 -1893 5827 -1863
rect 5842 -1881 5872 -1863
rect 5915 -1877 5929 -1863
rect 5965 -1877 6185 -1863
rect 5916 -1879 5929 -1877
rect 5882 -1891 5897 -1879
rect 5879 -1893 5901 -1891
rect 5906 -1893 5936 -1879
rect 5997 -1881 6150 -1877
rect 5979 -1893 6171 -1881
rect 6214 -1893 6244 -1879
rect 6250 -1893 6263 -1863
rect 6278 -1881 6308 -1863
rect 6351 -1893 6364 -1863
rect 6394 -1893 6407 -1863
rect 6422 -1881 6452 -1863
rect 6495 -1877 6509 -1863
rect 6545 -1877 6765 -1863
rect 6496 -1879 6509 -1877
rect 6462 -1891 6477 -1879
rect 6459 -1893 6481 -1891
rect 6486 -1893 6516 -1879
rect 6577 -1881 6730 -1877
rect 6559 -1893 6751 -1881
rect 6794 -1893 6824 -1879
rect 6830 -1893 6843 -1863
rect 6858 -1881 6888 -1863
rect 6931 -1893 6944 -1863
rect 0 -1906 6944 -1893
rect 14 -2010 27 -1906
rect 72 -1928 73 -1918
rect 88 -1928 101 -1918
rect 72 -1932 101 -1928
rect 106 -1932 136 -1906
rect 154 -1920 170 -1918
rect 242 -1920 295 -1906
rect 243 -1922 307 -1920
rect 154 -1932 169 -1928
rect 72 -1934 169 -1932
rect 56 -1942 107 -1934
rect 56 -1954 81 -1942
rect 88 -1954 107 -1942
rect 138 -1942 188 -1934
rect 138 -1950 154 -1942
rect 161 -1944 188 -1942
rect 197 -1942 212 -1938
rect 259 -1942 291 -1922
rect 350 -1934 365 -1906
rect 414 -1909 444 -1906
rect 414 -1912 450 -1909
rect 380 -1920 396 -1918
rect 381 -1932 396 -1928
rect 414 -1931 453 -1912
rect 472 -1918 479 -1917
rect 478 -1925 479 -1918
rect 462 -1928 463 -1925
rect 478 -1928 491 -1925
rect 414 -1932 444 -1931
rect 453 -1932 459 -1931
rect 462 -1932 491 -1928
rect 381 -1933 491 -1932
rect 381 -1934 497 -1933
rect 350 -1942 418 -1934
rect 197 -1944 266 -1942
rect 284 -1944 418 -1942
rect 161 -1948 233 -1944
rect 161 -1950 286 -1948
rect 161 -1954 233 -1950
rect 56 -1962 107 -1954
rect 154 -1958 233 -1954
rect 314 -1958 418 -1944
rect 447 -1942 497 -1934
rect 447 -1951 463 -1942
rect 154 -1962 418 -1958
rect 444 -1954 463 -1951
rect 470 -1954 497 -1942
rect 444 -1962 497 -1954
rect 72 -1970 73 -1962
rect 88 -1970 101 -1962
rect 72 -1978 88 -1970
rect 69 -1985 88 -1982
rect 69 -1994 91 -1985
rect 42 -2004 91 -1994
rect 42 -2010 72 -2004
rect 91 -2009 96 -2004
rect 14 -2026 88 -2010
rect 106 -2018 136 -1962
rect 171 -1972 379 -1962
rect 414 -1966 459 -1962
rect 462 -1963 463 -1962
rect 478 -1963 491 -1962
rect 338 -1976 386 -1972
rect 221 -1998 251 -1989
rect 314 -1996 329 -1989
rect 350 -1998 386 -1976
rect 197 -2002 386 -1998
rect 212 -2005 386 -2002
rect 205 -2008 386 -2005
rect 14 -2028 27 -2026
rect 42 -2028 76 -2026
rect 14 -2044 88 -2028
rect 115 -2032 128 -2018
rect 143 -2032 159 -2016
rect 205 -2021 216 -2008
rect 14 -2066 27 -2044
rect 42 -2066 72 -2044
rect 115 -2048 177 -2032
rect 205 -2039 216 -2023
rect 221 -2028 231 -2008
rect 241 -2028 255 -2008
rect 258 -2021 267 -2008
rect 283 -2021 292 -2008
rect 221 -2039 255 -2028
rect 258 -2039 266 -2023
rect 283 -2039 292 -2023
rect 299 -2028 309 -2008
rect 319 -2028 333 -2008
rect 334 -2021 345 -2008
rect 299 -2039 333 -2028
rect 334 -2039 345 -2023
rect 391 -2032 407 -2016
rect 414 -2018 444 -1966
rect 478 -1970 479 -1963
rect 463 -1978 479 -1970
rect 450 -2010 463 -1991
rect 478 -2010 508 -1994
rect 450 -2026 524 -2010
rect 450 -2028 463 -2026
rect 478 -2028 512 -2026
rect 115 -2050 128 -2048
rect 143 -2050 177 -2048
rect 115 -2066 177 -2050
rect 221 -2055 234 -2052
rect 299 -2055 329 -2044
rect 377 -2048 423 -2032
rect 450 -2044 524 -2028
rect 377 -2050 411 -2048
rect 376 -2066 423 -2050
rect 450 -2066 463 -2044
rect 478 -2066 508 -2044
rect 535 -2066 536 -2050
rect 551 -2066 564 -1906
rect 594 -2010 607 -1906
rect 652 -1928 653 -1918
rect 668 -1928 681 -1918
rect 652 -1932 681 -1928
rect 686 -1932 716 -1906
rect 734 -1920 750 -1918
rect 822 -1920 875 -1906
rect 823 -1922 887 -1920
rect 734 -1932 749 -1928
rect 652 -1934 749 -1932
rect 636 -1942 687 -1934
rect 636 -1954 661 -1942
rect 668 -1954 687 -1942
rect 718 -1942 768 -1934
rect 718 -1950 734 -1942
rect 741 -1944 768 -1942
rect 777 -1942 792 -1938
rect 839 -1942 871 -1922
rect 930 -1934 945 -1906
rect 994 -1909 1024 -1906
rect 994 -1912 1030 -1909
rect 960 -1920 976 -1918
rect 961 -1932 976 -1928
rect 994 -1931 1033 -1912
rect 1052 -1918 1059 -1917
rect 1058 -1925 1059 -1918
rect 1042 -1928 1043 -1925
rect 1058 -1928 1071 -1925
rect 994 -1932 1024 -1931
rect 1033 -1932 1039 -1931
rect 1042 -1932 1071 -1928
rect 961 -1933 1071 -1932
rect 961 -1934 1077 -1933
rect 930 -1942 998 -1934
rect 777 -1944 846 -1942
rect 864 -1944 998 -1942
rect 741 -1948 813 -1944
rect 741 -1950 866 -1948
rect 741 -1954 813 -1950
rect 636 -1962 687 -1954
rect 734 -1958 813 -1954
rect 894 -1958 998 -1944
rect 1027 -1942 1077 -1934
rect 1027 -1951 1043 -1942
rect 734 -1962 998 -1958
rect 1024 -1954 1043 -1951
rect 1050 -1954 1077 -1942
rect 1024 -1962 1077 -1954
rect 652 -1970 653 -1962
rect 668 -1970 681 -1962
rect 652 -1978 668 -1970
rect 649 -1985 668 -1982
rect 649 -1994 671 -1985
rect 622 -2004 671 -1994
rect 622 -2010 652 -2004
rect 671 -2009 676 -2004
rect 594 -2026 668 -2010
rect 686 -2018 716 -1962
rect 751 -1972 959 -1962
rect 994 -1966 1039 -1962
rect 1042 -1963 1043 -1962
rect 1058 -1963 1071 -1962
rect 918 -1976 966 -1972
rect 801 -1998 831 -1989
rect 894 -1996 909 -1989
rect 930 -1998 966 -1976
rect 777 -2002 966 -1998
rect 792 -2005 966 -2002
rect 785 -2008 966 -2005
rect 594 -2028 607 -2026
rect 622 -2028 656 -2026
rect 594 -2044 668 -2028
rect 695 -2032 708 -2018
rect 723 -2032 739 -2016
rect 785 -2021 796 -2008
rect 578 -2066 579 -2050
rect 594 -2066 607 -2044
rect 622 -2066 652 -2044
rect 695 -2048 757 -2032
rect 785 -2039 796 -2023
rect 801 -2028 811 -2008
rect 821 -2028 835 -2008
rect 838 -2021 847 -2008
rect 863 -2021 872 -2008
rect 801 -2039 835 -2028
rect 838 -2039 846 -2023
rect 863 -2039 872 -2023
rect 879 -2028 889 -2008
rect 899 -2028 913 -2008
rect 914 -2021 925 -2008
rect 879 -2039 913 -2028
rect 914 -2039 925 -2023
rect 971 -2032 987 -2016
rect 994 -2018 1024 -1966
rect 1058 -1970 1059 -1963
rect 1043 -1978 1059 -1970
rect 1030 -2010 1043 -1991
rect 1058 -2010 1088 -1994
rect 1030 -2026 1104 -2010
rect 1030 -2028 1043 -2026
rect 1058 -2028 1092 -2026
rect 695 -2050 708 -2048
rect 723 -2050 757 -2048
rect 695 -2066 757 -2050
rect 801 -2055 814 -2052
rect 879 -2055 909 -2044
rect 957 -2048 1003 -2032
rect 1030 -2044 1104 -2028
rect 957 -2050 991 -2048
rect 956 -2066 1003 -2050
rect 1030 -2066 1043 -2044
rect 1058 -2066 1088 -2044
rect 1115 -2066 1116 -2050
rect 1131 -2066 1144 -1906
rect 1174 -2010 1187 -1906
rect 1232 -1928 1233 -1918
rect 1248 -1928 1261 -1918
rect 1232 -1932 1261 -1928
rect 1266 -1932 1296 -1906
rect 1314 -1920 1330 -1918
rect 1402 -1920 1455 -1906
rect 1403 -1922 1467 -1920
rect 1314 -1932 1329 -1928
rect 1232 -1934 1329 -1932
rect 1216 -1942 1267 -1934
rect 1216 -1954 1241 -1942
rect 1248 -1954 1267 -1942
rect 1298 -1942 1348 -1934
rect 1298 -1950 1314 -1942
rect 1321 -1944 1348 -1942
rect 1357 -1942 1372 -1938
rect 1419 -1942 1451 -1922
rect 1510 -1934 1525 -1906
rect 1574 -1909 1604 -1906
rect 1574 -1912 1610 -1909
rect 1540 -1920 1556 -1918
rect 1541 -1932 1556 -1928
rect 1574 -1931 1613 -1912
rect 1632 -1918 1639 -1917
rect 1638 -1925 1639 -1918
rect 1622 -1928 1623 -1925
rect 1638 -1928 1651 -1925
rect 1574 -1932 1604 -1931
rect 1613 -1932 1619 -1931
rect 1622 -1932 1651 -1928
rect 1541 -1933 1651 -1932
rect 1541 -1934 1657 -1933
rect 1510 -1942 1578 -1934
rect 1357 -1944 1426 -1942
rect 1444 -1944 1578 -1942
rect 1321 -1948 1393 -1944
rect 1321 -1950 1446 -1948
rect 1321 -1954 1393 -1950
rect 1216 -1962 1267 -1954
rect 1314 -1958 1393 -1954
rect 1474 -1958 1578 -1944
rect 1607 -1942 1657 -1934
rect 1607 -1951 1623 -1942
rect 1314 -1962 1578 -1958
rect 1604 -1954 1623 -1951
rect 1630 -1954 1657 -1942
rect 1604 -1962 1657 -1954
rect 1232 -1970 1233 -1962
rect 1248 -1970 1261 -1962
rect 1232 -1978 1248 -1970
rect 1229 -1985 1248 -1982
rect 1229 -1994 1251 -1985
rect 1202 -2004 1251 -1994
rect 1202 -2010 1232 -2004
rect 1251 -2009 1256 -2004
rect 1174 -2026 1248 -2010
rect 1266 -2018 1296 -1962
rect 1331 -1972 1539 -1962
rect 1574 -1966 1619 -1962
rect 1622 -1963 1623 -1962
rect 1638 -1963 1651 -1962
rect 1498 -1976 1546 -1972
rect 1381 -1998 1411 -1989
rect 1474 -1996 1489 -1989
rect 1510 -1998 1546 -1976
rect 1357 -2002 1546 -1998
rect 1372 -2005 1546 -2002
rect 1365 -2008 1546 -2005
rect 1174 -2028 1187 -2026
rect 1202 -2028 1236 -2026
rect 1174 -2044 1248 -2028
rect 1275 -2032 1288 -2018
rect 1303 -2032 1319 -2016
rect 1365 -2021 1376 -2008
rect 1158 -2066 1159 -2050
rect 1174 -2066 1187 -2044
rect 1202 -2066 1232 -2044
rect 1275 -2048 1337 -2032
rect 1365 -2039 1376 -2023
rect 1381 -2028 1391 -2008
rect 1401 -2028 1415 -2008
rect 1418 -2021 1427 -2008
rect 1443 -2021 1452 -2008
rect 1381 -2039 1415 -2028
rect 1418 -2039 1426 -2023
rect 1443 -2039 1452 -2023
rect 1459 -2028 1469 -2008
rect 1479 -2028 1493 -2008
rect 1494 -2021 1505 -2008
rect 1459 -2039 1493 -2028
rect 1494 -2039 1505 -2023
rect 1551 -2032 1567 -2016
rect 1574 -2018 1604 -1966
rect 1638 -1970 1639 -1963
rect 1623 -1978 1639 -1970
rect 1610 -2010 1623 -1991
rect 1638 -2010 1668 -1994
rect 1610 -2026 1684 -2010
rect 1610 -2028 1623 -2026
rect 1638 -2028 1672 -2026
rect 1275 -2050 1288 -2048
rect 1303 -2050 1337 -2048
rect 1275 -2066 1337 -2050
rect 1381 -2055 1394 -2052
rect 1459 -2055 1489 -2044
rect 1537 -2048 1583 -2032
rect 1610 -2044 1684 -2028
rect 1537 -2050 1571 -2048
rect 1536 -2066 1583 -2050
rect 1610 -2066 1623 -2044
rect 1638 -2066 1668 -2044
rect 1695 -2066 1696 -2050
rect 1711 -2066 1724 -1906
rect 1754 -2010 1767 -1906
rect 1812 -1928 1813 -1918
rect 1828 -1928 1841 -1918
rect 1812 -1932 1841 -1928
rect 1846 -1932 1876 -1906
rect 1894 -1920 1910 -1918
rect 1982 -1920 2035 -1906
rect 1983 -1922 2047 -1920
rect 1894 -1932 1909 -1928
rect 1812 -1934 1909 -1932
rect 1796 -1942 1847 -1934
rect 1796 -1954 1821 -1942
rect 1828 -1954 1847 -1942
rect 1878 -1942 1928 -1934
rect 1878 -1950 1894 -1942
rect 1901 -1944 1928 -1942
rect 1937 -1942 1952 -1938
rect 1999 -1942 2031 -1922
rect 2090 -1934 2105 -1906
rect 2154 -1909 2184 -1906
rect 2154 -1912 2190 -1909
rect 2120 -1920 2136 -1918
rect 2121 -1932 2136 -1928
rect 2154 -1931 2193 -1912
rect 2212 -1918 2219 -1917
rect 2218 -1925 2219 -1918
rect 2202 -1928 2203 -1925
rect 2218 -1928 2231 -1925
rect 2154 -1932 2184 -1931
rect 2193 -1932 2199 -1931
rect 2202 -1932 2231 -1928
rect 2121 -1933 2231 -1932
rect 2121 -1934 2237 -1933
rect 2090 -1942 2158 -1934
rect 1937 -1944 2006 -1942
rect 2024 -1944 2158 -1942
rect 1901 -1948 1973 -1944
rect 1901 -1950 2026 -1948
rect 1901 -1954 1973 -1950
rect 1796 -1962 1847 -1954
rect 1894 -1958 1973 -1954
rect 2054 -1958 2158 -1944
rect 2187 -1942 2237 -1934
rect 2187 -1951 2203 -1942
rect 1894 -1962 2158 -1958
rect 2184 -1954 2203 -1951
rect 2210 -1954 2237 -1942
rect 2184 -1962 2237 -1954
rect 1812 -1970 1813 -1962
rect 1828 -1970 1841 -1962
rect 1812 -1978 1828 -1970
rect 1809 -1985 1828 -1982
rect 1809 -1994 1831 -1985
rect 1782 -2004 1831 -1994
rect 1782 -2010 1812 -2004
rect 1831 -2009 1836 -2004
rect 1754 -2026 1828 -2010
rect 1846 -2018 1876 -1962
rect 1911 -1972 2119 -1962
rect 2154 -1966 2199 -1962
rect 2202 -1963 2203 -1962
rect 2218 -1963 2231 -1962
rect 2078 -1976 2126 -1972
rect 1961 -1998 1991 -1989
rect 2054 -1996 2069 -1989
rect 2090 -1998 2126 -1976
rect 1937 -2002 2126 -1998
rect 1952 -2005 2126 -2002
rect 1945 -2008 2126 -2005
rect 1754 -2028 1767 -2026
rect 1782 -2028 1816 -2026
rect 1754 -2044 1828 -2028
rect 1855 -2032 1868 -2018
rect 1883 -2032 1899 -2016
rect 1945 -2021 1956 -2008
rect 1738 -2066 1739 -2050
rect 1754 -2066 1767 -2044
rect 1782 -2066 1812 -2044
rect 1855 -2048 1917 -2032
rect 1945 -2039 1956 -2023
rect 1961 -2028 1971 -2008
rect 1981 -2028 1995 -2008
rect 1998 -2021 2007 -2008
rect 2023 -2021 2032 -2008
rect 1961 -2039 1995 -2028
rect 1998 -2039 2006 -2023
rect 2023 -2039 2032 -2023
rect 2039 -2028 2049 -2008
rect 2059 -2028 2073 -2008
rect 2074 -2021 2085 -2008
rect 2039 -2039 2073 -2028
rect 2074 -2039 2085 -2023
rect 2131 -2032 2147 -2016
rect 2154 -2018 2184 -1966
rect 2218 -1970 2219 -1963
rect 2203 -1978 2219 -1970
rect 2190 -2010 2203 -1991
rect 2218 -2010 2248 -1994
rect 2190 -2026 2264 -2010
rect 2190 -2028 2203 -2026
rect 2218 -2028 2252 -2026
rect 1855 -2050 1868 -2048
rect 1883 -2050 1917 -2048
rect 1855 -2066 1917 -2050
rect 1961 -2055 1974 -2052
rect 2039 -2055 2069 -2044
rect 2117 -2048 2163 -2032
rect 2190 -2044 2264 -2028
rect 2117 -2050 2151 -2048
rect 2116 -2066 2163 -2050
rect 2190 -2066 2203 -2044
rect 2218 -2066 2248 -2044
rect 2275 -2066 2276 -2050
rect 2291 -2066 2304 -1906
rect 2334 -2010 2347 -1906
rect 2392 -1928 2393 -1918
rect 2408 -1928 2421 -1918
rect 2392 -1932 2421 -1928
rect 2426 -1932 2456 -1906
rect 2474 -1920 2490 -1918
rect 2562 -1920 2615 -1906
rect 2563 -1922 2627 -1920
rect 2474 -1932 2489 -1928
rect 2392 -1934 2489 -1932
rect 2376 -1942 2427 -1934
rect 2376 -1954 2401 -1942
rect 2408 -1954 2427 -1942
rect 2458 -1942 2508 -1934
rect 2458 -1950 2474 -1942
rect 2481 -1944 2508 -1942
rect 2517 -1942 2532 -1938
rect 2579 -1942 2611 -1922
rect 2670 -1934 2685 -1906
rect 2734 -1909 2764 -1906
rect 2734 -1912 2770 -1909
rect 2700 -1920 2716 -1918
rect 2701 -1932 2716 -1928
rect 2734 -1931 2773 -1912
rect 2792 -1918 2799 -1917
rect 2798 -1925 2799 -1918
rect 2782 -1928 2783 -1925
rect 2798 -1928 2811 -1925
rect 2734 -1932 2764 -1931
rect 2773 -1932 2779 -1931
rect 2782 -1932 2811 -1928
rect 2701 -1933 2811 -1932
rect 2701 -1934 2817 -1933
rect 2670 -1942 2738 -1934
rect 2517 -1944 2586 -1942
rect 2604 -1944 2738 -1942
rect 2481 -1948 2553 -1944
rect 2481 -1950 2606 -1948
rect 2481 -1954 2553 -1950
rect 2376 -1962 2427 -1954
rect 2474 -1958 2553 -1954
rect 2634 -1958 2738 -1944
rect 2767 -1942 2817 -1934
rect 2767 -1951 2783 -1942
rect 2474 -1962 2738 -1958
rect 2764 -1954 2783 -1951
rect 2790 -1954 2817 -1942
rect 2764 -1962 2817 -1954
rect 2392 -1970 2393 -1962
rect 2408 -1970 2421 -1962
rect 2392 -1978 2408 -1970
rect 2389 -1985 2408 -1982
rect 2389 -1994 2411 -1985
rect 2362 -2004 2411 -1994
rect 2362 -2010 2392 -2004
rect 2411 -2009 2416 -2004
rect 2334 -2026 2408 -2010
rect 2426 -2018 2456 -1962
rect 2491 -1972 2699 -1962
rect 2734 -1966 2779 -1962
rect 2782 -1963 2783 -1962
rect 2798 -1963 2811 -1962
rect 2658 -1976 2706 -1972
rect 2541 -1998 2571 -1989
rect 2634 -1996 2649 -1989
rect 2670 -1998 2706 -1976
rect 2517 -2002 2706 -1998
rect 2532 -2005 2706 -2002
rect 2525 -2008 2706 -2005
rect 2334 -2028 2347 -2026
rect 2362 -2028 2396 -2026
rect 2334 -2044 2408 -2028
rect 2435 -2032 2448 -2018
rect 2463 -2032 2479 -2016
rect 2525 -2021 2536 -2008
rect 2318 -2066 2319 -2050
rect 2334 -2066 2347 -2044
rect 2362 -2066 2392 -2044
rect 2435 -2048 2497 -2032
rect 2525 -2039 2536 -2023
rect 2541 -2028 2551 -2008
rect 2561 -2028 2575 -2008
rect 2578 -2021 2587 -2008
rect 2603 -2021 2612 -2008
rect 2541 -2039 2575 -2028
rect 2578 -2039 2586 -2023
rect 2603 -2039 2612 -2023
rect 2619 -2028 2629 -2008
rect 2639 -2028 2653 -2008
rect 2654 -2021 2665 -2008
rect 2619 -2039 2653 -2028
rect 2654 -2039 2665 -2023
rect 2711 -2032 2727 -2016
rect 2734 -2018 2764 -1966
rect 2798 -1970 2799 -1963
rect 2783 -1978 2799 -1970
rect 2770 -2010 2783 -1991
rect 2798 -2010 2828 -1994
rect 2770 -2026 2844 -2010
rect 2770 -2028 2783 -2026
rect 2798 -2028 2832 -2026
rect 2435 -2050 2448 -2048
rect 2463 -2050 2497 -2048
rect 2435 -2066 2497 -2050
rect 2541 -2055 2554 -2052
rect 2619 -2055 2649 -2044
rect 2697 -2048 2743 -2032
rect 2770 -2044 2844 -2028
rect 2697 -2050 2731 -2048
rect 2696 -2066 2743 -2050
rect 2770 -2066 2783 -2044
rect 2798 -2066 2828 -2044
rect 2855 -2066 2856 -2050
rect 2871 -2066 2884 -1906
rect 2914 -2010 2927 -1906
rect 2972 -1928 2973 -1918
rect 2988 -1928 3001 -1918
rect 2972 -1932 3001 -1928
rect 3006 -1932 3036 -1906
rect 3054 -1920 3070 -1918
rect 3142 -1920 3195 -1906
rect 3143 -1922 3205 -1920
rect 3054 -1932 3069 -1928
rect 2972 -1934 3069 -1932
rect 2956 -1942 3007 -1934
rect 2956 -1954 2981 -1942
rect 2988 -1954 3007 -1942
rect 3038 -1942 3088 -1934
rect 3038 -1950 3054 -1942
rect 3061 -1944 3088 -1942
rect 3097 -1942 3112 -1938
rect 3159 -1942 3191 -1922
rect 3250 -1934 3265 -1906
rect 3314 -1909 3344 -1906
rect 3314 -1912 3350 -1909
rect 3280 -1920 3296 -1918
rect 3281 -1932 3296 -1928
rect 3314 -1931 3353 -1912
rect 3372 -1918 3379 -1917
rect 3378 -1925 3379 -1918
rect 3362 -1928 3363 -1925
rect 3378 -1928 3391 -1925
rect 3314 -1932 3344 -1931
rect 3353 -1932 3359 -1931
rect 3362 -1932 3391 -1928
rect 3281 -1933 3391 -1932
rect 3281 -1934 3397 -1933
rect 3250 -1942 3318 -1934
rect 3097 -1944 3166 -1942
rect 3184 -1944 3318 -1942
rect 3061 -1948 3133 -1944
rect 3061 -1950 3186 -1948
rect 3061 -1954 3133 -1950
rect 2956 -1962 3007 -1954
rect 3054 -1958 3133 -1954
rect 3214 -1958 3318 -1944
rect 3347 -1942 3397 -1934
rect 3347 -1951 3363 -1942
rect 3054 -1962 3318 -1958
rect 3344 -1954 3363 -1951
rect 3370 -1954 3397 -1942
rect 3344 -1962 3397 -1954
rect 2972 -1970 2973 -1962
rect 2988 -1970 3001 -1962
rect 2972 -1978 2988 -1970
rect 2969 -1985 2988 -1982
rect 2969 -1994 2991 -1985
rect 2942 -2004 2991 -1994
rect 2942 -2010 2972 -2004
rect 2991 -2009 2996 -2004
rect 2914 -2026 2988 -2010
rect 3006 -2018 3036 -1962
rect 3071 -1972 3279 -1962
rect 3314 -1966 3359 -1962
rect 3362 -1963 3363 -1962
rect 3378 -1963 3391 -1962
rect 3238 -1976 3286 -1972
rect 3121 -1998 3151 -1989
rect 3214 -1996 3229 -1989
rect 3250 -1998 3286 -1976
rect 3097 -2002 3286 -1998
rect 3112 -2005 3286 -2002
rect 3105 -2008 3286 -2005
rect 2914 -2028 2927 -2026
rect 2942 -2028 2976 -2026
rect 2914 -2044 2988 -2028
rect 3015 -2032 3028 -2018
rect 3043 -2032 3059 -2016
rect 3105 -2021 3116 -2008
rect 2898 -2066 2899 -2050
rect 2914 -2066 2927 -2044
rect 2942 -2066 2972 -2044
rect 3015 -2048 3077 -2032
rect 3105 -2039 3116 -2023
rect 3121 -2028 3131 -2008
rect 3141 -2028 3155 -2008
rect 3158 -2021 3167 -2008
rect 3183 -2021 3192 -2008
rect 3121 -2039 3155 -2028
rect 3158 -2039 3166 -2023
rect 3183 -2039 3192 -2023
rect 3199 -2028 3209 -2008
rect 3219 -2028 3233 -2008
rect 3234 -2021 3245 -2008
rect 3199 -2039 3233 -2028
rect 3234 -2039 3245 -2023
rect 3291 -2032 3307 -2016
rect 3314 -2018 3344 -1966
rect 3378 -1970 3379 -1963
rect 3363 -1978 3379 -1970
rect 3350 -2010 3363 -1991
rect 3378 -2010 3408 -1994
rect 3350 -2026 3424 -2010
rect 3350 -2028 3363 -2026
rect 3378 -2028 3412 -2026
rect 3015 -2050 3028 -2048
rect 3043 -2050 3077 -2048
rect 3015 -2066 3077 -2050
rect 3121 -2055 3134 -2052
rect 3199 -2055 3229 -2044
rect 3277 -2048 3323 -2032
rect 3350 -2044 3424 -2028
rect 3277 -2050 3311 -2048
rect 3276 -2066 3323 -2050
rect 3350 -2066 3363 -2044
rect 3378 -2066 3408 -2044
rect 3435 -2066 3436 -2050
rect 3451 -2066 3464 -1906
rect 3494 -2010 3507 -1906
rect 3552 -1928 3553 -1918
rect 3568 -1928 3581 -1918
rect 3552 -1932 3581 -1928
rect 3586 -1932 3616 -1906
rect 3634 -1920 3650 -1918
rect 3722 -1920 3775 -1906
rect 3723 -1922 3787 -1920
rect 3634 -1932 3649 -1928
rect 3552 -1934 3649 -1932
rect 3536 -1942 3587 -1934
rect 3536 -1954 3561 -1942
rect 3568 -1954 3587 -1942
rect 3618 -1942 3668 -1934
rect 3618 -1950 3634 -1942
rect 3641 -1944 3668 -1942
rect 3677 -1942 3692 -1938
rect 3739 -1942 3771 -1922
rect 3830 -1934 3845 -1906
rect 3894 -1909 3924 -1906
rect 3894 -1912 3930 -1909
rect 3860 -1920 3876 -1918
rect 3861 -1932 3876 -1928
rect 3894 -1931 3933 -1912
rect 3952 -1918 3959 -1917
rect 3958 -1925 3959 -1918
rect 3942 -1928 3943 -1925
rect 3958 -1928 3971 -1925
rect 3894 -1932 3924 -1931
rect 3933 -1932 3939 -1931
rect 3942 -1932 3971 -1928
rect 3861 -1933 3971 -1932
rect 3861 -1934 3977 -1933
rect 3830 -1942 3898 -1934
rect 3677 -1944 3746 -1942
rect 3764 -1944 3898 -1942
rect 3641 -1948 3713 -1944
rect 3641 -1950 3766 -1948
rect 3641 -1954 3713 -1950
rect 3536 -1962 3587 -1954
rect 3634 -1958 3713 -1954
rect 3794 -1958 3898 -1944
rect 3927 -1942 3977 -1934
rect 3927 -1951 3943 -1942
rect 3634 -1962 3898 -1958
rect 3924 -1954 3943 -1951
rect 3950 -1954 3977 -1942
rect 3924 -1962 3977 -1954
rect 3552 -1970 3553 -1962
rect 3568 -1970 3581 -1962
rect 3552 -1978 3568 -1970
rect 3549 -1985 3568 -1982
rect 3549 -1994 3571 -1985
rect 3522 -2004 3571 -1994
rect 3522 -2010 3552 -2004
rect 3571 -2009 3576 -2004
rect 3494 -2026 3568 -2010
rect 3586 -2018 3616 -1962
rect 3651 -1972 3859 -1962
rect 3894 -1966 3939 -1962
rect 3942 -1963 3943 -1962
rect 3958 -1963 3971 -1962
rect 3818 -1976 3866 -1972
rect 3701 -1998 3731 -1989
rect 3794 -1996 3809 -1989
rect 3830 -1998 3866 -1976
rect 3677 -2002 3866 -1998
rect 3692 -2005 3866 -2002
rect 3685 -2008 3866 -2005
rect 3494 -2028 3507 -2026
rect 3522 -2028 3556 -2026
rect 3494 -2044 3568 -2028
rect 3595 -2032 3608 -2018
rect 3623 -2032 3639 -2016
rect 3685 -2021 3696 -2008
rect 3478 -2066 3479 -2050
rect 3494 -2066 3507 -2044
rect 3522 -2066 3552 -2044
rect 3595 -2048 3657 -2032
rect 3685 -2039 3696 -2023
rect 3701 -2028 3711 -2008
rect 3721 -2028 3735 -2008
rect 3738 -2021 3747 -2008
rect 3763 -2021 3772 -2008
rect 3701 -2039 3735 -2028
rect 3738 -2039 3746 -2023
rect 3763 -2039 3772 -2023
rect 3779 -2028 3789 -2008
rect 3799 -2028 3813 -2008
rect 3814 -2021 3825 -2008
rect 3779 -2039 3813 -2028
rect 3814 -2039 3825 -2023
rect 3871 -2032 3887 -2016
rect 3894 -2018 3924 -1966
rect 3958 -1970 3959 -1963
rect 3943 -1978 3959 -1970
rect 3930 -2010 3943 -1991
rect 3958 -2010 3988 -1994
rect 3930 -2026 4004 -2010
rect 3930 -2028 3943 -2026
rect 3958 -2028 3992 -2026
rect 3595 -2050 3608 -2048
rect 3623 -2050 3657 -2048
rect 3595 -2066 3657 -2050
rect 3701 -2055 3714 -2052
rect 3779 -2055 3809 -2044
rect 3857 -2048 3903 -2032
rect 3930 -2044 4004 -2028
rect 3857 -2050 3891 -2048
rect 3856 -2066 3903 -2050
rect 3930 -2066 3943 -2044
rect 3958 -2066 3988 -2044
rect 4015 -2066 4016 -2050
rect 4031 -2066 4044 -1906
rect 4074 -2010 4087 -1906
rect 4132 -1928 4133 -1918
rect 4148 -1928 4161 -1918
rect 4132 -1932 4161 -1928
rect 4166 -1932 4196 -1906
rect 4214 -1920 4230 -1918
rect 4302 -1920 4355 -1906
rect 4303 -1922 4367 -1920
rect 4214 -1932 4229 -1928
rect 4132 -1934 4229 -1932
rect 4116 -1942 4167 -1934
rect 4116 -1954 4141 -1942
rect 4148 -1954 4167 -1942
rect 4198 -1942 4248 -1934
rect 4198 -1950 4214 -1942
rect 4221 -1944 4248 -1942
rect 4257 -1942 4272 -1938
rect 4319 -1942 4351 -1922
rect 4410 -1934 4425 -1906
rect 4474 -1909 4504 -1906
rect 4611 -1907 6944 -1906
rect 4474 -1912 4510 -1909
rect 4440 -1920 4456 -1918
rect 4441 -1932 4456 -1928
rect 4474 -1931 4513 -1912
rect 4532 -1918 4539 -1917
rect 4538 -1925 4539 -1918
rect 4522 -1928 4523 -1925
rect 4538 -1928 4551 -1925
rect 4474 -1932 4504 -1931
rect 4513 -1932 4519 -1931
rect 4522 -1932 4551 -1928
rect 4441 -1933 4551 -1932
rect 4441 -1934 4557 -1933
rect 4410 -1942 4478 -1934
rect 4257 -1944 4326 -1942
rect 4344 -1944 4478 -1942
rect 4221 -1948 4293 -1944
rect 4221 -1950 4346 -1948
rect 4221 -1954 4293 -1950
rect 4116 -1962 4167 -1954
rect 4214 -1958 4293 -1954
rect 4374 -1958 4478 -1944
rect 4507 -1942 4557 -1934
rect 4507 -1951 4523 -1942
rect 4214 -1962 4478 -1958
rect 4504 -1954 4523 -1951
rect 4530 -1954 4557 -1942
rect 4504 -1962 4557 -1954
rect 4132 -1970 4133 -1962
rect 4148 -1970 4161 -1962
rect 4132 -1978 4148 -1970
rect 4129 -1985 4148 -1982
rect 4129 -1994 4151 -1985
rect 4102 -2004 4151 -1994
rect 4102 -2010 4132 -2004
rect 4151 -2009 4156 -2004
rect 4074 -2026 4148 -2010
rect 4166 -2018 4196 -1962
rect 4231 -1972 4439 -1962
rect 4474 -1966 4519 -1962
rect 4522 -1963 4523 -1962
rect 4538 -1963 4551 -1962
rect 4398 -1976 4446 -1972
rect 4281 -1998 4311 -1989
rect 4374 -1996 4389 -1989
rect 4410 -1998 4446 -1976
rect 4257 -2002 4446 -1998
rect 4272 -2005 4446 -2002
rect 4265 -2008 4446 -2005
rect 4074 -2028 4087 -2026
rect 4102 -2028 4136 -2026
rect 4074 -2044 4148 -2028
rect 4175 -2032 4188 -2018
rect 4203 -2032 4219 -2016
rect 4265 -2021 4276 -2008
rect 4058 -2066 4059 -2050
rect 4074 -2066 4087 -2044
rect 4102 -2066 4132 -2044
rect 4175 -2048 4237 -2032
rect 4265 -2039 4276 -2023
rect 4281 -2028 4291 -2008
rect 4301 -2028 4315 -2008
rect 4318 -2021 4327 -2008
rect 4343 -2021 4352 -2008
rect 4281 -2039 4315 -2028
rect 4318 -2039 4326 -2023
rect 4343 -2039 4352 -2023
rect 4359 -2028 4369 -2008
rect 4379 -2028 4393 -2008
rect 4394 -2021 4405 -2008
rect 4359 -2039 4393 -2028
rect 4394 -2039 4405 -2023
rect 4451 -2032 4467 -2016
rect 4474 -2018 4504 -1966
rect 4538 -1970 4539 -1963
rect 4523 -1978 4539 -1970
rect 4510 -2010 4523 -1991
rect 4538 -2010 4568 -1994
rect 4510 -2026 4584 -2010
rect 4510 -2028 4523 -2026
rect 4538 -2028 4572 -2026
rect 4175 -2050 4188 -2048
rect 4203 -2050 4237 -2048
rect 4175 -2066 4237 -2050
rect 4281 -2055 4294 -2052
rect 4359 -2055 4389 -2044
rect 4437 -2048 4483 -2032
rect 4510 -2044 4584 -2028
rect 4437 -2050 4471 -2048
rect 4436 -2066 4483 -2050
rect 4510 -2066 4523 -2044
rect 4538 -2066 4568 -2044
rect 4595 -2066 4596 -2050
rect 4611 -2066 4624 -1907
rect 4654 -2011 4667 -1907
rect 4712 -1929 4713 -1919
rect 4733 -1921 4741 -1919
rect 4731 -1923 4741 -1921
rect 4728 -1929 4741 -1923
rect 4712 -1933 4741 -1929
rect 4746 -1933 4776 -1907
rect 4794 -1921 4810 -1919
rect 4882 -1921 4933 -1907
rect 4883 -1923 4947 -1921
rect 4794 -1933 4809 -1929
rect 4712 -1935 4809 -1933
rect 4696 -1943 4747 -1935
rect 4696 -1955 4721 -1943
rect 4728 -1955 4747 -1943
rect 4778 -1943 4828 -1935
rect 4778 -1951 4794 -1943
rect 4801 -1945 4828 -1943
rect 4837 -1943 4852 -1939
rect 4899 -1943 4931 -1923
rect 4990 -1935 5005 -1907
rect 5054 -1910 5084 -1907
rect 5054 -1913 5090 -1910
rect 5020 -1921 5036 -1919
rect 5021 -1933 5036 -1929
rect 5054 -1932 5093 -1913
rect 5112 -1919 5119 -1918
rect 5118 -1926 5119 -1919
rect 5102 -1929 5103 -1926
rect 5118 -1929 5131 -1926
rect 5054 -1933 5084 -1932
rect 5093 -1933 5099 -1932
rect 5102 -1933 5131 -1929
rect 5021 -1934 5131 -1933
rect 5021 -1935 5137 -1934
rect 4990 -1943 5058 -1935
rect 4837 -1945 4906 -1943
rect 4924 -1945 5058 -1943
rect 4801 -1949 4873 -1945
rect 4801 -1951 4926 -1949
rect 4801 -1955 4873 -1951
rect 4696 -1963 4747 -1955
rect 4794 -1959 4873 -1955
rect 4954 -1959 5058 -1945
rect 5087 -1943 5137 -1935
rect 5087 -1952 5103 -1943
rect 4794 -1963 5058 -1959
rect 5084 -1955 5103 -1952
rect 5110 -1955 5137 -1943
rect 5084 -1963 5137 -1955
rect 4712 -1971 4713 -1963
rect 4728 -1971 4741 -1963
rect 4712 -1979 4728 -1971
rect 4709 -1986 4728 -1983
rect 4709 -1995 4731 -1986
rect 4682 -2005 4731 -1995
rect 4682 -2011 4712 -2005
rect 4731 -2010 4736 -2005
rect 4654 -2027 4728 -2011
rect 4746 -2019 4776 -1963
rect 4811 -1973 5019 -1963
rect 5054 -1967 5099 -1963
rect 5102 -1964 5103 -1963
rect 5118 -1964 5131 -1963
rect 4978 -1977 5026 -1973
rect 4861 -1999 4891 -1990
rect 4954 -1997 4969 -1990
rect 4990 -1999 5026 -1977
rect 4837 -2003 5026 -1999
rect 4852 -2006 5026 -2003
rect 4845 -2009 5026 -2006
rect 4654 -2029 4667 -2027
rect 4682 -2029 4716 -2027
rect 4654 -2045 4728 -2029
rect 4755 -2033 4768 -2019
rect 4783 -2033 4799 -2017
rect 4845 -2022 4856 -2009
rect 0 -2074 33 -2066
rect 0 -2100 7 -2074
rect 14 -2100 33 -2074
rect 97 -2078 159 -2066
rect 171 -2078 246 -2066
rect 304 -2078 379 -2066
rect 391 -2078 422 -2066
rect 428 -2078 463 -2066
rect 97 -2080 259 -2078
rect 0 -2108 33 -2100
rect 115 -2108 128 -2080
rect 143 -2082 158 -2080
rect 182 -2107 189 -2100
rect 192 -2108 259 -2080
rect 291 -2080 463 -2078
rect 261 -2102 289 -2098
rect 291 -2102 371 -2080
rect 392 -2082 407 -2080
rect 261 -2104 371 -2102
rect 261 -2108 289 -2104
rect 291 -2108 371 -2104
rect 14 -2118 27 -2108
rect 42 -2118 72 -2108
rect 115 -2118 158 -2108
rect 165 -2118 173 -2108
rect 192 -2116 195 -2108
rect 259 -2116 291 -2108
rect 192 -2118 358 -2116
rect 377 -2118 388 -2108
rect 392 -2118 422 -2108
rect 450 -2118 463 -2080
rect 535 -2074 570 -2066
rect 535 -2100 536 -2074
rect 543 -2100 570 -2074
rect 535 -2108 570 -2100
rect 572 -2074 613 -2066
rect 572 -2100 587 -2074
rect 594 -2100 613 -2074
rect 677 -2078 739 -2066
rect 751 -2078 826 -2066
rect 884 -2078 959 -2066
rect 971 -2078 1002 -2066
rect 1008 -2078 1043 -2066
rect 677 -2080 839 -2078
rect 572 -2108 613 -2100
rect 695 -2108 708 -2080
rect 723 -2082 738 -2080
rect 762 -2107 769 -2100
rect 772 -2108 839 -2080
rect 871 -2080 1043 -2078
rect 841 -2102 869 -2098
rect 871 -2102 951 -2080
rect 972 -2082 987 -2080
rect 841 -2104 951 -2102
rect 841 -2108 869 -2104
rect 871 -2108 951 -2104
rect 478 -2118 508 -2108
rect 535 -2118 536 -2108
rect 551 -2118 564 -2108
rect 578 -2118 579 -2108
rect 594 -2118 607 -2108
rect 622 -2118 652 -2108
rect 695 -2118 738 -2108
rect 745 -2118 753 -2108
rect 772 -2116 775 -2108
rect 839 -2116 871 -2108
rect 772 -2118 938 -2116
rect 957 -2118 968 -2108
rect 972 -2118 1002 -2108
rect 1030 -2118 1043 -2080
rect 1115 -2074 1150 -2066
rect 1115 -2100 1116 -2074
rect 1123 -2100 1150 -2074
rect 1115 -2108 1150 -2100
rect 1152 -2074 1193 -2066
rect 1152 -2100 1167 -2074
rect 1174 -2100 1193 -2074
rect 1257 -2078 1319 -2066
rect 1331 -2078 1406 -2066
rect 1464 -2078 1539 -2066
rect 1551 -2078 1582 -2066
rect 1588 -2078 1623 -2066
rect 1257 -2080 1419 -2078
rect 1152 -2108 1193 -2100
rect 1275 -2108 1288 -2080
rect 1303 -2082 1318 -2080
rect 1342 -2107 1349 -2100
rect 1352 -2108 1419 -2080
rect 1451 -2080 1623 -2078
rect 1421 -2102 1449 -2098
rect 1451 -2102 1531 -2080
rect 1552 -2082 1567 -2080
rect 1421 -2104 1531 -2102
rect 1421 -2108 1449 -2104
rect 1451 -2108 1531 -2104
rect 1058 -2118 1088 -2108
rect 1115 -2118 1116 -2108
rect 1131 -2118 1144 -2108
rect 1158 -2118 1159 -2108
rect 1174 -2118 1187 -2108
rect 1202 -2118 1232 -2108
rect 1275 -2118 1318 -2108
rect 1325 -2118 1333 -2108
rect 1352 -2116 1355 -2108
rect 1419 -2116 1451 -2108
rect 1352 -2118 1518 -2116
rect 1537 -2118 1548 -2108
rect 1552 -2118 1582 -2108
rect 1610 -2118 1623 -2080
rect 1695 -2074 1730 -2066
rect 1695 -2100 1696 -2074
rect 1703 -2100 1730 -2074
rect 1695 -2108 1730 -2100
rect 1732 -2074 1773 -2066
rect 1732 -2100 1747 -2074
rect 1754 -2100 1773 -2074
rect 1837 -2078 1899 -2066
rect 1911 -2078 1986 -2066
rect 2044 -2078 2119 -2066
rect 2131 -2078 2162 -2066
rect 2168 -2078 2203 -2066
rect 1837 -2080 1999 -2078
rect 1732 -2108 1773 -2100
rect 1855 -2108 1868 -2080
rect 1883 -2082 1898 -2080
rect 1922 -2107 1929 -2100
rect 1932 -2108 1999 -2080
rect 2031 -2080 2203 -2078
rect 2001 -2102 2029 -2098
rect 2031 -2102 2111 -2080
rect 2132 -2082 2147 -2080
rect 2001 -2104 2111 -2102
rect 2001 -2108 2029 -2104
rect 2031 -2108 2111 -2104
rect 1638 -2118 1668 -2108
rect 1695 -2118 1696 -2108
rect 1711 -2118 1724 -2108
rect 1738 -2118 1739 -2108
rect 1754 -2118 1767 -2108
rect 1782 -2118 1812 -2108
rect 1855 -2118 1898 -2108
rect 1905 -2118 1913 -2108
rect 1932 -2116 1935 -2108
rect 1999 -2116 2031 -2108
rect 1932 -2118 2098 -2116
rect 2117 -2118 2128 -2108
rect 2132 -2118 2162 -2108
rect 2190 -2118 2203 -2080
rect 2275 -2074 2310 -2066
rect 2275 -2100 2276 -2074
rect 2283 -2100 2310 -2074
rect 2275 -2108 2310 -2100
rect 2312 -2074 2353 -2066
rect 2312 -2100 2327 -2074
rect 2334 -2100 2353 -2074
rect 2417 -2078 2479 -2066
rect 2491 -2078 2566 -2066
rect 2624 -2078 2699 -2066
rect 2711 -2078 2742 -2066
rect 2748 -2078 2783 -2066
rect 2417 -2080 2579 -2078
rect 2312 -2108 2353 -2100
rect 2435 -2108 2448 -2080
rect 2463 -2082 2478 -2080
rect 2502 -2107 2509 -2100
rect 2512 -2108 2579 -2080
rect 2611 -2080 2783 -2078
rect 2581 -2102 2609 -2098
rect 2611 -2102 2691 -2080
rect 2712 -2082 2727 -2080
rect 2581 -2104 2691 -2102
rect 2581 -2108 2609 -2104
rect 2611 -2108 2691 -2104
rect 2218 -2118 2248 -2108
rect 2275 -2118 2276 -2108
rect 2291 -2118 2304 -2108
rect 2318 -2118 2319 -2108
rect 2334 -2118 2347 -2108
rect 2362 -2118 2392 -2108
rect 2435 -2118 2478 -2108
rect 2485 -2118 2493 -2108
rect 2512 -2116 2515 -2108
rect 2579 -2116 2611 -2108
rect 2512 -2118 2678 -2116
rect 2697 -2118 2708 -2108
rect 2712 -2118 2742 -2108
rect 2770 -2118 2783 -2080
rect 2855 -2074 2890 -2066
rect 2855 -2100 2856 -2074
rect 2863 -2100 2890 -2074
rect 2855 -2108 2890 -2100
rect 2892 -2074 2933 -2066
rect 2892 -2100 2907 -2074
rect 2914 -2100 2933 -2074
rect 2997 -2078 3059 -2066
rect 3071 -2078 3146 -2066
rect 3204 -2078 3279 -2066
rect 3291 -2078 3322 -2066
rect 3328 -2078 3363 -2066
rect 2997 -2080 3159 -2078
rect 2892 -2108 2933 -2100
rect 3015 -2108 3028 -2080
rect 3043 -2082 3058 -2080
rect 3082 -2107 3089 -2100
rect 3092 -2108 3159 -2080
rect 3191 -2080 3363 -2078
rect 3161 -2102 3189 -2098
rect 3191 -2102 3271 -2080
rect 3292 -2082 3307 -2080
rect 3161 -2104 3271 -2102
rect 3161 -2108 3189 -2104
rect 3191 -2108 3271 -2104
rect 2798 -2118 2828 -2108
rect 2855 -2118 2856 -2108
rect 2871 -2118 2884 -2108
rect 2898 -2118 2899 -2108
rect 2914 -2118 2927 -2108
rect 2942 -2118 2972 -2108
rect 3015 -2118 3058 -2108
rect 3065 -2118 3073 -2108
rect 3092 -2116 3095 -2108
rect 3159 -2116 3191 -2108
rect 3092 -2118 3258 -2116
rect 3277 -2118 3288 -2108
rect 3292 -2118 3322 -2108
rect 3350 -2118 3363 -2080
rect 3435 -2074 3470 -2066
rect 3435 -2100 3436 -2074
rect 3443 -2100 3470 -2074
rect 3435 -2108 3470 -2100
rect 3472 -2074 3513 -2066
rect 3472 -2100 3487 -2074
rect 3494 -2100 3513 -2074
rect 3577 -2078 3639 -2066
rect 3651 -2078 3726 -2066
rect 3784 -2078 3859 -2066
rect 3871 -2078 3902 -2066
rect 3908 -2078 3943 -2066
rect 3577 -2080 3739 -2078
rect 3472 -2108 3513 -2100
rect 3595 -2108 3608 -2080
rect 3623 -2082 3638 -2080
rect 3662 -2107 3669 -2100
rect 3672 -2108 3739 -2080
rect 3771 -2080 3943 -2078
rect 3741 -2102 3769 -2098
rect 3771 -2102 3851 -2080
rect 3872 -2082 3887 -2080
rect 3741 -2104 3851 -2102
rect 3741 -2108 3769 -2104
rect 3771 -2108 3851 -2104
rect 3378 -2118 3408 -2108
rect 3435 -2118 3436 -2108
rect 3451 -2118 3464 -2108
rect 3478 -2118 3479 -2108
rect 3494 -2118 3507 -2108
rect 3522 -2118 3552 -2108
rect 3595 -2118 3638 -2108
rect 3645 -2118 3653 -2108
rect 3672 -2116 3675 -2108
rect 3739 -2116 3771 -2108
rect 3672 -2118 3838 -2116
rect 3857 -2118 3868 -2108
rect 3872 -2118 3902 -2108
rect 3930 -2118 3943 -2080
rect 4015 -2074 4050 -2066
rect 4015 -2100 4016 -2074
rect 4023 -2100 4050 -2074
rect 4015 -2108 4050 -2100
rect 4052 -2074 4093 -2066
rect 4052 -2100 4067 -2074
rect 4074 -2100 4093 -2074
rect 4157 -2078 4219 -2066
rect 4231 -2078 4306 -2066
rect 4364 -2078 4439 -2066
rect 4451 -2078 4482 -2066
rect 4488 -2078 4523 -2066
rect 4157 -2080 4319 -2078
rect 4052 -2108 4093 -2100
rect 4175 -2108 4188 -2080
rect 4203 -2082 4218 -2080
rect 4242 -2107 4249 -2100
rect 4252 -2108 4319 -2080
rect 4351 -2080 4523 -2078
rect 4321 -2102 4349 -2098
rect 4351 -2102 4431 -2080
rect 4452 -2082 4467 -2080
rect 4321 -2104 4431 -2102
rect 4321 -2108 4349 -2104
rect 4351 -2108 4431 -2104
rect 3958 -2118 3988 -2108
rect 4015 -2118 4016 -2108
rect 4031 -2118 4044 -2108
rect 4058 -2118 4059 -2108
rect 4074 -2118 4087 -2108
rect 4102 -2118 4132 -2108
rect 4175 -2118 4218 -2108
rect 4225 -2118 4233 -2108
rect 4252 -2116 4255 -2108
rect 4319 -2116 4351 -2108
rect 4252 -2118 4418 -2116
rect 4437 -2118 4448 -2108
rect 4452 -2118 4482 -2108
rect 4510 -2118 4523 -2080
rect 4595 -2074 4630 -2066
rect 4638 -2067 4639 -2051
rect 4654 -2067 4667 -2045
rect 4682 -2067 4712 -2045
rect 4755 -2049 4817 -2033
rect 4845 -2040 4856 -2024
rect 4861 -2029 4871 -2009
rect 4881 -2029 4895 -2009
rect 4898 -2022 4907 -2009
rect 4923 -2022 4932 -2009
rect 4861 -2040 4895 -2029
rect 4898 -2040 4907 -2024
rect 4923 -2040 4932 -2024
rect 4939 -2029 4949 -2009
rect 4959 -2029 4973 -2009
rect 4974 -2022 4985 -2009
rect 4939 -2040 4973 -2029
rect 4974 -2040 4985 -2024
rect 5031 -2033 5047 -2017
rect 5054 -2019 5084 -1967
rect 5118 -1971 5119 -1964
rect 5103 -1979 5119 -1971
rect 5090 -2011 5103 -1992
rect 5118 -2011 5148 -1995
rect 5090 -2027 5164 -2011
rect 5090 -2029 5103 -2027
rect 5118 -2029 5152 -2027
rect 4755 -2051 4768 -2049
rect 4783 -2051 4817 -2049
rect 4755 -2067 4817 -2051
rect 4861 -2056 4877 -2053
rect 4939 -2056 4969 -2045
rect 5017 -2049 5063 -2033
rect 5090 -2045 5164 -2029
rect 5017 -2051 5051 -2049
rect 5016 -2067 5063 -2051
rect 5090 -2067 5103 -2045
rect 5118 -2067 5148 -2045
rect 5175 -2067 5176 -2051
rect 5191 -2067 5204 -1907
rect 5234 -2011 5247 -1907
rect 5292 -1929 5293 -1919
rect 5313 -1921 5321 -1919
rect 5311 -1923 5321 -1921
rect 5308 -1929 5321 -1923
rect 5292 -1933 5321 -1929
rect 5326 -1933 5356 -1907
rect 5374 -1921 5390 -1919
rect 5462 -1921 5513 -1907
rect 5463 -1923 5527 -1921
rect 5374 -1933 5389 -1929
rect 5292 -1935 5389 -1933
rect 5276 -1943 5327 -1935
rect 5276 -1955 5301 -1943
rect 5308 -1955 5327 -1943
rect 5358 -1943 5408 -1935
rect 5358 -1951 5374 -1943
rect 5381 -1945 5408 -1943
rect 5417 -1943 5432 -1939
rect 5479 -1943 5511 -1923
rect 5570 -1935 5585 -1907
rect 5634 -1910 5664 -1907
rect 5634 -1913 5670 -1910
rect 5600 -1921 5616 -1919
rect 5601 -1933 5616 -1929
rect 5634 -1932 5673 -1913
rect 5692 -1919 5699 -1918
rect 5698 -1926 5699 -1919
rect 5682 -1929 5683 -1926
rect 5698 -1929 5711 -1926
rect 5634 -1933 5664 -1932
rect 5673 -1933 5679 -1932
rect 5682 -1933 5711 -1929
rect 5601 -1934 5711 -1933
rect 5601 -1935 5717 -1934
rect 5570 -1943 5638 -1935
rect 5417 -1945 5486 -1943
rect 5504 -1945 5638 -1943
rect 5381 -1949 5453 -1945
rect 5381 -1951 5506 -1949
rect 5381 -1955 5453 -1951
rect 5276 -1963 5327 -1955
rect 5374 -1959 5453 -1955
rect 5534 -1959 5638 -1945
rect 5667 -1943 5717 -1935
rect 5667 -1952 5683 -1943
rect 5374 -1963 5638 -1959
rect 5664 -1955 5683 -1952
rect 5690 -1955 5717 -1943
rect 5664 -1963 5717 -1955
rect 5292 -1971 5293 -1963
rect 5308 -1971 5321 -1963
rect 5292 -1979 5308 -1971
rect 5289 -1986 5308 -1983
rect 5289 -1995 5311 -1986
rect 5262 -2005 5311 -1995
rect 5262 -2011 5292 -2005
rect 5311 -2010 5316 -2005
rect 5234 -2027 5308 -2011
rect 5326 -2019 5356 -1963
rect 5391 -1973 5599 -1963
rect 5634 -1967 5679 -1963
rect 5682 -1964 5683 -1963
rect 5698 -1964 5711 -1963
rect 5558 -1977 5606 -1973
rect 5441 -1999 5471 -1990
rect 5534 -1997 5549 -1990
rect 5570 -1999 5606 -1977
rect 5417 -2003 5606 -1999
rect 5432 -2006 5606 -2003
rect 5425 -2009 5606 -2006
rect 5234 -2029 5247 -2027
rect 5262 -2029 5296 -2027
rect 5234 -2045 5308 -2029
rect 5335 -2033 5348 -2019
rect 5363 -2033 5379 -2017
rect 5425 -2022 5436 -2009
rect 5218 -2067 5219 -2051
rect 5234 -2067 5247 -2045
rect 5262 -2067 5292 -2045
rect 5335 -2049 5397 -2033
rect 5425 -2040 5436 -2024
rect 5441 -2029 5451 -2009
rect 5461 -2029 5475 -2009
rect 5478 -2022 5487 -2009
rect 5503 -2022 5512 -2009
rect 5441 -2040 5475 -2029
rect 5478 -2040 5487 -2024
rect 5503 -2040 5512 -2024
rect 5519 -2029 5529 -2009
rect 5539 -2029 5553 -2009
rect 5554 -2022 5565 -2009
rect 5519 -2040 5553 -2029
rect 5554 -2040 5565 -2024
rect 5611 -2033 5627 -2017
rect 5634 -2019 5664 -1967
rect 5698 -1971 5699 -1964
rect 5683 -1979 5699 -1971
rect 5670 -2011 5683 -1992
rect 5698 -2011 5728 -1995
rect 5670 -2027 5744 -2011
rect 5670 -2029 5683 -2027
rect 5698 -2029 5732 -2027
rect 5335 -2051 5348 -2049
rect 5363 -2051 5397 -2049
rect 5335 -2067 5397 -2051
rect 5441 -2056 5457 -2053
rect 5519 -2056 5549 -2045
rect 5597 -2049 5643 -2033
rect 5670 -2045 5744 -2029
rect 5597 -2051 5631 -2049
rect 5596 -2067 5643 -2051
rect 5670 -2067 5683 -2045
rect 5698 -2067 5728 -2045
rect 5755 -2067 5756 -2051
rect 5771 -2067 5784 -1907
rect 5814 -2011 5827 -1907
rect 5872 -1929 5873 -1919
rect 5893 -1921 5901 -1919
rect 5891 -1923 5901 -1921
rect 5888 -1929 5901 -1923
rect 5872 -1933 5901 -1929
rect 5906 -1933 5936 -1907
rect 5954 -1921 5970 -1919
rect 6042 -1921 6093 -1907
rect 6043 -1923 6107 -1921
rect 5954 -1933 5969 -1929
rect 5872 -1935 5969 -1933
rect 5856 -1943 5907 -1935
rect 5856 -1955 5881 -1943
rect 5888 -1955 5907 -1943
rect 5938 -1943 5988 -1935
rect 5938 -1951 5954 -1943
rect 5961 -1945 5988 -1943
rect 5997 -1943 6012 -1939
rect 6059 -1943 6091 -1923
rect 6150 -1935 6165 -1907
rect 6214 -1910 6244 -1907
rect 6214 -1913 6250 -1910
rect 6180 -1921 6196 -1919
rect 6181 -1933 6196 -1929
rect 6214 -1932 6253 -1913
rect 6272 -1919 6279 -1918
rect 6278 -1926 6279 -1919
rect 6262 -1929 6263 -1926
rect 6278 -1929 6291 -1926
rect 6214 -1933 6244 -1932
rect 6253 -1933 6259 -1932
rect 6262 -1933 6291 -1929
rect 6181 -1934 6291 -1933
rect 6181 -1935 6297 -1934
rect 6150 -1943 6218 -1935
rect 5997 -1945 6066 -1943
rect 6084 -1945 6218 -1943
rect 5961 -1949 6033 -1945
rect 5961 -1951 6086 -1949
rect 5961 -1955 6033 -1951
rect 5856 -1963 5907 -1955
rect 5954 -1959 6033 -1955
rect 6114 -1959 6218 -1945
rect 6247 -1943 6297 -1935
rect 6247 -1952 6263 -1943
rect 5954 -1963 6218 -1959
rect 6244 -1955 6263 -1952
rect 6270 -1955 6297 -1943
rect 6244 -1963 6297 -1955
rect 5872 -1971 5873 -1963
rect 5888 -1971 5901 -1963
rect 5872 -1979 5888 -1971
rect 5869 -1986 5888 -1983
rect 5869 -1995 5891 -1986
rect 5842 -2005 5891 -1995
rect 5842 -2011 5872 -2005
rect 5891 -2010 5896 -2005
rect 5814 -2027 5888 -2011
rect 5906 -2019 5936 -1963
rect 5971 -1973 6179 -1963
rect 6214 -1967 6259 -1963
rect 6262 -1964 6263 -1963
rect 6278 -1964 6291 -1963
rect 6138 -1977 6186 -1973
rect 6021 -1999 6051 -1990
rect 6114 -1997 6129 -1990
rect 6150 -1999 6186 -1977
rect 5997 -2003 6186 -1999
rect 6012 -2006 6186 -2003
rect 6005 -2009 6186 -2006
rect 5814 -2029 5827 -2027
rect 5842 -2029 5876 -2027
rect 5814 -2045 5888 -2029
rect 5915 -2033 5928 -2019
rect 5943 -2033 5959 -2017
rect 6005 -2022 6016 -2009
rect 5798 -2067 5799 -2051
rect 5814 -2067 5827 -2045
rect 5842 -2067 5872 -2045
rect 5915 -2049 5977 -2033
rect 6005 -2040 6016 -2024
rect 6021 -2029 6031 -2009
rect 6041 -2029 6055 -2009
rect 6058 -2022 6067 -2009
rect 6083 -2022 6092 -2009
rect 6021 -2040 6055 -2029
rect 6058 -2040 6067 -2024
rect 6083 -2040 6092 -2024
rect 6099 -2029 6109 -2009
rect 6119 -2029 6133 -2009
rect 6134 -2022 6145 -2009
rect 6099 -2040 6133 -2029
rect 6134 -2040 6145 -2024
rect 6191 -2033 6207 -2017
rect 6214 -2019 6244 -1967
rect 6278 -1971 6279 -1964
rect 6263 -1979 6279 -1971
rect 6250 -2011 6263 -1992
rect 6278 -2011 6308 -1995
rect 6250 -2027 6324 -2011
rect 6250 -2029 6263 -2027
rect 6278 -2029 6312 -2027
rect 5915 -2051 5928 -2049
rect 5943 -2051 5977 -2049
rect 5915 -2067 5977 -2051
rect 6021 -2056 6037 -2053
rect 6099 -2056 6129 -2045
rect 6177 -2049 6223 -2033
rect 6250 -2045 6324 -2029
rect 6177 -2051 6211 -2049
rect 6176 -2067 6223 -2051
rect 6250 -2067 6263 -2045
rect 6278 -2067 6308 -2045
rect 6335 -2067 6336 -2051
rect 6351 -2067 6364 -1907
rect 6394 -2011 6407 -1907
rect 6452 -1929 6453 -1919
rect 6473 -1921 6481 -1919
rect 6471 -1923 6481 -1921
rect 6468 -1929 6481 -1923
rect 6452 -1933 6481 -1929
rect 6486 -1933 6516 -1907
rect 6534 -1921 6550 -1919
rect 6622 -1921 6673 -1907
rect 6623 -1923 6687 -1921
rect 6534 -1933 6549 -1929
rect 6452 -1935 6549 -1933
rect 6436 -1943 6487 -1935
rect 6436 -1955 6461 -1943
rect 6468 -1955 6487 -1943
rect 6518 -1943 6568 -1935
rect 6518 -1951 6534 -1943
rect 6541 -1945 6568 -1943
rect 6577 -1943 6592 -1939
rect 6639 -1943 6671 -1923
rect 6730 -1935 6745 -1907
rect 6794 -1910 6824 -1907
rect 6794 -1913 6830 -1910
rect 6760 -1921 6776 -1919
rect 6761 -1933 6776 -1929
rect 6794 -1932 6833 -1913
rect 6852 -1919 6859 -1918
rect 6858 -1926 6859 -1919
rect 6842 -1929 6843 -1926
rect 6858 -1929 6871 -1926
rect 6794 -1933 6824 -1932
rect 6833 -1933 6839 -1932
rect 6842 -1933 6871 -1929
rect 6761 -1934 6871 -1933
rect 6761 -1935 6877 -1934
rect 6730 -1943 6798 -1935
rect 6577 -1945 6646 -1943
rect 6664 -1945 6798 -1943
rect 6541 -1949 6613 -1945
rect 6541 -1951 6666 -1949
rect 6541 -1955 6613 -1951
rect 6436 -1963 6487 -1955
rect 6534 -1959 6613 -1955
rect 6694 -1959 6798 -1945
rect 6827 -1943 6877 -1935
rect 6827 -1952 6843 -1943
rect 6534 -1963 6798 -1959
rect 6824 -1955 6843 -1952
rect 6850 -1955 6877 -1943
rect 6824 -1963 6877 -1955
rect 6452 -1971 6453 -1963
rect 6468 -1971 6481 -1963
rect 6452 -1979 6468 -1971
rect 6449 -1986 6468 -1983
rect 6449 -1995 6471 -1986
rect 6422 -2005 6471 -1995
rect 6422 -2011 6452 -2005
rect 6471 -2010 6476 -2005
rect 6394 -2027 6468 -2011
rect 6486 -2019 6516 -1963
rect 6551 -1973 6759 -1963
rect 6794 -1967 6839 -1963
rect 6842 -1964 6843 -1963
rect 6858 -1964 6871 -1963
rect 6718 -1977 6766 -1973
rect 6601 -1999 6631 -1990
rect 6694 -1997 6709 -1990
rect 6730 -1999 6766 -1977
rect 6577 -2003 6766 -1999
rect 6592 -2006 6766 -2003
rect 6585 -2009 6766 -2006
rect 6394 -2029 6407 -2027
rect 6422 -2029 6456 -2027
rect 6394 -2045 6468 -2029
rect 6495 -2033 6508 -2019
rect 6523 -2033 6539 -2017
rect 6585 -2022 6596 -2009
rect 6378 -2067 6379 -2051
rect 6394 -2067 6407 -2045
rect 6422 -2067 6452 -2045
rect 6495 -2049 6557 -2033
rect 6585 -2040 6596 -2024
rect 6601 -2029 6611 -2009
rect 6621 -2029 6635 -2009
rect 6638 -2022 6647 -2009
rect 6663 -2022 6672 -2009
rect 6601 -2040 6635 -2029
rect 6638 -2040 6647 -2024
rect 6663 -2040 6672 -2024
rect 6679 -2029 6689 -2009
rect 6699 -2029 6713 -2009
rect 6714 -2022 6725 -2009
rect 6679 -2040 6713 -2029
rect 6714 -2040 6725 -2024
rect 6771 -2033 6787 -2017
rect 6794 -2019 6824 -1967
rect 6858 -1971 6859 -1964
rect 6843 -1979 6859 -1971
rect 6830 -2011 6843 -1992
rect 6858 -2011 6888 -1995
rect 6830 -2027 6904 -2011
rect 6830 -2029 6843 -2027
rect 6858 -2029 6892 -2027
rect 6495 -2051 6508 -2049
rect 6523 -2051 6557 -2049
rect 6495 -2067 6557 -2051
rect 6601 -2056 6617 -2053
rect 6679 -2056 6709 -2045
rect 6757 -2049 6803 -2033
rect 6830 -2045 6904 -2029
rect 6757 -2051 6791 -2049
rect 6756 -2067 6803 -2051
rect 6830 -2067 6843 -2045
rect 6858 -2067 6888 -2045
rect 6915 -2067 6916 -2051
rect 6931 -2067 6944 -1907
rect 4595 -2100 4596 -2074
rect 4603 -2100 4630 -2074
rect 4595 -2108 4630 -2100
rect 4632 -2075 4673 -2067
rect 4632 -2101 4647 -2075
rect 4654 -2101 4673 -2075
rect 4737 -2079 4799 -2067
rect 4811 -2079 4886 -2067
rect 4944 -2079 5019 -2067
rect 5031 -2079 5062 -2067
rect 5068 -2079 5103 -2067
rect 4737 -2081 4899 -2079
rect 4538 -2118 4568 -2108
rect 4595 -2118 4596 -2108
rect 4611 -2118 4624 -2108
rect 4632 -2109 4673 -2101
rect 4755 -2109 4768 -2081
rect 4783 -2083 4798 -2081
rect 4832 -2099 4899 -2081
rect 4931 -2081 5103 -2079
rect 4931 -2099 5011 -2081
rect 5032 -2083 5047 -2081
rect 4822 -2108 4829 -2101
rect 4832 -2109 5011 -2099
rect 0 -2119 4624 -2118
rect 4638 -2119 4639 -2109
rect 4654 -2119 4667 -2109
rect 4682 -2119 4712 -2109
rect 4755 -2119 4798 -2109
rect 4805 -2119 4813 -2109
rect 4832 -2117 4835 -2109
rect 4899 -2117 4931 -2109
rect 4832 -2119 4998 -2117
rect 5017 -2119 5028 -2109
rect 5032 -2119 5062 -2109
rect 5090 -2119 5103 -2081
rect 5175 -2075 5210 -2067
rect 5175 -2101 5176 -2075
rect 5183 -2101 5210 -2075
rect 5175 -2109 5210 -2101
rect 5212 -2075 5253 -2067
rect 5212 -2101 5227 -2075
rect 5234 -2101 5253 -2075
rect 5317 -2079 5379 -2067
rect 5391 -2079 5466 -2067
rect 5524 -2079 5599 -2067
rect 5611 -2079 5642 -2067
rect 5648 -2079 5683 -2067
rect 5317 -2081 5479 -2079
rect 5212 -2109 5253 -2101
rect 5335 -2109 5348 -2081
rect 5363 -2083 5378 -2081
rect 5412 -2099 5479 -2081
rect 5511 -2081 5683 -2079
rect 5511 -2099 5591 -2081
rect 5612 -2083 5627 -2081
rect 5402 -2108 5409 -2101
rect 5412 -2109 5591 -2099
rect 5118 -2119 5148 -2109
rect 5175 -2119 5176 -2109
rect 5191 -2119 5204 -2109
rect 5218 -2119 5219 -2109
rect 5234 -2119 5247 -2109
rect 5262 -2119 5292 -2109
rect 5335 -2119 5378 -2109
rect 5385 -2119 5393 -2109
rect 5412 -2117 5415 -2109
rect 5479 -2117 5511 -2109
rect 5412 -2119 5578 -2117
rect 5597 -2119 5608 -2109
rect 5612 -2119 5642 -2109
rect 5670 -2119 5683 -2081
rect 5755 -2075 5790 -2067
rect 5755 -2101 5756 -2075
rect 5763 -2101 5790 -2075
rect 5755 -2109 5790 -2101
rect 5792 -2075 5833 -2067
rect 5792 -2101 5807 -2075
rect 5814 -2101 5833 -2075
rect 5897 -2079 5959 -2067
rect 5971 -2079 6046 -2067
rect 6104 -2079 6179 -2067
rect 6191 -2079 6222 -2067
rect 6228 -2079 6263 -2067
rect 5897 -2081 6059 -2079
rect 5792 -2109 5833 -2101
rect 5915 -2109 5928 -2081
rect 5943 -2083 5958 -2081
rect 5992 -2099 6059 -2081
rect 6091 -2081 6263 -2079
rect 6091 -2099 6171 -2081
rect 6192 -2083 6207 -2081
rect 5982 -2108 5989 -2101
rect 5992 -2109 6171 -2099
rect 5698 -2119 5728 -2109
rect 5755 -2119 5756 -2109
rect 5771 -2119 5784 -2109
rect 5798 -2119 5799 -2109
rect 5814 -2119 5827 -2109
rect 5842 -2119 5872 -2109
rect 5915 -2119 5958 -2109
rect 5965 -2119 5973 -2109
rect 5992 -2117 5995 -2109
rect 6059 -2117 6091 -2109
rect 5992 -2119 6158 -2117
rect 6177 -2119 6188 -2109
rect 6192 -2119 6222 -2109
rect 6250 -2119 6263 -2081
rect 6335 -2075 6370 -2067
rect 6335 -2101 6336 -2075
rect 6343 -2101 6370 -2075
rect 6335 -2109 6370 -2101
rect 6372 -2075 6413 -2067
rect 6372 -2101 6387 -2075
rect 6394 -2101 6413 -2075
rect 6477 -2079 6539 -2067
rect 6551 -2079 6626 -2067
rect 6684 -2079 6759 -2067
rect 6771 -2079 6802 -2067
rect 6808 -2079 6843 -2067
rect 6477 -2081 6639 -2079
rect 6372 -2109 6413 -2101
rect 6495 -2109 6508 -2081
rect 6523 -2083 6538 -2081
rect 6572 -2099 6639 -2081
rect 6671 -2081 6843 -2079
rect 6671 -2099 6751 -2081
rect 6772 -2083 6787 -2081
rect 6562 -2108 6569 -2101
rect 6572 -2109 6751 -2099
rect 6278 -2119 6308 -2109
rect 6335 -2119 6336 -2109
rect 6351 -2119 6364 -2109
rect 6378 -2119 6379 -2109
rect 6394 -2119 6407 -2109
rect 6422 -2119 6452 -2109
rect 6495 -2119 6538 -2109
rect 6545 -2119 6553 -2109
rect 6572 -2117 6575 -2109
rect 6639 -2117 6671 -2109
rect 6572 -2119 6738 -2117
rect 6757 -2119 6768 -2109
rect 6772 -2119 6802 -2109
rect 6830 -2119 6843 -2081
rect 6915 -2075 6950 -2067
rect 6915 -2101 6916 -2075
rect 6923 -2101 6950 -2075
rect 6915 -2109 6950 -2101
rect 6858 -2119 6888 -2109
rect 6915 -2119 6916 -2109
rect 6931 -2119 6944 -2109
rect 0 -2132 6944 -2119
rect 14 -2146 27 -2132
rect 42 -2150 72 -2132
rect 115 -2146 128 -2132
rect 165 -2145 173 -2132
rect 206 -2145 344 -2132
rect 377 -2145 385 -2132
rect 242 -2146 293 -2145
rect 450 -2146 463 -2132
rect 243 -2148 307 -2146
rect 478 -2150 508 -2132
rect 551 -2146 564 -2132
rect 594 -2146 607 -2132
rect 622 -2150 652 -2132
rect 695 -2146 708 -2132
rect 745 -2145 753 -2132
rect 786 -2145 924 -2132
rect 957 -2145 965 -2132
rect 822 -2146 873 -2145
rect 1030 -2146 1043 -2132
rect 823 -2148 887 -2146
rect 1058 -2150 1088 -2132
rect 1131 -2146 1144 -2132
rect 1174 -2146 1187 -2132
rect 1202 -2150 1232 -2132
rect 1275 -2146 1288 -2132
rect 1325 -2145 1333 -2132
rect 1366 -2145 1504 -2132
rect 1537 -2145 1545 -2132
rect 1402 -2146 1453 -2145
rect 1610 -2146 1623 -2132
rect 1403 -2148 1467 -2146
rect 1638 -2150 1668 -2132
rect 1711 -2146 1724 -2132
rect 1754 -2146 1767 -2132
rect 1782 -2150 1812 -2132
rect 1855 -2146 1868 -2132
rect 1905 -2145 1913 -2132
rect 1946 -2145 2084 -2132
rect 2117 -2145 2125 -2132
rect 1982 -2146 2033 -2145
rect 2190 -2146 2203 -2132
rect 1983 -2148 2047 -2146
rect 2218 -2150 2248 -2132
rect 2291 -2146 2304 -2132
rect 2334 -2146 2347 -2132
rect 2362 -2150 2392 -2132
rect 2435 -2146 2448 -2132
rect 2485 -2145 2493 -2132
rect 2526 -2145 2664 -2132
rect 2697 -2145 2705 -2132
rect 2562 -2146 2613 -2145
rect 2770 -2146 2783 -2132
rect 2563 -2148 2627 -2146
rect 2798 -2150 2828 -2132
rect 2871 -2146 2884 -2132
rect 2914 -2146 2927 -2132
rect 2942 -2150 2972 -2132
rect 3015 -2146 3028 -2132
rect 3065 -2145 3073 -2132
rect 3106 -2145 3244 -2132
rect 3277 -2145 3285 -2132
rect 3142 -2146 3193 -2145
rect 3350 -2146 3363 -2132
rect 3143 -2148 3205 -2146
rect 3378 -2150 3408 -2132
rect 3451 -2146 3464 -2132
rect 3494 -2146 3507 -2132
rect 3522 -2150 3552 -2132
rect 3595 -2146 3608 -2132
rect 3645 -2145 3653 -2132
rect 3686 -2145 3824 -2132
rect 3857 -2145 3865 -2132
rect 3722 -2146 3773 -2145
rect 3930 -2146 3943 -2132
rect 3723 -2148 3787 -2146
rect 3958 -2150 3988 -2132
rect 4031 -2146 4044 -2132
rect 4074 -2146 4087 -2132
rect 4102 -2150 4132 -2132
rect 4175 -2146 4188 -2132
rect 4225 -2145 4233 -2132
rect 4266 -2145 4404 -2132
rect 4437 -2145 4445 -2132
rect 4302 -2146 4353 -2145
rect 4510 -2146 4523 -2132
rect 4303 -2148 4367 -2146
rect 4538 -2150 4568 -2132
rect 4611 -2133 6944 -2132
rect 4611 -2146 4624 -2133
rect 4654 -2195 4667 -2133
rect 4682 -2151 4712 -2133
rect 4755 -2147 4768 -2133
rect 4805 -2146 4813 -2133
rect 4846 -2146 4984 -2133
rect 5017 -2146 5025 -2133
rect 4882 -2147 4933 -2146
rect 5090 -2147 5103 -2133
rect 4899 -2149 4931 -2147
rect 5118 -2151 5148 -2133
rect 5191 -2195 5204 -2133
rect 5234 -2195 5247 -2133
rect 5262 -2151 5292 -2133
rect 5335 -2147 5348 -2133
rect 5385 -2146 5393 -2133
rect 5426 -2146 5564 -2133
rect 5597 -2146 5605 -2133
rect 5462 -2147 5513 -2146
rect 5670 -2147 5683 -2133
rect 5479 -2149 5511 -2147
rect 5698 -2151 5728 -2133
rect 5771 -2195 5784 -2133
rect 5814 -2195 5827 -2133
rect 5842 -2151 5872 -2133
rect 5915 -2147 5928 -2133
rect 5965 -2146 5973 -2133
rect 6006 -2146 6144 -2133
rect 6177 -2146 6185 -2133
rect 6042 -2147 6093 -2146
rect 6250 -2147 6263 -2133
rect 6059 -2149 6091 -2147
rect 6278 -2151 6308 -2133
rect 6351 -2195 6364 -2133
rect 6394 -2195 6407 -2133
rect 6422 -2151 6452 -2133
rect 6495 -2147 6508 -2133
rect 6545 -2146 6553 -2133
rect 6586 -2146 6724 -2133
rect 6757 -2146 6765 -2133
rect 6622 -2147 6673 -2146
rect 6830 -2147 6843 -2133
rect 6639 -2149 6671 -2147
rect 6858 -2151 6888 -2133
rect 6931 -2195 6944 -2133
<< pwell >>
rect 4568 2006 4593 2040
rect 4568 1736 4591 1770
<< metal1 >>
rect 4568 2006 4593 2040
rect 4568 1736 4591 1770
use 10T_4x4_magic  10T_4x4_magic_0
timestamp 1667336911
transform 1 0 4645 0 1 819
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_1
timestamp 1667336911
transform 1 0 4645 0 1 1900
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_2
timestamp 1667336911
transform 1 0 4645 0 1 1360
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_3
timestamp 1667336911
transform 1 0 4645 0 1 279
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_4
timestamp 1667336911
transform 1 0 4645 0 1 -261
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_5
timestamp 1667336911
transform 1 0 4645 0 1 -801
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_6
timestamp 1667336911
transform 1 0 4645 0 1 -1341
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_7
timestamp 1667336911
transform 1 0 4645 0 1 -1881
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_8
timestamp 1667336911
transform 1 0 5805 0 1 279
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_9
timestamp 1667336911
transform 1 0 5805 0 1 -261
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_10
timestamp 1667336911
transform 1 0 5805 0 1 -801
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_11
timestamp 1667336911
transform 1 0 5805 0 1 -1341
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_12
timestamp 1667336911
transform 1 0 5805 0 1 -1881
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_13
timestamp 1667336911
transform 1 0 5805 0 1 819
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_14
timestamp 1667336911
transform 1 0 5805 0 1 1900
box -54 -314 1145 322
use 10T_4x4_magic  10T_4x4_magic_15
timestamp 1667336911
transform 1 0 5805 0 1 1360
box -54 -314 1145 322
use 10T_8x8_magic  10T_8x8_magic_0
timestamp 1667336911
transform 1 0 -1 0 1 1094
box -7 -1084 4631 1122
use 10T_8x8_magic  10T_8x8_magic_1
timestamp 1667336911
transform 1 0 -1 0 1 -1066
box -7 -1084 4631 1122
<< end >>
