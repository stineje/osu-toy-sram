** sch_path: /home/rjridle/osu-toy-sram/custom_layout/xschsky130_fd_bd_sram__sram_sp_cell.sch

** INV 0
Mppu_2   left_net  right_net VPWR      PWELL ppu   L=0.15  W=0.14
Mnpd_1   left_net  right_net VGND      VSUBS npd   L=0.15  W=0.21

** INV 1
Mppu_1   right_net left_net  VPWR      PWELL ppu   L=0.15  W=0.14
Mnpd_0   right_net left_net  VGND      VSUBS npd   L=0.15  W=0.21

** Left side
Mppu_3   left_net  WL1       left_net  PWELL ppu   L=0.095 W=0.07 
Mnpass_1 left_net  WL1       bit_v     VSUBS npass L=0.15  W=0.14 

** Right Side
Mppu_0   right_net WL2       right_net PWELL ppu   L=0.095 W=0.07
Mnpass_0 right_net WL2       bit_b_v   VSUBS npass L=0.15  W=0.14
