magic
tech sky130A
magscale 1 2
timestamp 1675183705
<< nwell >>
rect 191 4187 344 4283
rect 771 4187 924 4283
rect 191 3917 344 4013
rect 771 3917 924 4013
rect 191 3647 344 3743
rect 771 3647 924 3743
rect 191 3377 344 3473
rect 771 3377 924 3473
rect 191 3107 344 3203
rect 771 3107 924 3203
rect 191 2837 344 2933
rect 771 2837 924 2933
rect 191 2567 344 2663
rect 771 2567 924 2663
rect 191 2297 344 2393
rect 771 2297 924 2393
rect 191 2027 344 2123
rect 771 2027 924 2123
rect 191 1757 344 1853
rect 771 1757 924 1853
rect 191 1487 344 1583
rect 771 1487 924 1583
rect 191 1217 344 1313
rect 771 1217 924 1313
rect 191 947 344 1043
rect 771 947 924 1043
rect 191 677 344 773
rect 771 677 924 773
rect 191 407 344 503
rect 771 407 924 503
rect 191 137 344 233
rect 771 137 924 233
rect 1351 4187 1504 4283
rect 1931 4187 2084 4283
rect 1351 3917 1504 4013
rect 1931 3917 2084 4013
rect 1351 3647 1504 3743
rect 1931 3647 2084 3743
rect 1351 3377 1504 3473
rect 1931 3377 2084 3473
rect 1351 3107 1504 3203
rect 1931 3107 2084 3203
rect 1351 2837 1504 2933
rect 1931 2837 2084 2933
rect 1351 2567 1504 2663
rect 1931 2567 2084 2663
rect 1351 2297 1504 2393
rect 1931 2297 2084 2393
rect 1351 2027 1504 2123
rect 1931 2027 2084 2123
rect 1351 1757 1504 1853
rect 1931 1757 2084 1853
rect 1351 1487 1504 1583
rect 1931 1487 2084 1583
rect 1351 1217 1504 1313
rect 1931 1217 2084 1313
rect 1351 947 1504 1043
rect 1931 947 2084 1043
rect 1351 677 1504 773
rect 1931 677 2084 773
rect 1351 407 1504 503
rect 1931 407 2084 503
rect 1351 137 1504 233
rect 1931 137 2084 233
rect 2511 4187 2664 4283
rect 3091 4187 3244 4283
rect 2511 3917 2664 4013
rect 3091 3917 3244 4013
rect 2511 3647 2664 3743
rect 3091 3647 3244 3743
rect 2511 3377 2664 3473
rect 3091 3377 3244 3473
rect 2511 3107 2664 3203
rect 3091 3107 3244 3203
rect 2511 2837 2664 2933
rect 3091 2837 3244 2933
rect 2511 2567 2664 2663
rect 3091 2567 3244 2663
rect 2511 2297 2664 2393
rect 3091 2297 3244 2393
rect 2511 2027 2664 2123
rect 3091 2027 3244 2123
rect 2511 1757 2664 1853
rect 3091 1757 3244 1853
rect 2511 1487 2664 1583
rect 3091 1487 3244 1583
rect 2511 1217 2664 1313
rect 3091 1217 3244 1313
rect 2511 947 2664 1043
rect 3091 947 3244 1043
rect 2511 677 2664 773
rect 3091 677 3244 773
rect 2511 407 2664 503
rect 3091 407 3244 503
rect 2511 137 2664 233
rect 3091 137 3244 233
rect 3671 4187 3824 4283
rect 4251 4187 4404 4283
rect 3671 3917 3824 4013
rect 4251 3917 4404 4013
rect 3671 3647 3824 3743
rect 4251 3647 4404 3743
rect 3671 3377 3824 3473
rect 4251 3377 4404 3473
rect 3671 3107 3824 3203
rect 4251 3107 4404 3203
rect 3671 2837 3824 2933
rect 4251 2837 4404 2933
rect 3671 2567 3824 2663
rect 4251 2567 4404 2663
rect 3671 2297 3824 2393
rect 4251 2297 4404 2393
rect 3671 2027 3824 2123
rect 4251 2027 4404 2123
rect 3671 1757 3824 1853
rect 4251 1757 4404 1853
rect 3671 1487 3824 1583
rect 4251 1487 4404 1583
rect 3671 1217 3824 1313
rect 4251 1217 4404 1313
rect 3671 947 3824 1043
rect 4251 947 4404 1043
rect 3671 677 3824 773
rect 4251 677 4404 773
rect 3671 407 3824 503
rect 4251 407 4404 503
rect 3671 137 3824 233
rect 4251 137 4404 233
rect 4831 4187 4984 4283
rect 5411 4187 5564 4283
rect 4831 3917 4984 4013
rect 5411 3917 5564 4013
rect 4831 3647 4984 3743
rect 5411 3647 5564 3743
rect 4831 3377 4984 3473
rect 5411 3377 5564 3473
rect 4831 3107 4984 3203
rect 5411 3107 5564 3203
rect 4831 2837 4984 2933
rect 5411 2837 5564 2933
rect 4831 2567 4984 2663
rect 5411 2567 5564 2663
rect 4831 2297 4984 2393
rect 5411 2297 5564 2393
rect 4831 2027 4984 2123
rect 5411 2027 5564 2123
rect 4831 1757 4984 1853
rect 5411 1757 5564 1853
rect 4831 1487 4984 1583
rect 5411 1487 5564 1583
rect 4831 1217 4984 1313
rect 5411 1217 5564 1313
rect 4831 947 4984 1043
rect 5411 947 5564 1043
rect 4831 677 4984 773
rect 5411 677 5564 773
rect 4831 407 4984 503
rect 5411 407 5564 503
rect 4831 137 4984 233
rect 5411 137 5564 233
rect 5991 4187 6144 4283
rect 6571 4187 6724 4283
rect 5991 3917 6144 4013
rect 6571 3917 6724 4013
rect 5991 3647 6144 3743
rect 6571 3647 6724 3743
rect 5991 3377 6144 3473
rect 6571 3377 6724 3473
rect 5991 3107 6144 3203
rect 6571 3107 6724 3203
rect 5991 2837 6144 2933
rect 6571 2837 6724 2933
rect 5991 2567 6144 2663
rect 6571 2567 6724 2663
rect 5991 2297 6144 2393
rect 6571 2297 6724 2393
rect 5991 2027 6144 2123
rect 6571 2027 6724 2123
rect 5991 1757 6144 1853
rect 6571 1757 6724 1853
rect 5991 1487 6144 1583
rect 6571 1487 6724 1583
rect 5991 1217 6144 1313
rect 6571 1217 6724 1313
rect 5991 947 6144 1043
rect 6571 947 6724 1043
rect 5991 677 6144 773
rect 6571 677 6724 773
rect 5991 407 6144 503
rect 6571 407 6724 503
rect 5991 137 6144 233
rect 6571 137 6724 233
<< pwell >>
rect -7 4141 163 4313
rect 375 4141 743 4313
rect 955 4141 1125 4313
rect -7 4043 1125 4141
rect -7 3871 163 4043
rect 375 3871 743 4043
rect 955 3871 1125 4043
rect -7 3773 1125 3871
rect -7 3601 163 3773
rect 375 3601 743 3773
rect 955 3601 1125 3773
rect -7 3503 1125 3601
rect -7 3331 163 3503
rect 375 3331 743 3503
rect 955 3331 1125 3503
rect -7 3233 1125 3331
rect -7 3061 163 3233
rect 375 3061 743 3233
rect 955 3061 1125 3233
rect -7 2963 1125 3061
rect -7 2791 163 2963
rect 375 2791 743 2963
rect 955 2791 1125 2963
rect -7 2693 1125 2791
rect -7 2521 163 2693
rect 375 2521 743 2693
rect 955 2521 1125 2693
rect -7 2423 1125 2521
rect -7 2251 163 2423
rect 375 2251 743 2423
rect 955 2251 1125 2423
rect -7 2153 1125 2251
rect -7 1981 163 2153
rect 375 1981 743 2153
rect 955 1981 1125 2153
rect -7 1883 1125 1981
rect -7 1711 163 1883
rect 375 1711 743 1883
rect 955 1711 1125 1883
rect -7 1613 1125 1711
rect -7 1441 163 1613
rect 375 1441 743 1613
rect 955 1441 1125 1613
rect -7 1343 1125 1441
rect -7 1171 163 1343
rect 375 1171 743 1343
rect 955 1171 1125 1343
rect -7 1073 1125 1171
rect -7 901 163 1073
rect 375 901 743 1073
rect 955 901 1125 1073
rect -7 803 1125 901
rect -7 631 163 803
rect 375 631 743 803
rect 955 631 1125 803
rect -7 533 1125 631
rect -7 361 163 533
rect 375 361 743 533
rect 955 361 1125 533
rect -7 263 1125 361
rect -7 91 163 263
rect 375 91 743 263
rect 955 91 1125 263
rect -7 -7 1125 91
rect 1153 4141 1323 4313
rect 1535 4141 1903 4313
rect 2115 4141 2285 4313
rect 1153 4043 2285 4141
rect 1153 3871 1323 4043
rect 1535 3871 1903 4043
rect 2115 3871 2285 4043
rect 1153 3773 2285 3871
rect 1153 3601 1323 3773
rect 1535 3601 1903 3773
rect 2115 3601 2285 3773
rect 1153 3503 2285 3601
rect 1153 3331 1323 3503
rect 1535 3331 1903 3503
rect 2115 3331 2285 3503
rect 1153 3233 2285 3331
rect 1153 3061 1323 3233
rect 1535 3061 1903 3233
rect 2115 3061 2285 3233
rect 1153 2963 2285 3061
rect 1153 2791 1323 2963
rect 1535 2791 1903 2963
rect 2115 2791 2285 2963
rect 1153 2693 2285 2791
rect 1153 2521 1323 2693
rect 1535 2521 1903 2693
rect 2115 2521 2285 2693
rect 1153 2423 2285 2521
rect 1153 2251 1323 2423
rect 1535 2251 1903 2423
rect 2115 2251 2285 2423
rect 1153 2153 2285 2251
rect 1153 1981 1323 2153
rect 1535 1981 1903 2153
rect 2115 1981 2285 2153
rect 1153 1883 2285 1981
rect 1153 1711 1323 1883
rect 1535 1711 1903 1883
rect 2115 1711 2285 1883
rect 1153 1613 2285 1711
rect 1153 1441 1323 1613
rect 1535 1441 1903 1613
rect 2115 1441 2285 1613
rect 1153 1343 2285 1441
rect 1153 1171 1323 1343
rect 1535 1171 1903 1343
rect 2115 1171 2285 1343
rect 1153 1073 2285 1171
rect 1153 901 1323 1073
rect 1535 901 1903 1073
rect 2115 901 2285 1073
rect 1153 803 2285 901
rect 1153 631 1323 803
rect 1535 631 1903 803
rect 2115 631 2285 803
rect 1153 533 2285 631
rect 1153 361 1323 533
rect 1535 361 1903 533
rect 2115 361 2285 533
rect 1153 263 2285 361
rect 1153 91 1323 263
rect 1535 91 1903 263
rect 2115 91 2285 263
rect 1153 -7 2285 91
rect 2313 4141 2483 4313
rect 2695 4141 3063 4313
rect 3275 4141 3445 4313
rect 2313 4043 3445 4141
rect 2313 3871 2483 4043
rect 2695 3871 3063 4043
rect 3275 3871 3445 4043
rect 2313 3773 3445 3871
rect 2313 3601 2483 3773
rect 2695 3601 3063 3773
rect 3275 3601 3445 3773
rect 2313 3503 3445 3601
rect 2313 3331 2483 3503
rect 2695 3331 3063 3503
rect 3275 3331 3445 3503
rect 2313 3233 3445 3331
rect 2313 3061 2483 3233
rect 2695 3061 3063 3233
rect 3275 3061 3445 3233
rect 2313 2963 3445 3061
rect 2313 2791 2483 2963
rect 2695 2791 3063 2963
rect 3275 2791 3445 2963
rect 2313 2693 3445 2791
rect 2313 2521 2483 2693
rect 2695 2521 3063 2693
rect 3275 2521 3445 2693
rect 2313 2423 3445 2521
rect 2313 2251 2483 2423
rect 2695 2251 3063 2423
rect 3275 2251 3445 2423
rect 2313 2153 3445 2251
rect 2313 1981 2483 2153
rect 2695 1981 3063 2153
rect 3275 1981 3445 2153
rect 2313 1883 3445 1981
rect 2313 1711 2483 1883
rect 2695 1711 3063 1883
rect 3275 1711 3445 1883
rect 2313 1613 3445 1711
rect 2313 1441 2483 1613
rect 2695 1441 3063 1613
rect 3275 1441 3445 1613
rect 2313 1343 3445 1441
rect 2313 1171 2483 1343
rect 2695 1171 3063 1343
rect 3275 1171 3445 1343
rect 2313 1073 3445 1171
rect 2313 901 2483 1073
rect 2695 901 3063 1073
rect 3275 901 3445 1073
rect 2313 803 3445 901
rect 2313 631 2483 803
rect 2695 631 3063 803
rect 3275 631 3445 803
rect 2313 533 3445 631
rect 2313 361 2483 533
rect 2695 361 3063 533
rect 3275 361 3445 533
rect 2313 263 3445 361
rect 2313 91 2483 263
rect 2695 91 3063 263
rect 3275 91 3445 263
rect 2313 -7 3445 91
rect 3473 4141 3643 4313
rect 3855 4141 4223 4313
rect 4435 4141 4605 4313
rect 3473 4043 4605 4141
rect 3473 3871 3643 4043
rect 3855 3871 4223 4043
rect 4435 3871 4605 4043
rect 3473 3773 4605 3871
rect 3473 3601 3643 3773
rect 3855 3601 4223 3773
rect 4435 3601 4605 3773
rect 3473 3503 4605 3601
rect 3473 3331 3643 3503
rect 3855 3331 4223 3503
rect 4435 3331 4605 3503
rect 3473 3233 4605 3331
rect 3473 3061 3643 3233
rect 3855 3061 4223 3233
rect 4435 3061 4605 3233
rect 3473 2963 4605 3061
rect 3473 2791 3643 2963
rect 3855 2791 4223 2963
rect 4435 2791 4605 2963
rect 3473 2693 4605 2791
rect 3473 2521 3643 2693
rect 3855 2521 4223 2693
rect 4435 2521 4605 2693
rect 3473 2423 4605 2521
rect 3473 2251 3643 2423
rect 3855 2251 4223 2423
rect 4435 2251 4605 2423
rect 3473 2153 4605 2251
rect 3473 1981 3643 2153
rect 3855 1981 4223 2153
rect 4435 1981 4605 2153
rect 3473 1883 4605 1981
rect 3473 1711 3643 1883
rect 3855 1711 4223 1883
rect 4435 1711 4605 1883
rect 3473 1613 4605 1711
rect 3473 1441 3643 1613
rect 3855 1441 4223 1613
rect 4435 1441 4605 1613
rect 3473 1343 4605 1441
rect 3473 1171 3643 1343
rect 3855 1171 4223 1343
rect 4435 1171 4605 1343
rect 3473 1073 4605 1171
rect 3473 901 3643 1073
rect 3855 901 4223 1073
rect 4435 901 4605 1073
rect 3473 803 4605 901
rect 3473 631 3643 803
rect 3855 631 4223 803
rect 4435 631 4605 803
rect 3473 533 4605 631
rect 3473 361 3643 533
rect 3855 361 4223 533
rect 4435 361 4605 533
rect 3473 263 4605 361
rect 3473 91 3643 263
rect 3855 91 4223 263
rect 4435 91 4605 263
rect 3473 -7 4605 91
rect 4633 4141 4803 4313
rect 5015 4141 5383 4313
rect 5595 4141 5765 4313
rect 4633 4043 5765 4141
rect 4633 3871 4803 4043
rect 5015 3871 5383 4043
rect 5595 3871 5765 4043
rect 4633 3773 5765 3871
rect 4633 3601 4803 3773
rect 5015 3601 5383 3773
rect 5595 3601 5765 3773
rect 4633 3503 5765 3601
rect 4633 3331 4803 3503
rect 5015 3331 5383 3503
rect 5595 3331 5765 3503
rect 4633 3233 5765 3331
rect 4633 3061 4803 3233
rect 5015 3061 5383 3233
rect 5595 3061 5765 3233
rect 4633 2963 5765 3061
rect 4633 2791 4803 2963
rect 5015 2791 5383 2963
rect 5595 2791 5765 2963
rect 4633 2693 5765 2791
rect 4633 2521 4803 2693
rect 5015 2521 5383 2693
rect 5595 2521 5765 2693
rect 4633 2423 5765 2521
rect 4633 2251 4803 2423
rect 5015 2251 5383 2423
rect 5595 2251 5765 2423
rect 4633 2153 5765 2251
rect 4633 1981 4803 2153
rect 5015 1981 5383 2153
rect 5595 1981 5765 2153
rect 4633 1883 5765 1981
rect 4633 1711 4803 1883
rect 5015 1711 5383 1883
rect 5595 1711 5765 1883
rect 4633 1613 5765 1711
rect 4633 1441 4803 1613
rect 5015 1441 5383 1613
rect 5595 1441 5765 1613
rect 4633 1343 5765 1441
rect 4633 1171 4803 1343
rect 5015 1171 5383 1343
rect 5595 1171 5765 1343
rect 4633 1073 5765 1171
rect 4633 901 4803 1073
rect 5015 901 5383 1073
rect 5595 901 5765 1073
rect 4633 803 5765 901
rect 4633 631 4803 803
rect 5015 631 5383 803
rect 5595 631 5765 803
rect 4633 533 5765 631
rect 4633 361 4803 533
rect 5015 361 5383 533
rect 5595 361 5765 533
rect 4633 263 5765 361
rect 4633 91 4803 263
rect 5015 91 5383 263
rect 5595 91 5765 263
rect 4633 -7 5765 91
rect 5793 4141 5963 4313
rect 6175 4141 6543 4313
rect 6755 4141 6925 4313
rect 5793 4043 6925 4141
rect 5793 3871 5963 4043
rect 6175 3871 6543 4043
rect 6755 3871 6925 4043
rect 5793 3773 6925 3871
rect 5793 3601 5963 3773
rect 6175 3601 6543 3773
rect 6755 3601 6925 3773
rect 5793 3503 6925 3601
rect 5793 3331 5963 3503
rect 6175 3331 6543 3503
rect 6755 3331 6925 3503
rect 5793 3233 6925 3331
rect 5793 3061 5963 3233
rect 6175 3061 6543 3233
rect 6755 3061 6925 3233
rect 5793 2963 6925 3061
rect 5793 2791 5963 2963
rect 6175 2791 6543 2963
rect 6755 2791 6925 2963
rect 5793 2693 6925 2791
rect 5793 2521 5963 2693
rect 6175 2521 6543 2693
rect 6755 2521 6925 2693
rect 5793 2423 6925 2521
rect 5793 2251 5963 2423
rect 6175 2251 6543 2423
rect 6755 2251 6925 2423
rect 5793 2153 6925 2251
rect 5793 1981 5963 2153
rect 6175 1981 6543 2153
rect 6755 1981 6925 2153
rect 5793 1883 6925 1981
rect 5793 1711 5963 1883
rect 6175 1711 6543 1883
rect 6755 1711 6925 1883
rect 5793 1613 6925 1711
rect 5793 1441 5963 1613
rect 6175 1441 6543 1613
rect 6755 1441 6925 1613
rect 5793 1343 6925 1441
rect 5793 1171 5963 1343
rect 6175 1171 6543 1343
rect 6755 1171 6925 1343
rect 5793 1073 6925 1171
rect 5793 901 5963 1073
rect 6175 901 6543 1073
rect 6755 901 6925 1073
rect 5793 803 6925 901
rect 5793 631 5963 803
rect 6175 631 6543 803
rect 6755 631 6925 803
rect 5793 533 6925 631
rect 5793 361 5963 533
rect 6175 361 6543 533
rect 6755 361 6925 533
rect 5793 263 6925 361
rect 5793 91 5963 263
rect 6175 91 6543 263
rect 6755 91 6925 263
rect 5793 -7 6925 91
<< nmos >>
rect 100 4227 130 4255
rect 408 4227 438 4255
rect 680 4227 710 4255
rect 988 4227 1018 4255
rect 1260 4227 1290 4255
rect 1568 4227 1598 4255
rect 1840 4227 1870 4255
rect 2148 4227 2178 4255
rect 2420 4227 2450 4255
rect 2728 4227 2758 4255
rect 3000 4227 3030 4255
rect 3308 4227 3338 4255
rect 3580 4227 3610 4255
rect 3888 4227 3918 4255
rect 4160 4227 4190 4255
rect 4468 4227 4498 4255
rect 4740 4227 4770 4255
rect 5048 4227 5078 4255
rect 5320 4227 5350 4255
rect 5628 4227 5658 4255
rect 5900 4227 5930 4255
rect 6208 4227 6238 4255
rect 6480 4227 6510 4255
rect 6788 4227 6818 4255
rect 36 4081 66 4123
rect 472 4081 502 4123
rect 616 4081 646 4123
rect 1052 4081 1082 4123
rect 1196 4081 1226 4123
rect 1632 4081 1662 4123
rect 1776 4081 1806 4123
rect 2212 4081 2242 4123
rect 2356 4081 2386 4123
rect 2792 4081 2822 4123
rect 2936 4081 2966 4123
rect 3372 4081 3402 4123
rect 3516 4081 3546 4123
rect 3952 4081 3982 4123
rect 4096 4081 4126 4123
rect 4532 4081 4562 4123
rect 4676 4081 4706 4123
rect 5112 4081 5142 4123
rect 5256 4081 5286 4123
rect 5692 4081 5722 4123
rect 5836 4081 5866 4123
rect 6272 4081 6302 4123
rect 6416 4081 6446 4123
rect 6852 4081 6882 4123
rect 100 3957 130 3985
rect 408 3957 438 3985
rect 680 3957 710 3985
rect 988 3957 1018 3985
rect 1260 3957 1290 3985
rect 1568 3957 1598 3985
rect 1840 3957 1870 3985
rect 2148 3957 2178 3985
rect 2420 3957 2450 3985
rect 2728 3957 2758 3985
rect 3000 3957 3030 3985
rect 3308 3957 3338 3985
rect 3580 3957 3610 3985
rect 3888 3957 3918 3985
rect 4160 3957 4190 3985
rect 4468 3957 4498 3985
rect 4740 3957 4770 3985
rect 5048 3957 5078 3985
rect 5320 3957 5350 3985
rect 5628 3957 5658 3985
rect 5900 3957 5930 3985
rect 6208 3957 6238 3985
rect 6480 3957 6510 3985
rect 6788 3957 6818 3985
rect 36 3811 66 3853
rect 472 3811 502 3853
rect 616 3811 646 3853
rect 1052 3811 1082 3853
rect 1196 3811 1226 3853
rect 1632 3811 1662 3853
rect 1776 3811 1806 3853
rect 2212 3811 2242 3853
rect 2356 3811 2386 3853
rect 2792 3811 2822 3853
rect 2936 3811 2966 3853
rect 3372 3811 3402 3853
rect 3516 3811 3546 3853
rect 3952 3811 3982 3853
rect 4096 3811 4126 3853
rect 4532 3811 4562 3853
rect 4676 3811 4706 3853
rect 5112 3811 5142 3853
rect 5256 3811 5286 3853
rect 5692 3811 5722 3853
rect 5836 3811 5866 3853
rect 6272 3811 6302 3853
rect 6416 3811 6446 3853
rect 6852 3811 6882 3853
rect 100 3687 130 3715
rect 408 3687 438 3715
rect 680 3687 710 3715
rect 988 3687 1018 3715
rect 1260 3687 1290 3715
rect 1568 3687 1598 3715
rect 1840 3687 1870 3715
rect 2148 3687 2178 3715
rect 2420 3687 2450 3715
rect 2728 3687 2758 3715
rect 3000 3687 3030 3715
rect 3308 3687 3338 3715
rect 3580 3687 3610 3715
rect 3888 3687 3918 3715
rect 4160 3687 4190 3715
rect 4468 3687 4498 3715
rect 4740 3687 4770 3715
rect 5048 3687 5078 3715
rect 5320 3687 5350 3715
rect 5628 3687 5658 3715
rect 5900 3687 5930 3715
rect 6208 3687 6238 3715
rect 6480 3687 6510 3715
rect 6788 3687 6818 3715
rect 36 3541 66 3583
rect 472 3541 502 3583
rect 616 3541 646 3583
rect 1052 3541 1082 3583
rect 1196 3541 1226 3583
rect 1632 3541 1662 3583
rect 1776 3541 1806 3583
rect 2212 3541 2242 3583
rect 2356 3541 2386 3583
rect 2792 3541 2822 3583
rect 2936 3541 2966 3583
rect 3372 3541 3402 3583
rect 3516 3541 3546 3583
rect 3952 3541 3982 3583
rect 4096 3541 4126 3583
rect 4532 3541 4562 3583
rect 4676 3541 4706 3583
rect 5112 3541 5142 3583
rect 5256 3541 5286 3583
rect 5692 3541 5722 3583
rect 5836 3541 5866 3583
rect 6272 3541 6302 3583
rect 6416 3541 6446 3583
rect 6852 3541 6882 3583
rect 100 3417 130 3445
rect 408 3417 438 3445
rect 680 3417 710 3445
rect 988 3417 1018 3445
rect 1260 3417 1290 3445
rect 1568 3417 1598 3445
rect 1840 3417 1870 3445
rect 2148 3417 2178 3445
rect 2420 3417 2450 3445
rect 2728 3417 2758 3445
rect 3000 3417 3030 3445
rect 3308 3417 3338 3445
rect 3580 3417 3610 3445
rect 3888 3417 3918 3445
rect 4160 3417 4190 3445
rect 4468 3417 4498 3445
rect 4740 3417 4770 3445
rect 5048 3417 5078 3445
rect 5320 3417 5350 3445
rect 5628 3417 5658 3445
rect 5900 3417 5930 3445
rect 6208 3417 6238 3445
rect 6480 3417 6510 3445
rect 6788 3417 6818 3445
rect 36 3271 66 3313
rect 472 3271 502 3313
rect 616 3271 646 3313
rect 1052 3271 1082 3313
rect 1196 3271 1226 3313
rect 1632 3271 1662 3313
rect 1776 3271 1806 3313
rect 2212 3271 2242 3313
rect 2356 3271 2386 3313
rect 2792 3271 2822 3313
rect 2936 3271 2966 3313
rect 3372 3271 3402 3313
rect 3516 3271 3546 3313
rect 3952 3271 3982 3313
rect 4096 3271 4126 3313
rect 4532 3271 4562 3313
rect 4676 3271 4706 3313
rect 5112 3271 5142 3313
rect 5256 3271 5286 3313
rect 5692 3271 5722 3313
rect 5836 3271 5866 3313
rect 6272 3271 6302 3313
rect 6416 3271 6446 3313
rect 6852 3271 6882 3313
rect 100 3147 130 3175
rect 408 3147 438 3175
rect 680 3147 710 3175
rect 988 3147 1018 3175
rect 1260 3147 1290 3175
rect 1568 3147 1598 3175
rect 1840 3147 1870 3175
rect 2148 3147 2178 3175
rect 2420 3147 2450 3175
rect 2728 3147 2758 3175
rect 3000 3147 3030 3175
rect 3308 3147 3338 3175
rect 3580 3147 3610 3175
rect 3888 3147 3918 3175
rect 4160 3147 4190 3175
rect 4468 3147 4498 3175
rect 4740 3147 4770 3175
rect 5048 3147 5078 3175
rect 5320 3147 5350 3175
rect 5628 3147 5658 3175
rect 5900 3147 5930 3175
rect 6208 3147 6238 3175
rect 6480 3147 6510 3175
rect 6788 3147 6818 3175
rect 36 3001 66 3043
rect 472 3001 502 3043
rect 616 3001 646 3043
rect 1052 3001 1082 3043
rect 1196 3001 1226 3043
rect 1632 3001 1662 3043
rect 1776 3001 1806 3043
rect 2212 3001 2242 3043
rect 2356 3001 2386 3043
rect 2792 3001 2822 3043
rect 2936 3001 2966 3043
rect 3372 3001 3402 3043
rect 3516 3001 3546 3043
rect 3952 3001 3982 3043
rect 4096 3001 4126 3043
rect 4532 3001 4562 3043
rect 4676 3001 4706 3043
rect 5112 3001 5142 3043
rect 5256 3001 5286 3043
rect 5692 3001 5722 3043
rect 5836 3001 5866 3043
rect 6272 3001 6302 3043
rect 6416 3001 6446 3043
rect 6852 3001 6882 3043
rect 100 2877 130 2905
rect 408 2877 438 2905
rect 680 2877 710 2905
rect 988 2877 1018 2905
rect 1260 2877 1290 2905
rect 1568 2877 1598 2905
rect 1840 2877 1870 2905
rect 2148 2877 2178 2905
rect 2420 2877 2450 2905
rect 2728 2877 2758 2905
rect 3000 2877 3030 2905
rect 3308 2877 3338 2905
rect 3580 2877 3610 2905
rect 3888 2877 3918 2905
rect 4160 2877 4190 2905
rect 4468 2877 4498 2905
rect 4740 2877 4770 2905
rect 5048 2877 5078 2905
rect 5320 2877 5350 2905
rect 5628 2877 5658 2905
rect 5900 2877 5930 2905
rect 6208 2877 6238 2905
rect 6480 2877 6510 2905
rect 6788 2877 6818 2905
rect 36 2731 66 2773
rect 472 2731 502 2773
rect 616 2731 646 2773
rect 1052 2731 1082 2773
rect 1196 2731 1226 2773
rect 1632 2731 1662 2773
rect 1776 2731 1806 2773
rect 2212 2731 2242 2773
rect 2356 2731 2386 2773
rect 2792 2731 2822 2773
rect 2936 2731 2966 2773
rect 3372 2731 3402 2773
rect 3516 2731 3546 2773
rect 3952 2731 3982 2773
rect 4096 2731 4126 2773
rect 4532 2731 4562 2773
rect 4676 2731 4706 2773
rect 5112 2731 5142 2773
rect 5256 2731 5286 2773
rect 5692 2731 5722 2773
rect 5836 2731 5866 2773
rect 6272 2731 6302 2773
rect 6416 2731 6446 2773
rect 6852 2731 6882 2773
rect 100 2607 130 2635
rect 408 2607 438 2635
rect 680 2607 710 2635
rect 988 2607 1018 2635
rect 1260 2607 1290 2635
rect 1568 2607 1598 2635
rect 1840 2607 1870 2635
rect 2148 2607 2178 2635
rect 2420 2607 2450 2635
rect 2728 2607 2758 2635
rect 3000 2607 3030 2635
rect 3308 2607 3338 2635
rect 3580 2607 3610 2635
rect 3888 2607 3918 2635
rect 4160 2607 4190 2635
rect 4468 2607 4498 2635
rect 4740 2607 4770 2635
rect 5048 2607 5078 2635
rect 5320 2607 5350 2635
rect 5628 2607 5658 2635
rect 5900 2607 5930 2635
rect 6208 2607 6238 2635
rect 6480 2607 6510 2635
rect 6788 2607 6818 2635
rect 36 2461 66 2503
rect 472 2461 502 2503
rect 616 2461 646 2503
rect 1052 2461 1082 2503
rect 1196 2461 1226 2503
rect 1632 2461 1662 2503
rect 1776 2461 1806 2503
rect 2212 2461 2242 2503
rect 2356 2461 2386 2503
rect 2792 2461 2822 2503
rect 2936 2461 2966 2503
rect 3372 2461 3402 2503
rect 3516 2461 3546 2503
rect 3952 2461 3982 2503
rect 4096 2461 4126 2503
rect 4532 2461 4562 2503
rect 4676 2461 4706 2503
rect 5112 2461 5142 2503
rect 5256 2461 5286 2503
rect 5692 2461 5722 2503
rect 5836 2461 5866 2503
rect 6272 2461 6302 2503
rect 6416 2461 6446 2503
rect 6852 2461 6882 2503
rect 100 2337 130 2365
rect 408 2337 438 2365
rect 680 2337 710 2365
rect 988 2337 1018 2365
rect 1260 2337 1290 2365
rect 1568 2337 1598 2365
rect 1840 2337 1870 2365
rect 2148 2337 2178 2365
rect 2420 2337 2450 2365
rect 2728 2337 2758 2365
rect 3000 2337 3030 2365
rect 3308 2337 3338 2365
rect 3580 2337 3610 2365
rect 3888 2337 3918 2365
rect 4160 2337 4190 2365
rect 4468 2337 4498 2365
rect 4740 2337 4770 2365
rect 5048 2337 5078 2365
rect 5320 2337 5350 2365
rect 5628 2337 5658 2365
rect 5900 2337 5930 2365
rect 6208 2337 6238 2365
rect 6480 2337 6510 2365
rect 6788 2337 6818 2365
rect 36 2191 66 2233
rect 472 2191 502 2233
rect 616 2191 646 2233
rect 1052 2191 1082 2233
rect 1196 2191 1226 2233
rect 1632 2191 1662 2233
rect 1776 2191 1806 2233
rect 2212 2191 2242 2233
rect 2356 2191 2386 2233
rect 2792 2191 2822 2233
rect 2936 2191 2966 2233
rect 3372 2191 3402 2233
rect 3516 2191 3546 2233
rect 3952 2191 3982 2233
rect 4096 2191 4126 2233
rect 4532 2191 4562 2233
rect 4676 2191 4706 2233
rect 5112 2191 5142 2233
rect 5256 2191 5286 2233
rect 5692 2191 5722 2233
rect 5836 2191 5866 2233
rect 6272 2191 6302 2233
rect 6416 2191 6446 2233
rect 6852 2191 6882 2233
rect 100 2067 130 2095
rect 408 2067 438 2095
rect 680 2067 710 2095
rect 988 2067 1018 2095
rect 1260 2067 1290 2095
rect 1568 2067 1598 2095
rect 1840 2067 1870 2095
rect 2148 2067 2178 2095
rect 2420 2067 2450 2095
rect 2728 2067 2758 2095
rect 3000 2067 3030 2095
rect 3308 2067 3338 2095
rect 3580 2067 3610 2095
rect 3888 2067 3918 2095
rect 4160 2067 4190 2095
rect 4468 2067 4498 2095
rect 4740 2067 4770 2095
rect 5048 2067 5078 2095
rect 5320 2067 5350 2095
rect 5628 2067 5658 2095
rect 5900 2067 5930 2095
rect 6208 2067 6238 2095
rect 6480 2067 6510 2095
rect 6788 2067 6818 2095
rect 36 1921 66 1963
rect 472 1921 502 1963
rect 616 1921 646 1963
rect 1052 1921 1082 1963
rect 1196 1921 1226 1963
rect 1632 1921 1662 1963
rect 1776 1921 1806 1963
rect 2212 1921 2242 1963
rect 2356 1921 2386 1963
rect 2792 1921 2822 1963
rect 2936 1921 2966 1963
rect 3372 1921 3402 1963
rect 3516 1921 3546 1963
rect 3952 1921 3982 1963
rect 4096 1921 4126 1963
rect 4532 1921 4562 1963
rect 4676 1921 4706 1963
rect 5112 1921 5142 1963
rect 5256 1921 5286 1963
rect 5692 1921 5722 1963
rect 5836 1921 5866 1963
rect 6272 1921 6302 1963
rect 6416 1921 6446 1963
rect 6852 1921 6882 1963
rect 100 1797 130 1825
rect 408 1797 438 1825
rect 680 1797 710 1825
rect 988 1797 1018 1825
rect 1260 1797 1290 1825
rect 1568 1797 1598 1825
rect 1840 1797 1870 1825
rect 2148 1797 2178 1825
rect 2420 1797 2450 1825
rect 2728 1797 2758 1825
rect 3000 1797 3030 1825
rect 3308 1797 3338 1825
rect 3580 1797 3610 1825
rect 3888 1797 3918 1825
rect 4160 1797 4190 1825
rect 4468 1797 4498 1825
rect 4740 1797 4770 1825
rect 5048 1797 5078 1825
rect 5320 1797 5350 1825
rect 5628 1797 5658 1825
rect 5900 1797 5930 1825
rect 6208 1797 6238 1825
rect 6480 1797 6510 1825
rect 6788 1797 6818 1825
rect 36 1651 66 1693
rect 472 1651 502 1693
rect 616 1651 646 1693
rect 1052 1651 1082 1693
rect 1196 1651 1226 1693
rect 1632 1651 1662 1693
rect 1776 1651 1806 1693
rect 2212 1651 2242 1693
rect 2356 1651 2386 1693
rect 2792 1651 2822 1693
rect 2936 1651 2966 1693
rect 3372 1651 3402 1693
rect 3516 1651 3546 1693
rect 3952 1651 3982 1693
rect 4096 1651 4126 1693
rect 4532 1651 4562 1693
rect 4676 1651 4706 1693
rect 5112 1651 5142 1693
rect 5256 1651 5286 1693
rect 5692 1651 5722 1693
rect 5836 1651 5866 1693
rect 6272 1651 6302 1693
rect 6416 1651 6446 1693
rect 6852 1651 6882 1693
rect 100 1527 130 1555
rect 408 1527 438 1555
rect 680 1527 710 1555
rect 988 1527 1018 1555
rect 1260 1527 1290 1555
rect 1568 1527 1598 1555
rect 1840 1527 1870 1555
rect 2148 1527 2178 1555
rect 2420 1527 2450 1555
rect 2728 1527 2758 1555
rect 3000 1527 3030 1555
rect 3308 1527 3338 1555
rect 3580 1527 3610 1555
rect 3888 1527 3918 1555
rect 4160 1527 4190 1555
rect 4468 1527 4498 1555
rect 4740 1527 4770 1555
rect 5048 1527 5078 1555
rect 5320 1527 5350 1555
rect 5628 1527 5658 1555
rect 5900 1527 5930 1555
rect 6208 1527 6238 1555
rect 6480 1527 6510 1555
rect 6788 1527 6818 1555
rect 36 1381 66 1423
rect 472 1381 502 1423
rect 616 1381 646 1423
rect 1052 1381 1082 1423
rect 1196 1381 1226 1423
rect 1632 1381 1662 1423
rect 1776 1381 1806 1423
rect 2212 1381 2242 1423
rect 2356 1381 2386 1423
rect 2792 1381 2822 1423
rect 2936 1381 2966 1423
rect 3372 1381 3402 1423
rect 3516 1381 3546 1423
rect 3952 1381 3982 1423
rect 4096 1381 4126 1423
rect 4532 1381 4562 1423
rect 4676 1381 4706 1423
rect 5112 1381 5142 1423
rect 5256 1381 5286 1423
rect 5692 1381 5722 1423
rect 5836 1381 5866 1423
rect 6272 1381 6302 1423
rect 6416 1381 6446 1423
rect 6852 1381 6882 1423
rect 100 1257 130 1285
rect 408 1257 438 1285
rect 680 1257 710 1285
rect 988 1257 1018 1285
rect 1260 1257 1290 1285
rect 1568 1257 1598 1285
rect 1840 1257 1870 1285
rect 2148 1257 2178 1285
rect 2420 1257 2450 1285
rect 2728 1257 2758 1285
rect 3000 1257 3030 1285
rect 3308 1257 3338 1285
rect 3580 1257 3610 1285
rect 3888 1257 3918 1285
rect 4160 1257 4190 1285
rect 4468 1257 4498 1285
rect 4740 1257 4770 1285
rect 5048 1257 5078 1285
rect 5320 1257 5350 1285
rect 5628 1257 5658 1285
rect 5900 1257 5930 1285
rect 6208 1257 6238 1285
rect 6480 1257 6510 1285
rect 6788 1257 6818 1285
rect 36 1111 66 1153
rect 472 1111 502 1153
rect 616 1111 646 1153
rect 1052 1111 1082 1153
rect 1196 1111 1226 1153
rect 1632 1111 1662 1153
rect 1776 1111 1806 1153
rect 2212 1111 2242 1153
rect 2356 1111 2386 1153
rect 2792 1111 2822 1153
rect 2936 1111 2966 1153
rect 3372 1111 3402 1153
rect 3516 1111 3546 1153
rect 3952 1111 3982 1153
rect 4096 1111 4126 1153
rect 4532 1111 4562 1153
rect 4676 1111 4706 1153
rect 5112 1111 5142 1153
rect 5256 1111 5286 1153
rect 5692 1111 5722 1153
rect 5836 1111 5866 1153
rect 6272 1111 6302 1153
rect 6416 1111 6446 1153
rect 6852 1111 6882 1153
rect 100 987 130 1015
rect 408 987 438 1015
rect 680 987 710 1015
rect 988 987 1018 1015
rect 1260 987 1290 1015
rect 1568 987 1598 1015
rect 1840 987 1870 1015
rect 2148 987 2178 1015
rect 2420 987 2450 1015
rect 2728 987 2758 1015
rect 3000 987 3030 1015
rect 3308 987 3338 1015
rect 3580 987 3610 1015
rect 3888 987 3918 1015
rect 4160 987 4190 1015
rect 4468 987 4498 1015
rect 4740 987 4770 1015
rect 5048 987 5078 1015
rect 5320 987 5350 1015
rect 5628 987 5658 1015
rect 5900 987 5930 1015
rect 6208 987 6238 1015
rect 6480 987 6510 1015
rect 6788 987 6818 1015
rect 36 841 66 883
rect 472 841 502 883
rect 616 841 646 883
rect 1052 841 1082 883
rect 1196 841 1226 883
rect 1632 841 1662 883
rect 1776 841 1806 883
rect 2212 841 2242 883
rect 2356 841 2386 883
rect 2792 841 2822 883
rect 2936 841 2966 883
rect 3372 841 3402 883
rect 3516 841 3546 883
rect 3952 841 3982 883
rect 4096 841 4126 883
rect 4532 841 4562 883
rect 4676 841 4706 883
rect 5112 841 5142 883
rect 5256 841 5286 883
rect 5692 841 5722 883
rect 5836 841 5866 883
rect 6272 841 6302 883
rect 6416 841 6446 883
rect 6852 841 6882 883
rect 100 717 130 745
rect 408 717 438 745
rect 680 717 710 745
rect 988 717 1018 745
rect 1260 717 1290 745
rect 1568 717 1598 745
rect 1840 717 1870 745
rect 2148 717 2178 745
rect 2420 717 2450 745
rect 2728 717 2758 745
rect 3000 717 3030 745
rect 3308 717 3338 745
rect 3580 717 3610 745
rect 3888 717 3918 745
rect 4160 717 4190 745
rect 4468 717 4498 745
rect 4740 717 4770 745
rect 5048 717 5078 745
rect 5320 717 5350 745
rect 5628 717 5658 745
rect 5900 717 5930 745
rect 6208 717 6238 745
rect 6480 717 6510 745
rect 6788 717 6818 745
rect 36 571 66 613
rect 472 571 502 613
rect 616 571 646 613
rect 1052 571 1082 613
rect 1196 571 1226 613
rect 1632 571 1662 613
rect 1776 571 1806 613
rect 2212 571 2242 613
rect 2356 571 2386 613
rect 2792 571 2822 613
rect 2936 571 2966 613
rect 3372 571 3402 613
rect 3516 571 3546 613
rect 3952 571 3982 613
rect 4096 571 4126 613
rect 4532 571 4562 613
rect 4676 571 4706 613
rect 5112 571 5142 613
rect 5256 571 5286 613
rect 5692 571 5722 613
rect 5836 571 5866 613
rect 6272 571 6302 613
rect 6416 571 6446 613
rect 6852 571 6882 613
rect 100 447 130 475
rect 408 447 438 475
rect 680 447 710 475
rect 988 447 1018 475
rect 1260 447 1290 475
rect 1568 447 1598 475
rect 1840 447 1870 475
rect 2148 447 2178 475
rect 2420 447 2450 475
rect 2728 447 2758 475
rect 3000 447 3030 475
rect 3308 447 3338 475
rect 3580 447 3610 475
rect 3888 447 3918 475
rect 4160 447 4190 475
rect 4468 447 4498 475
rect 4740 447 4770 475
rect 5048 447 5078 475
rect 5320 447 5350 475
rect 5628 447 5658 475
rect 5900 447 5930 475
rect 6208 447 6238 475
rect 6480 447 6510 475
rect 6788 447 6818 475
rect 36 301 66 343
rect 472 301 502 343
rect 616 301 646 343
rect 1052 301 1082 343
rect 1196 301 1226 343
rect 1632 301 1662 343
rect 1776 301 1806 343
rect 2212 301 2242 343
rect 2356 301 2386 343
rect 2792 301 2822 343
rect 2936 301 2966 343
rect 3372 301 3402 343
rect 3516 301 3546 343
rect 3952 301 3982 343
rect 4096 301 4126 343
rect 4532 301 4562 343
rect 4676 301 4706 343
rect 5112 301 5142 343
rect 5256 301 5286 343
rect 5692 301 5722 343
rect 5836 301 5866 343
rect 6272 301 6302 343
rect 6416 301 6446 343
rect 6852 301 6882 343
rect 100 177 130 205
rect 408 177 438 205
rect 680 177 710 205
rect 988 177 1018 205
rect 1260 177 1290 205
rect 1568 177 1598 205
rect 1840 177 1870 205
rect 2148 177 2178 205
rect 2420 177 2450 205
rect 2728 177 2758 205
rect 3000 177 3030 205
rect 3308 177 3338 205
rect 3580 177 3610 205
rect 3888 177 3918 205
rect 4160 177 4190 205
rect 4468 177 4498 205
rect 4740 177 4770 205
rect 5048 177 5078 205
rect 5320 177 5350 205
rect 5628 177 5658 205
rect 5900 177 5930 205
rect 6208 177 6238 205
rect 6480 177 6510 205
rect 6788 177 6818 205
rect 36 31 66 73
rect 472 31 502 73
rect 616 31 646 73
rect 1052 31 1082 73
rect 1196 31 1226 73
rect 1632 31 1662 73
rect 1776 31 1806 73
rect 2212 31 2242 73
rect 2356 31 2386 73
rect 2792 31 2822 73
rect 2936 31 2966 73
rect 3372 31 3402 73
rect 3516 31 3546 73
rect 3952 31 3982 73
rect 4096 31 4126 73
rect 4532 31 4562 73
rect 4676 31 4706 73
rect 5112 31 5142 73
rect 5256 31 5286 73
rect 5692 31 5722 73
rect 5836 31 5866 73
rect 6272 31 6302 73
rect 6416 31 6446 73
rect 6852 31 6882 73
<< npd >>
rect 215 4081 245 4123
rect 293 4081 323 4123
rect 795 4081 825 4123
rect 873 4081 903 4123
rect 1375 4081 1405 4123
rect 1453 4081 1483 4123
rect 1955 4081 1985 4123
rect 2033 4081 2063 4123
rect 2535 4081 2565 4123
rect 2613 4081 2643 4123
rect 3115 4081 3145 4123
rect 3193 4081 3223 4123
rect 3695 4081 3725 4123
rect 3773 4081 3803 4123
rect 4275 4081 4305 4123
rect 4353 4081 4383 4123
rect 4855 4081 4885 4123
rect 4933 4081 4963 4123
rect 5435 4081 5465 4123
rect 5513 4081 5543 4123
rect 6015 4081 6045 4123
rect 6093 4081 6123 4123
rect 6595 4081 6625 4123
rect 6673 4081 6703 4123
rect 215 3811 245 3853
rect 293 3811 323 3853
rect 795 3811 825 3853
rect 873 3811 903 3853
rect 1375 3811 1405 3853
rect 1453 3811 1483 3853
rect 1955 3811 1985 3853
rect 2033 3811 2063 3853
rect 2535 3811 2565 3853
rect 2613 3811 2643 3853
rect 3115 3811 3145 3853
rect 3193 3811 3223 3853
rect 3695 3811 3725 3853
rect 3773 3811 3803 3853
rect 4275 3811 4305 3853
rect 4353 3811 4383 3853
rect 4855 3811 4885 3853
rect 4933 3811 4963 3853
rect 5435 3811 5465 3853
rect 5513 3811 5543 3853
rect 6015 3811 6045 3853
rect 6093 3811 6123 3853
rect 6595 3811 6625 3853
rect 6673 3811 6703 3853
rect 215 3541 245 3583
rect 293 3541 323 3583
rect 795 3541 825 3583
rect 873 3541 903 3583
rect 1375 3541 1405 3583
rect 1453 3541 1483 3583
rect 1955 3541 1985 3583
rect 2033 3541 2063 3583
rect 2535 3541 2565 3583
rect 2613 3541 2643 3583
rect 3115 3541 3145 3583
rect 3193 3541 3223 3583
rect 3695 3541 3725 3583
rect 3773 3541 3803 3583
rect 4275 3541 4305 3583
rect 4353 3541 4383 3583
rect 4855 3541 4885 3583
rect 4933 3541 4963 3583
rect 5435 3541 5465 3583
rect 5513 3541 5543 3583
rect 6015 3541 6045 3583
rect 6093 3541 6123 3583
rect 6595 3541 6625 3583
rect 6673 3541 6703 3583
rect 215 3271 245 3313
rect 293 3271 323 3313
rect 795 3271 825 3313
rect 873 3271 903 3313
rect 1375 3271 1405 3313
rect 1453 3271 1483 3313
rect 1955 3271 1985 3313
rect 2033 3271 2063 3313
rect 2535 3271 2565 3313
rect 2613 3271 2643 3313
rect 3115 3271 3145 3313
rect 3193 3271 3223 3313
rect 3695 3271 3725 3313
rect 3773 3271 3803 3313
rect 4275 3271 4305 3313
rect 4353 3271 4383 3313
rect 4855 3271 4885 3313
rect 4933 3271 4963 3313
rect 5435 3271 5465 3313
rect 5513 3271 5543 3313
rect 6015 3271 6045 3313
rect 6093 3271 6123 3313
rect 6595 3271 6625 3313
rect 6673 3271 6703 3313
rect 215 3001 245 3043
rect 293 3001 323 3043
rect 795 3001 825 3043
rect 873 3001 903 3043
rect 1375 3001 1405 3043
rect 1453 3001 1483 3043
rect 1955 3001 1985 3043
rect 2033 3001 2063 3043
rect 2535 3001 2565 3043
rect 2613 3001 2643 3043
rect 3115 3001 3145 3043
rect 3193 3001 3223 3043
rect 3695 3001 3725 3043
rect 3773 3001 3803 3043
rect 4275 3001 4305 3043
rect 4353 3001 4383 3043
rect 4855 3001 4885 3043
rect 4933 3001 4963 3043
rect 5435 3001 5465 3043
rect 5513 3001 5543 3043
rect 6015 3001 6045 3043
rect 6093 3001 6123 3043
rect 6595 3001 6625 3043
rect 6673 3001 6703 3043
rect 215 2731 245 2773
rect 293 2731 323 2773
rect 795 2731 825 2773
rect 873 2731 903 2773
rect 1375 2731 1405 2773
rect 1453 2731 1483 2773
rect 1955 2731 1985 2773
rect 2033 2731 2063 2773
rect 2535 2731 2565 2773
rect 2613 2731 2643 2773
rect 3115 2731 3145 2773
rect 3193 2731 3223 2773
rect 3695 2731 3725 2773
rect 3773 2731 3803 2773
rect 4275 2731 4305 2773
rect 4353 2731 4383 2773
rect 4855 2731 4885 2773
rect 4933 2731 4963 2773
rect 5435 2731 5465 2773
rect 5513 2731 5543 2773
rect 6015 2731 6045 2773
rect 6093 2731 6123 2773
rect 6595 2731 6625 2773
rect 6673 2731 6703 2773
rect 215 2461 245 2503
rect 293 2461 323 2503
rect 795 2461 825 2503
rect 873 2461 903 2503
rect 1375 2461 1405 2503
rect 1453 2461 1483 2503
rect 1955 2461 1985 2503
rect 2033 2461 2063 2503
rect 2535 2461 2565 2503
rect 2613 2461 2643 2503
rect 3115 2461 3145 2503
rect 3193 2461 3223 2503
rect 3695 2461 3725 2503
rect 3773 2461 3803 2503
rect 4275 2461 4305 2503
rect 4353 2461 4383 2503
rect 4855 2461 4885 2503
rect 4933 2461 4963 2503
rect 5435 2461 5465 2503
rect 5513 2461 5543 2503
rect 6015 2461 6045 2503
rect 6093 2461 6123 2503
rect 6595 2461 6625 2503
rect 6673 2461 6703 2503
rect 215 2191 245 2233
rect 293 2191 323 2233
rect 795 2191 825 2233
rect 873 2191 903 2233
rect 1375 2191 1405 2233
rect 1453 2191 1483 2233
rect 1955 2191 1985 2233
rect 2033 2191 2063 2233
rect 2535 2191 2565 2233
rect 2613 2191 2643 2233
rect 3115 2191 3145 2233
rect 3193 2191 3223 2233
rect 3695 2191 3725 2233
rect 3773 2191 3803 2233
rect 4275 2191 4305 2233
rect 4353 2191 4383 2233
rect 4855 2191 4885 2233
rect 4933 2191 4963 2233
rect 5435 2191 5465 2233
rect 5513 2191 5543 2233
rect 6015 2191 6045 2233
rect 6093 2191 6123 2233
rect 6595 2191 6625 2233
rect 6673 2191 6703 2233
rect 215 1921 245 1963
rect 293 1921 323 1963
rect 795 1921 825 1963
rect 873 1921 903 1963
rect 1375 1921 1405 1963
rect 1453 1921 1483 1963
rect 1955 1921 1985 1963
rect 2033 1921 2063 1963
rect 2535 1921 2565 1963
rect 2613 1921 2643 1963
rect 3115 1921 3145 1963
rect 3193 1921 3223 1963
rect 3695 1921 3725 1963
rect 3773 1921 3803 1963
rect 4275 1921 4305 1963
rect 4353 1921 4383 1963
rect 4855 1921 4885 1963
rect 4933 1921 4963 1963
rect 5435 1921 5465 1963
rect 5513 1921 5543 1963
rect 6015 1921 6045 1963
rect 6093 1921 6123 1963
rect 6595 1921 6625 1963
rect 6673 1921 6703 1963
rect 215 1651 245 1693
rect 293 1651 323 1693
rect 795 1651 825 1693
rect 873 1651 903 1693
rect 1375 1651 1405 1693
rect 1453 1651 1483 1693
rect 1955 1651 1985 1693
rect 2033 1651 2063 1693
rect 2535 1651 2565 1693
rect 2613 1651 2643 1693
rect 3115 1651 3145 1693
rect 3193 1651 3223 1693
rect 3695 1651 3725 1693
rect 3773 1651 3803 1693
rect 4275 1651 4305 1693
rect 4353 1651 4383 1693
rect 4855 1651 4885 1693
rect 4933 1651 4963 1693
rect 5435 1651 5465 1693
rect 5513 1651 5543 1693
rect 6015 1651 6045 1693
rect 6093 1651 6123 1693
rect 6595 1651 6625 1693
rect 6673 1651 6703 1693
rect 215 1381 245 1423
rect 293 1381 323 1423
rect 795 1381 825 1423
rect 873 1381 903 1423
rect 1375 1381 1405 1423
rect 1453 1381 1483 1423
rect 1955 1381 1985 1423
rect 2033 1381 2063 1423
rect 2535 1381 2565 1423
rect 2613 1381 2643 1423
rect 3115 1381 3145 1423
rect 3193 1381 3223 1423
rect 3695 1381 3725 1423
rect 3773 1381 3803 1423
rect 4275 1381 4305 1423
rect 4353 1381 4383 1423
rect 4855 1381 4885 1423
rect 4933 1381 4963 1423
rect 5435 1381 5465 1423
rect 5513 1381 5543 1423
rect 6015 1381 6045 1423
rect 6093 1381 6123 1423
rect 6595 1381 6625 1423
rect 6673 1381 6703 1423
rect 215 1111 245 1153
rect 293 1111 323 1153
rect 795 1111 825 1153
rect 873 1111 903 1153
rect 1375 1111 1405 1153
rect 1453 1111 1483 1153
rect 1955 1111 1985 1153
rect 2033 1111 2063 1153
rect 2535 1111 2565 1153
rect 2613 1111 2643 1153
rect 3115 1111 3145 1153
rect 3193 1111 3223 1153
rect 3695 1111 3725 1153
rect 3773 1111 3803 1153
rect 4275 1111 4305 1153
rect 4353 1111 4383 1153
rect 4855 1111 4885 1153
rect 4933 1111 4963 1153
rect 5435 1111 5465 1153
rect 5513 1111 5543 1153
rect 6015 1111 6045 1153
rect 6093 1111 6123 1153
rect 6595 1111 6625 1153
rect 6673 1111 6703 1153
rect 215 841 245 883
rect 293 841 323 883
rect 795 841 825 883
rect 873 841 903 883
rect 1375 841 1405 883
rect 1453 841 1483 883
rect 1955 841 1985 883
rect 2033 841 2063 883
rect 2535 841 2565 883
rect 2613 841 2643 883
rect 3115 841 3145 883
rect 3193 841 3223 883
rect 3695 841 3725 883
rect 3773 841 3803 883
rect 4275 841 4305 883
rect 4353 841 4383 883
rect 4855 841 4885 883
rect 4933 841 4963 883
rect 5435 841 5465 883
rect 5513 841 5543 883
rect 6015 841 6045 883
rect 6093 841 6123 883
rect 6595 841 6625 883
rect 6673 841 6703 883
rect 215 571 245 613
rect 293 571 323 613
rect 795 571 825 613
rect 873 571 903 613
rect 1375 571 1405 613
rect 1453 571 1483 613
rect 1955 571 1985 613
rect 2033 571 2063 613
rect 2535 571 2565 613
rect 2613 571 2643 613
rect 3115 571 3145 613
rect 3193 571 3223 613
rect 3695 571 3725 613
rect 3773 571 3803 613
rect 4275 571 4305 613
rect 4353 571 4383 613
rect 4855 571 4885 613
rect 4933 571 4963 613
rect 5435 571 5465 613
rect 5513 571 5543 613
rect 6015 571 6045 613
rect 6093 571 6123 613
rect 6595 571 6625 613
rect 6673 571 6703 613
rect 215 301 245 343
rect 293 301 323 343
rect 795 301 825 343
rect 873 301 903 343
rect 1375 301 1405 343
rect 1453 301 1483 343
rect 1955 301 1985 343
rect 2033 301 2063 343
rect 2535 301 2565 343
rect 2613 301 2643 343
rect 3115 301 3145 343
rect 3193 301 3223 343
rect 3695 301 3725 343
rect 3773 301 3803 343
rect 4275 301 4305 343
rect 4353 301 4383 343
rect 4855 301 4885 343
rect 4933 301 4963 343
rect 5435 301 5465 343
rect 5513 301 5543 343
rect 6015 301 6045 343
rect 6093 301 6123 343
rect 6595 301 6625 343
rect 6673 301 6703 343
rect 215 31 245 73
rect 293 31 323 73
rect 795 31 825 73
rect 873 31 903 73
rect 1375 31 1405 73
rect 1453 31 1483 73
rect 1955 31 1985 73
rect 2033 31 2063 73
rect 2535 31 2565 73
rect 2613 31 2643 73
rect 3115 31 3145 73
rect 3193 31 3223 73
rect 3695 31 3725 73
rect 3773 31 3803 73
rect 4275 31 4305 73
rect 4353 31 4383 73
rect 4855 31 4885 73
rect 4933 31 4963 73
rect 5435 31 5465 73
rect 5513 31 5543 73
rect 6015 31 6045 73
rect 6093 31 6123 73
rect 6595 31 6625 73
rect 6673 31 6703 73
<< npass >>
rect 122 4081 152 4109
rect 386 4081 416 4109
rect 702 4081 732 4109
rect 966 4081 996 4109
rect 1282 4081 1312 4109
rect 1546 4081 1576 4109
rect 1862 4081 1892 4109
rect 2126 4081 2156 4109
rect 2442 4081 2472 4109
rect 2706 4081 2736 4109
rect 3022 4081 3052 4109
rect 3286 4081 3316 4109
rect 3602 4081 3632 4109
rect 3866 4081 3896 4109
rect 4182 4081 4212 4109
rect 4446 4081 4476 4109
rect 4762 4081 4792 4109
rect 5026 4081 5056 4109
rect 5342 4081 5372 4109
rect 5606 4081 5636 4109
rect 5922 4081 5952 4109
rect 6186 4081 6216 4109
rect 6502 4081 6532 4109
rect 6766 4081 6796 4109
rect 122 3811 152 3839
rect 386 3811 416 3839
rect 702 3811 732 3839
rect 966 3811 996 3839
rect 1282 3811 1312 3839
rect 1546 3811 1576 3839
rect 1862 3811 1892 3839
rect 2126 3811 2156 3839
rect 2442 3811 2472 3839
rect 2706 3811 2736 3839
rect 3022 3811 3052 3839
rect 3286 3811 3316 3839
rect 3602 3811 3632 3839
rect 3866 3811 3896 3839
rect 4182 3811 4212 3839
rect 4446 3811 4476 3839
rect 4762 3811 4792 3839
rect 5026 3811 5056 3839
rect 5342 3811 5372 3839
rect 5606 3811 5636 3839
rect 5922 3811 5952 3839
rect 6186 3811 6216 3839
rect 6502 3811 6532 3839
rect 6766 3811 6796 3839
rect 122 3541 152 3569
rect 386 3541 416 3569
rect 702 3541 732 3569
rect 966 3541 996 3569
rect 1282 3541 1312 3569
rect 1546 3541 1576 3569
rect 1862 3541 1892 3569
rect 2126 3541 2156 3569
rect 2442 3541 2472 3569
rect 2706 3541 2736 3569
rect 3022 3541 3052 3569
rect 3286 3541 3316 3569
rect 3602 3541 3632 3569
rect 3866 3541 3896 3569
rect 4182 3541 4212 3569
rect 4446 3541 4476 3569
rect 4762 3541 4792 3569
rect 5026 3541 5056 3569
rect 5342 3541 5372 3569
rect 5606 3541 5636 3569
rect 5922 3541 5952 3569
rect 6186 3541 6216 3569
rect 6502 3541 6532 3569
rect 6766 3541 6796 3569
rect 122 3271 152 3299
rect 386 3271 416 3299
rect 702 3271 732 3299
rect 966 3271 996 3299
rect 1282 3271 1312 3299
rect 1546 3271 1576 3299
rect 1862 3271 1892 3299
rect 2126 3271 2156 3299
rect 2442 3271 2472 3299
rect 2706 3271 2736 3299
rect 3022 3271 3052 3299
rect 3286 3271 3316 3299
rect 3602 3271 3632 3299
rect 3866 3271 3896 3299
rect 4182 3271 4212 3299
rect 4446 3271 4476 3299
rect 4762 3271 4792 3299
rect 5026 3271 5056 3299
rect 5342 3271 5372 3299
rect 5606 3271 5636 3299
rect 5922 3271 5952 3299
rect 6186 3271 6216 3299
rect 6502 3271 6532 3299
rect 6766 3271 6796 3299
rect 122 3001 152 3029
rect 386 3001 416 3029
rect 702 3001 732 3029
rect 966 3001 996 3029
rect 1282 3001 1312 3029
rect 1546 3001 1576 3029
rect 1862 3001 1892 3029
rect 2126 3001 2156 3029
rect 2442 3001 2472 3029
rect 2706 3001 2736 3029
rect 3022 3001 3052 3029
rect 3286 3001 3316 3029
rect 3602 3001 3632 3029
rect 3866 3001 3896 3029
rect 4182 3001 4212 3029
rect 4446 3001 4476 3029
rect 4762 3001 4792 3029
rect 5026 3001 5056 3029
rect 5342 3001 5372 3029
rect 5606 3001 5636 3029
rect 5922 3001 5952 3029
rect 6186 3001 6216 3029
rect 6502 3001 6532 3029
rect 6766 3001 6796 3029
rect 122 2731 152 2759
rect 386 2731 416 2759
rect 702 2731 732 2759
rect 966 2731 996 2759
rect 1282 2731 1312 2759
rect 1546 2731 1576 2759
rect 1862 2731 1892 2759
rect 2126 2731 2156 2759
rect 2442 2731 2472 2759
rect 2706 2731 2736 2759
rect 3022 2731 3052 2759
rect 3286 2731 3316 2759
rect 3602 2731 3632 2759
rect 3866 2731 3896 2759
rect 4182 2731 4212 2759
rect 4446 2731 4476 2759
rect 4762 2731 4792 2759
rect 5026 2731 5056 2759
rect 5342 2731 5372 2759
rect 5606 2731 5636 2759
rect 5922 2731 5952 2759
rect 6186 2731 6216 2759
rect 6502 2731 6532 2759
rect 6766 2731 6796 2759
rect 122 2461 152 2489
rect 386 2461 416 2489
rect 702 2461 732 2489
rect 966 2461 996 2489
rect 1282 2461 1312 2489
rect 1546 2461 1576 2489
rect 1862 2461 1892 2489
rect 2126 2461 2156 2489
rect 2442 2461 2472 2489
rect 2706 2461 2736 2489
rect 3022 2461 3052 2489
rect 3286 2461 3316 2489
rect 3602 2461 3632 2489
rect 3866 2461 3896 2489
rect 4182 2461 4212 2489
rect 4446 2461 4476 2489
rect 4762 2461 4792 2489
rect 5026 2461 5056 2489
rect 5342 2461 5372 2489
rect 5606 2461 5636 2489
rect 5922 2461 5952 2489
rect 6186 2461 6216 2489
rect 6502 2461 6532 2489
rect 6766 2461 6796 2489
rect 122 2191 152 2219
rect 386 2191 416 2219
rect 702 2191 732 2219
rect 966 2191 996 2219
rect 1282 2191 1312 2219
rect 1546 2191 1576 2219
rect 1862 2191 1892 2219
rect 2126 2191 2156 2219
rect 2442 2191 2472 2219
rect 2706 2191 2736 2219
rect 3022 2191 3052 2219
rect 3286 2191 3316 2219
rect 3602 2191 3632 2219
rect 3866 2191 3896 2219
rect 4182 2191 4212 2219
rect 4446 2191 4476 2219
rect 4762 2191 4792 2219
rect 5026 2191 5056 2219
rect 5342 2191 5372 2219
rect 5606 2191 5636 2219
rect 5922 2191 5952 2219
rect 6186 2191 6216 2219
rect 6502 2191 6532 2219
rect 6766 2191 6796 2219
rect 122 1921 152 1949
rect 386 1921 416 1949
rect 702 1921 732 1949
rect 966 1921 996 1949
rect 1282 1921 1312 1949
rect 1546 1921 1576 1949
rect 1862 1921 1892 1949
rect 2126 1921 2156 1949
rect 2442 1921 2472 1949
rect 2706 1921 2736 1949
rect 3022 1921 3052 1949
rect 3286 1921 3316 1949
rect 3602 1921 3632 1949
rect 3866 1921 3896 1949
rect 4182 1921 4212 1949
rect 4446 1921 4476 1949
rect 4762 1921 4792 1949
rect 5026 1921 5056 1949
rect 5342 1921 5372 1949
rect 5606 1921 5636 1949
rect 5922 1921 5952 1949
rect 6186 1921 6216 1949
rect 6502 1921 6532 1949
rect 6766 1921 6796 1949
rect 122 1651 152 1679
rect 386 1651 416 1679
rect 702 1651 732 1679
rect 966 1651 996 1679
rect 1282 1651 1312 1679
rect 1546 1651 1576 1679
rect 1862 1651 1892 1679
rect 2126 1651 2156 1679
rect 2442 1651 2472 1679
rect 2706 1651 2736 1679
rect 3022 1651 3052 1679
rect 3286 1651 3316 1679
rect 3602 1651 3632 1679
rect 3866 1651 3896 1679
rect 4182 1651 4212 1679
rect 4446 1651 4476 1679
rect 4762 1651 4792 1679
rect 5026 1651 5056 1679
rect 5342 1651 5372 1679
rect 5606 1651 5636 1679
rect 5922 1651 5952 1679
rect 6186 1651 6216 1679
rect 6502 1651 6532 1679
rect 6766 1651 6796 1679
rect 122 1381 152 1409
rect 386 1381 416 1409
rect 702 1381 732 1409
rect 966 1381 996 1409
rect 1282 1381 1312 1409
rect 1546 1381 1576 1409
rect 1862 1381 1892 1409
rect 2126 1381 2156 1409
rect 2442 1381 2472 1409
rect 2706 1381 2736 1409
rect 3022 1381 3052 1409
rect 3286 1381 3316 1409
rect 3602 1381 3632 1409
rect 3866 1381 3896 1409
rect 4182 1381 4212 1409
rect 4446 1381 4476 1409
rect 4762 1381 4792 1409
rect 5026 1381 5056 1409
rect 5342 1381 5372 1409
rect 5606 1381 5636 1409
rect 5922 1381 5952 1409
rect 6186 1381 6216 1409
rect 6502 1381 6532 1409
rect 6766 1381 6796 1409
rect 122 1111 152 1139
rect 386 1111 416 1139
rect 702 1111 732 1139
rect 966 1111 996 1139
rect 1282 1111 1312 1139
rect 1546 1111 1576 1139
rect 1862 1111 1892 1139
rect 2126 1111 2156 1139
rect 2442 1111 2472 1139
rect 2706 1111 2736 1139
rect 3022 1111 3052 1139
rect 3286 1111 3316 1139
rect 3602 1111 3632 1139
rect 3866 1111 3896 1139
rect 4182 1111 4212 1139
rect 4446 1111 4476 1139
rect 4762 1111 4792 1139
rect 5026 1111 5056 1139
rect 5342 1111 5372 1139
rect 5606 1111 5636 1139
rect 5922 1111 5952 1139
rect 6186 1111 6216 1139
rect 6502 1111 6532 1139
rect 6766 1111 6796 1139
rect 122 841 152 869
rect 386 841 416 869
rect 702 841 732 869
rect 966 841 996 869
rect 1282 841 1312 869
rect 1546 841 1576 869
rect 1862 841 1892 869
rect 2126 841 2156 869
rect 2442 841 2472 869
rect 2706 841 2736 869
rect 3022 841 3052 869
rect 3286 841 3316 869
rect 3602 841 3632 869
rect 3866 841 3896 869
rect 4182 841 4212 869
rect 4446 841 4476 869
rect 4762 841 4792 869
rect 5026 841 5056 869
rect 5342 841 5372 869
rect 5606 841 5636 869
rect 5922 841 5952 869
rect 6186 841 6216 869
rect 6502 841 6532 869
rect 6766 841 6796 869
rect 122 571 152 599
rect 386 571 416 599
rect 702 571 732 599
rect 966 571 996 599
rect 1282 571 1312 599
rect 1546 571 1576 599
rect 1862 571 1892 599
rect 2126 571 2156 599
rect 2442 571 2472 599
rect 2706 571 2736 599
rect 3022 571 3052 599
rect 3286 571 3316 599
rect 3602 571 3632 599
rect 3866 571 3896 599
rect 4182 571 4212 599
rect 4446 571 4476 599
rect 4762 571 4792 599
rect 5026 571 5056 599
rect 5342 571 5372 599
rect 5606 571 5636 599
rect 5922 571 5952 599
rect 6186 571 6216 599
rect 6502 571 6532 599
rect 6766 571 6796 599
rect 122 301 152 329
rect 386 301 416 329
rect 702 301 732 329
rect 966 301 996 329
rect 1282 301 1312 329
rect 1546 301 1576 329
rect 1862 301 1892 329
rect 2126 301 2156 329
rect 2442 301 2472 329
rect 2706 301 2736 329
rect 3022 301 3052 329
rect 3286 301 3316 329
rect 3602 301 3632 329
rect 3866 301 3896 329
rect 4182 301 4212 329
rect 4446 301 4476 329
rect 4762 301 4792 329
rect 5026 301 5056 329
rect 5342 301 5372 329
rect 5606 301 5636 329
rect 5922 301 5952 329
rect 6186 301 6216 329
rect 6502 301 6532 329
rect 6766 301 6796 329
rect 122 31 152 59
rect 386 31 416 59
rect 702 31 732 59
rect 966 31 996 59
rect 1282 31 1312 59
rect 1546 31 1576 59
rect 1862 31 1892 59
rect 2126 31 2156 59
rect 2442 31 2472 59
rect 2706 31 2736 59
rect 3022 31 3052 59
rect 3286 31 3316 59
rect 3602 31 3632 59
rect 3866 31 3896 59
rect 4182 31 4212 59
rect 4446 31 4476 59
rect 4762 31 4792 59
rect 5026 31 5056 59
rect 5342 31 5372 59
rect 5606 31 5636 59
rect 5922 31 5952 59
rect 6186 31 6216 59
rect 6502 31 6532 59
rect 6766 31 6796 59
<< ppu >>
rect 215 4217 245 4245
rect 293 4217 323 4245
rect 795 4217 825 4245
rect 873 4217 903 4245
rect 1375 4217 1405 4245
rect 1453 4217 1483 4245
rect 1955 4217 1985 4245
rect 2033 4217 2063 4245
rect 2535 4217 2565 4245
rect 2613 4217 2643 4245
rect 3115 4217 3145 4245
rect 3193 4217 3223 4245
rect 3695 4217 3725 4245
rect 3773 4217 3803 4245
rect 4275 4217 4305 4245
rect 4353 4217 4383 4245
rect 4855 4217 4885 4245
rect 4933 4217 4963 4245
rect 5435 4217 5465 4245
rect 5513 4217 5543 4245
rect 6015 4217 6045 4245
rect 6093 4217 6123 4245
rect 6595 4217 6625 4245
rect 6673 4217 6703 4245
rect 215 3947 245 3975
rect 293 3947 323 3975
rect 795 3947 825 3975
rect 873 3947 903 3975
rect 1375 3947 1405 3975
rect 1453 3947 1483 3975
rect 1955 3947 1985 3975
rect 2033 3947 2063 3975
rect 2535 3947 2565 3975
rect 2613 3947 2643 3975
rect 3115 3947 3145 3975
rect 3193 3947 3223 3975
rect 3695 3947 3725 3975
rect 3773 3947 3803 3975
rect 4275 3947 4305 3975
rect 4353 3947 4383 3975
rect 4855 3947 4885 3975
rect 4933 3947 4963 3975
rect 5435 3947 5465 3975
rect 5513 3947 5543 3975
rect 6015 3947 6045 3975
rect 6093 3947 6123 3975
rect 6595 3947 6625 3975
rect 6673 3947 6703 3975
rect 215 3677 245 3705
rect 293 3677 323 3705
rect 795 3677 825 3705
rect 873 3677 903 3705
rect 1375 3677 1405 3705
rect 1453 3677 1483 3705
rect 1955 3677 1985 3705
rect 2033 3677 2063 3705
rect 2535 3677 2565 3705
rect 2613 3677 2643 3705
rect 3115 3677 3145 3705
rect 3193 3677 3223 3705
rect 3695 3677 3725 3705
rect 3773 3677 3803 3705
rect 4275 3677 4305 3705
rect 4353 3677 4383 3705
rect 4855 3677 4885 3705
rect 4933 3677 4963 3705
rect 5435 3677 5465 3705
rect 5513 3677 5543 3705
rect 6015 3677 6045 3705
rect 6093 3677 6123 3705
rect 6595 3677 6625 3705
rect 6673 3677 6703 3705
rect 215 3407 245 3435
rect 293 3407 323 3435
rect 795 3407 825 3435
rect 873 3407 903 3435
rect 1375 3407 1405 3435
rect 1453 3407 1483 3435
rect 1955 3407 1985 3435
rect 2033 3407 2063 3435
rect 2535 3407 2565 3435
rect 2613 3407 2643 3435
rect 3115 3407 3145 3435
rect 3193 3407 3223 3435
rect 3695 3407 3725 3435
rect 3773 3407 3803 3435
rect 4275 3407 4305 3435
rect 4353 3407 4383 3435
rect 4855 3407 4885 3435
rect 4933 3407 4963 3435
rect 5435 3407 5465 3435
rect 5513 3407 5543 3435
rect 6015 3407 6045 3435
rect 6093 3407 6123 3435
rect 6595 3407 6625 3435
rect 6673 3407 6703 3435
rect 215 3137 245 3165
rect 293 3137 323 3165
rect 795 3137 825 3165
rect 873 3137 903 3165
rect 1375 3137 1405 3165
rect 1453 3137 1483 3165
rect 1955 3137 1985 3165
rect 2033 3137 2063 3165
rect 2535 3137 2565 3165
rect 2613 3137 2643 3165
rect 3115 3137 3145 3165
rect 3193 3137 3223 3165
rect 3695 3137 3725 3165
rect 3773 3137 3803 3165
rect 4275 3137 4305 3165
rect 4353 3137 4383 3165
rect 4855 3137 4885 3165
rect 4933 3137 4963 3165
rect 5435 3137 5465 3165
rect 5513 3137 5543 3165
rect 6015 3137 6045 3165
rect 6093 3137 6123 3165
rect 6595 3137 6625 3165
rect 6673 3137 6703 3165
rect 215 2867 245 2895
rect 293 2867 323 2895
rect 795 2867 825 2895
rect 873 2867 903 2895
rect 1375 2867 1405 2895
rect 1453 2867 1483 2895
rect 1955 2867 1985 2895
rect 2033 2867 2063 2895
rect 2535 2867 2565 2895
rect 2613 2867 2643 2895
rect 3115 2867 3145 2895
rect 3193 2867 3223 2895
rect 3695 2867 3725 2895
rect 3773 2867 3803 2895
rect 4275 2867 4305 2895
rect 4353 2867 4383 2895
rect 4855 2867 4885 2895
rect 4933 2867 4963 2895
rect 5435 2867 5465 2895
rect 5513 2867 5543 2895
rect 6015 2867 6045 2895
rect 6093 2867 6123 2895
rect 6595 2867 6625 2895
rect 6673 2867 6703 2895
rect 215 2597 245 2625
rect 293 2597 323 2625
rect 795 2597 825 2625
rect 873 2597 903 2625
rect 1375 2597 1405 2625
rect 1453 2597 1483 2625
rect 1955 2597 1985 2625
rect 2033 2597 2063 2625
rect 2535 2597 2565 2625
rect 2613 2597 2643 2625
rect 3115 2597 3145 2625
rect 3193 2597 3223 2625
rect 3695 2597 3725 2625
rect 3773 2597 3803 2625
rect 4275 2597 4305 2625
rect 4353 2597 4383 2625
rect 4855 2597 4885 2625
rect 4933 2597 4963 2625
rect 5435 2597 5465 2625
rect 5513 2597 5543 2625
rect 6015 2597 6045 2625
rect 6093 2597 6123 2625
rect 6595 2597 6625 2625
rect 6673 2597 6703 2625
rect 215 2327 245 2355
rect 293 2327 323 2355
rect 795 2327 825 2355
rect 873 2327 903 2355
rect 1375 2327 1405 2355
rect 1453 2327 1483 2355
rect 1955 2327 1985 2355
rect 2033 2327 2063 2355
rect 2535 2327 2565 2355
rect 2613 2327 2643 2355
rect 3115 2327 3145 2355
rect 3193 2327 3223 2355
rect 3695 2327 3725 2355
rect 3773 2327 3803 2355
rect 4275 2327 4305 2355
rect 4353 2327 4383 2355
rect 4855 2327 4885 2355
rect 4933 2327 4963 2355
rect 5435 2327 5465 2355
rect 5513 2327 5543 2355
rect 6015 2327 6045 2355
rect 6093 2327 6123 2355
rect 6595 2327 6625 2355
rect 6673 2327 6703 2355
rect 215 2057 245 2085
rect 293 2057 323 2085
rect 795 2057 825 2085
rect 873 2057 903 2085
rect 1375 2057 1405 2085
rect 1453 2057 1483 2085
rect 1955 2057 1985 2085
rect 2033 2057 2063 2085
rect 2535 2057 2565 2085
rect 2613 2057 2643 2085
rect 3115 2057 3145 2085
rect 3193 2057 3223 2085
rect 3695 2057 3725 2085
rect 3773 2057 3803 2085
rect 4275 2057 4305 2085
rect 4353 2057 4383 2085
rect 4855 2057 4885 2085
rect 4933 2057 4963 2085
rect 5435 2057 5465 2085
rect 5513 2057 5543 2085
rect 6015 2057 6045 2085
rect 6093 2057 6123 2085
rect 6595 2057 6625 2085
rect 6673 2057 6703 2085
rect 215 1787 245 1815
rect 293 1787 323 1815
rect 795 1787 825 1815
rect 873 1787 903 1815
rect 1375 1787 1405 1815
rect 1453 1787 1483 1815
rect 1955 1787 1985 1815
rect 2033 1787 2063 1815
rect 2535 1787 2565 1815
rect 2613 1787 2643 1815
rect 3115 1787 3145 1815
rect 3193 1787 3223 1815
rect 3695 1787 3725 1815
rect 3773 1787 3803 1815
rect 4275 1787 4305 1815
rect 4353 1787 4383 1815
rect 4855 1787 4885 1815
rect 4933 1787 4963 1815
rect 5435 1787 5465 1815
rect 5513 1787 5543 1815
rect 6015 1787 6045 1815
rect 6093 1787 6123 1815
rect 6595 1787 6625 1815
rect 6673 1787 6703 1815
rect 215 1517 245 1545
rect 293 1517 323 1545
rect 795 1517 825 1545
rect 873 1517 903 1545
rect 1375 1517 1405 1545
rect 1453 1517 1483 1545
rect 1955 1517 1985 1545
rect 2033 1517 2063 1545
rect 2535 1517 2565 1545
rect 2613 1517 2643 1545
rect 3115 1517 3145 1545
rect 3193 1517 3223 1545
rect 3695 1517 3725 1545
rect 3773 1517 3803 1545
rect 4275 1517 4305 1545
rect 4353 1517 4383 1545
rect 4855 1517 4885 1545
rect 4933 1517 4963 1545
rect 5435 1517 5465 1545
rect 5513 1517 5543 1545
rect 6015 1517 6045 1545
rect 6093 1517 6123 1545
rect 6595 1517 6625 1545
rect 6673 1517 6703 1545
rect 215 1247 245 1275
rect 293 1247 323 1275
rect 795 1247 825 1275
rect 873 1247 903 1275
rect 1375 1247 1405 1275
rect 1453 1247 1483 1275
rect 1955 1247 1985 1275
rect 2033 1247 2063 1275
rect 2535 1247 2565 1275
rect 2613 1247 2643 1275
rect 3115 1247 3145 1275
rect 3193 1247 3223 1275
rect 3695 1247 3725 1275
rect 3773 1247 3803 1275
rect 4275 1247 4305 1275
rect 4353 1247 4383 1275
rect 4855 1247 4885 1275
rect 4933 1247 4963 1275
rect 5435 1247 5465 1275
rect 5513 1247 5543 1275
rect 6015 1247 6045 1275
rect 6093 1247 6123 1275
rect 6595 1247 6625 1275
rect 6673 1247 6703 1275
rect 215 977 245 1005
rect 293 977 323 1005
rect 795 977 825 1005
rect 873 977 903 1005
rect 1375 977 1405 1005
rect 1453 977 1483 1005
rect 1955 977 1985 1005
rect 2033 977 2063 1005
rect 2535 977 2565 1005
rect 2613 977 2643 1005
rect 3115 977 3145 1005
rect 3193 977 3223 1005
rect 3695 977 3725 1005
rect 3773 977 3803 1005
rect 4275 977 4305 1005
rect 4353 977 4383 1005
rect 4855 977 4885 1005
rect 4933 977 4963 1005
rect 5435 977 5465 1005
rect 5513 977 5543 1005
rect 6015 977 6045 1005
rect 6093 977 6123 1005
rect 6595 977 6625 1005
rect 6673 977 6703 1005
rect 215 707 245 735
rect 293 707 323 735
rect 795 707 825 735
rect 873 707 903 735
rect 1375 707 1405 735
rect 1453 707 1483 735
rect 1955 707 1985 735
rect 2033 707 2063 735
rect 2535 707 2565 735
rect 2613 707 2643 735
rect 3115 707 3145 735
rect 3193 707 3223 735
rect 3695 707 3725 735
rect 3773 707 3803 735
rect 4275 707 4305 735
rect 4353 707 4383 735
rect 4855 707 4885 735
rect 4933 707 4963 735
rect 5435 707 5465 735
rect 5513 707 5543 735
rect 6015 707 6045 735
rect 6093 707 6123 735
rect 6595 707 6625 735
rect 6673 707 6703 735
rect 215 437 245 465
rect 293 437 323 465
rect 795 437 825 465
rect 873 437 903 465
rect 1375 437 1405 465
rect 1453 437 1483 465
rect 1955 437 1985 465
rect 2033 437 2063 465
rect 2535 437 2565 465
rect 2613 437 2643 465
rect 3115 437 3145 465
rect 3193 437 3223 465
rect 3695 437 3725 465
rect 3773 437 3803 465
rect 4275 437 4305 465
rect 4353 437 4383 465
rect 4855 437 4885 465
rect 4933 437 4963 465
rect 5435 437 5465 465
rect 5513 437 5543 465
rect 6015 437 6045 465
rect 6093 437 6123 465
rect 6595 437 6625 465
rect 6673 437 6703 465
rect 215 167 245 195
rect 293 167 323 195
rect 795 167 825 195
rect 873 167 903 195
rect 1375 167 1405 195
rect 1453 167 1483 195
rect 1955 167 1985 195
rect 2033 167 2063 195
rect 2535 167 2565 195
rect 2613 167 2643 195
rect 3115 167 3145 195
rect 3193 167 3223 195
rect 3695 167 3725 195
rect 3773 167 3803 195
rect 4275 167 4305 195
rect 4353 167 4383 195
rect 4855 167 4885 195
rect 4933 167 4963 195
rect 5435 167 5465 195
rect 5513 167 5543 195
rect 6015 167 6045 195
rect 6093 167 6123 195
rect 6595 167 6625 195
rect 6673 167 6703 195
<< ndiff >>
rect 82 4227 100 4255
rect 130 4227 148 4255
rect 390 4227 408 4255
rect 438 4227 457 4255
rect 662 4227 680 4255
rect 710 4227 728 4255
rect 970 4227 988 4255
rect 1018 4227 1037 4255
rect 1242 4227 1260 4255
rect 1290 4227 1308 4255
rect 1550 4227 1568 4255
rect 1598 4227 1617 4255
rect 1822 4227 1840 4255
rect 1870 4227 1888 4255
rect 2130 4227 2148 4255
rect 2178 4227 2197 4255
rect 2402 4227 2420 4255
rect 2450 4227 2468 4255
rect 2710 4227 2728 4255
rect 2758 4227 2777 4255
rect 2982 4227 3000 4255
rect 3030 4227 3048 4255
rect 3290 4227 3308 4255
rect 3338 4227 3357 4255
rect 3562 4227 3580 4255
rect 3610 4227 3628 4255
rect 3870 4227 3888 4255
rect 3918 4227 3937 4255
rect 4142 4227 4160 4255
rect 4190 4227 4208 4255
rect 4450 4227 4468 4255
rect 4498 4227 4517 4255
rect 4722 4227 4740 4255
rect 4770 4227 4788 4255
rect 5030 4227 5048 4255
rect 5078 4227 5097 4255
rect 5302 4227 5320 4255
rect 5350 4227 5368 4255
rect 5610 4227 5628 4255
rect 5658 4227 5677 4255
rect 5882 4227 5900 4255
rect 5930 4227 5948 4255
rect 6190 4227 6208 4255
rect 6238 4227 6257 4255
rect 6462 4227 6480 4255
rect 6510 4227 6528 4255
rect 6770 4227 6788 4255
rect 6818 4227 6837 4255
rect 8 4081 36 4123
rect 66 4109 91 4123
rect 190 4113 215 4123
rect 66 4081 122 4109
rect 152 4081 186 4109
tri 200 4106 207 4113 ne
rect 207 4081 215 4113
rect 245 4081 293 4123
rect 323 4113 348 4123
rect 323 4081 331 4113
rect 447 4109 472 4123
rect 352 4081 386 4109
rect 416 4081 472 4109
rect 502 4081 530 4123
rect 588 4081 616 4123
rect 646 4109 671 4123
rect 770 4113 795 4123
rect 646 4081 702 4109
rect 732 4081 766 4109
tri 780 4106 787 4113 ne
rect 787 4081 795 4113
rect 825 4081 873 4123
rect 903 4113 928 4123
rect 903 4081 911 4113
rect 1027 4109 1052 4123
rect 932 4081 966 4109
rect 996 4081 1052 4109
rect 1082 4081 1110 4123
rect 1168 4081 1196 4123
rect 1226 4109 1251 4123
rect 1350 4113 1375 4123
rect 1226 4081 1282 4109
rect 1312 4081 1346 4109
tri 1360 4106 1367 4113 ne
rect 1367 4081 1375 4113
rect 1405 4081 1453 4123
rect 1483 4113 1508 4123
rect 1483 4081 1491 4113
rect 1607 4109 1632 4123
rect 1512 4081 1546 4109
rect 1576 4081 1632 4109
rect 1662 4081 1690 4123
rect 1748 4081 1776 4123
rect 1806 4109 1831 4123
rect 1930 4113 1955 4123
rect 1806 4081 1862 4109
rect 1892 4081 1926 4109
tri 1940 4106 1947 4113 ne
rect 1947 4081 1955 4113
rect 1985 4081 2033 4123
rect 2063 4113 2088 4123
rect 2063 4081 2071 4113
rect 2187 4109 2212 4123
rect 2092 4081 2126 4109
rect 2156 4081 2212 4109
rect 2242 4081 2270 4123
rect 2328 4081 2356 4123
rect 2386 4109 2411 4123
rect 2510 4113 2535 4123
rect 2386 4081 2442 4109
rect 2472 4081 2506 4109
tri 2520 4106 2527 4113 ne
rect 2527 4081 2535 4113
rect 2565 4081 2613 4123
rect 2643 4113 2668 4123
rect 2643 4081 2651 4113
rect 2767 4109 2792 4123
rect 2672 4081 2706 4109
rect 2736 4081 2792 4109
rect 2822 4081 2850 4123
rect 2908 4081 2936 4123
rect 2966 4109 2991 4123
rect 3090 4113 3115 4123
rect 2966 4081 3022 4109
rect 3052 4081 3086 4109
tri 3100 4106 3107 4113 ne
rect 3107 4081 3115 4113
rect 3145 4081 3193 4123
rect 3223 4113 3248 4123
rect 3223 4081 3231 4113
rect 3347 4109 3372 4123
rect 3252 4081 3286 4109
rect 3316 4081 3372 4109
rect 3402 4081 3430 4123
rect 3488 4081 3516 4123
rect 3546 4109 3571 4123
rect 3670 4113 3695 4123
rect 3546 4081 3602 4109
rect 3632 4081 3666 4109
tri 3680 4106 3687 4113 ne
rect 3687 4081 3695 4113
rect 3725 4081 3773 4123
rect 3803 4113 3828 4123
rect 3803 4081 3811 4113
rect 3927 4109 3952 4123
rect 3832 4081 3866 4109
rect 3896 4081 3952 4109
rect 3982 4081 4010 4123
rect 4068 4081 4096 4123
rect 4126 4109 4151 4123
rect 4250 4113 4275 4123
rect 4126 4081 4182 4109
rect 4212 4081 4246 4109
tri 4260 4106 4267 4113 ne
rect 4267 4081 4275 4113
rect 4305 4081 4353 4123
rect 4383 4113 4408 4123
rect 4383 4081 4391 4113
rect 4507 4109 4532 4123
rect 4412 4081 4446 4109
rect 4476 4081 4532 4109
rect 4562 4081 4590 4123
rect 4648 4081 4676 4123
rect 4706 4109 4731 4123
rect 4830 4113 4855 4123
rect 4706 4081 4762 4109
rect 4792 4081 4826 4109
tri 4840 4106 4847 4113 ne
rect 4847 4081 4855 4113
rect 4885 4081 4933 4123
rect 4963 4113 4988 4123
rect 4963 4081 4971 4113
rect 5087 4109 5112 4123
rect 4992 4081 5026 4109
rect 5056 4081 5112 4109
rect 5142 4081 5170 4123
rect 5228 4081 5256 4123
rect 5286 4109 5311 4123
rect 5410 4113 5435 4123
rect 5286 4081 5342 4109
rect 5372 4081 5406 4109
tri 5420 4106 5427 4113 ne
rect 5427 4081 5435 4113
rect 5465 4081 5513 4123
rect 5543 4113 5568 4123
rect 5543 4081 5551 4113
rect 5667 4109 5692 4123
rect 5572 4081 5606 4109
rect 5636 4081 5692 4109
rect 5722 4081 5750 4123
rect 5808 4081 5836 4123
rect 5866 4109 5891 4123
rect 5990 4113 6015 4123
rect 5866 4081 5922 4109
rect 5952 4081 5986 4109
tri 6000 4106 6007 4113 ne
rect 6007 4081 6015 4113
rect 6045 4081 6093 4123
rect 6123 4113 6148 4123
rect 6123 4081 6131 4113
rect 6247 4109 6272 4123
rect 6152 4081 6186 4109
rect 6216 4081 6272 4109
rect 6302 4081 6330 4123
rect 6388 4081 6416 4123
rect 6446 4109 6471 4123
rect 6570 4113 6595 4123
rect 6446 4081 6502 4109
rect 6532 4081 6566 4109
tri 6580 4106 6587 4113 ne
rect 6587 4081 6595 4113
rect 6625 4081 6673 4123
rect 6703 4113 6728 4123
rect 6703 4081 6711 4113
rect 6827 4109 6852 4123
rect 6732 4081 6766 4109
rect 6796 4081 6852 4109
rect 6882 4081 6910 4123
rect 159 4057 186 4081
rect 253 4059 285 4081
rect 253 4057 255 4059
rect 283 4057 285 4059
rect 352 4057 379 4081
rect 159 4043 253 4057
rect 285 4043 379 4057
rect 739 4057 766 4081
rect 833 4059 865 4081
rect 833 4057 835 4059
rect 863 4057 865 4059
rect 932 4057 959 4081
rect 739 4043 833 4057
rect 865 4043 959 4057
rect 1319 4057 1346 4081
rect 1413 4059 1445 4081
rect 1413 4057 1415 4059
rect 1443 4057 1445 4059
rect 1512 4057 1539 4081
rect 1319 4043 1413 4057
rect 1445 4043 1539 4057
rect 1899 4057 1926 4081
rect 1993 4059 2025 4081
rect 1993 4057 1995 4059
rect 2023 4057 2025 4059
rect 2092 4057 2119 4081
rect 1899 4043 1993 4057
rect 2025 4043 2119 4057
rect 2479 4057 2506 4081
rect 2573 4059 2605 4081
rect 2573 4057 2575 4059
rect 2603 4057 2605 4059
rect 2672 4057 2699 4081
rect 2479 4043 2573 4057
rect 2605 4043 2699 4057
rect 3059 4057 3086 4081
rect 3153 4059 3185 4081
rect 3153 4057 3155 4059
rect 3183 4057 3185 4059
rect 3252 4057 3279 4081
rect 3059 4043 3153 4057
rect 3185 4043 3279 4057
rect 3639 4057 3666 4081
rect 3733 4059 3765 4081
rect 3733 4057 3735 4059
rect 3763 4057 3765 4059
rect 3832 4057 3859 4081
rect 3639 4043 3733 4057
rect 3765 4043 3859 4057
rect 4219 4057 4246 4081
rect 4313 4059 4345 4081
rect 4313 4057 4315 4059
rect 4343 4057 4345 4059
rect 4412 4057 4439 4081
rect 4219 4043 4313 4057
rect 4345 4043 4439 4057
rect 4799 4057 4826 4081
rect 4893 4059 4925 4081
rect 4893 4057 4895 4059
rect 4923 4057 4925 4059
rect 4992 4057 5019 4081
rect 4799 4043 4893 4057
rect 4925 4043 5019 4057
rect 5379 4057 5406 4081
rect 5473 4059 5505 4081
rect 5473 4057 5475 4059
rect 5503 4057 5505 4059
rect 5572 4057 5599 4081
rect 5379 4043 5473 4057
rect 5505 4043 5599 4057
rect 5959 4057 5986 4081
rect 6053 4059 6085 4081
rect 6053 4057 6055 4059
rect 6083 4057 6085 4059
rect 6152 4057 6179 4081
rect 5959 4043 6053 4057
rect 6085 4043 6179 4057
rect 6539 4057 6566 4081
rect 6633 4059 6665 4081
rect 6633 4057 6635 4059
rect 6663 4057 6665 4059
rect 6732 4057 6759 4081
rect 6539 4043 6633 4057
rect 6665 4043 6759 4057
rect 82 3957 100 3985
rect 130 3957 148 3985
rect 390 3957 408 3985
rect 438 3957 457 3985
rect 662 3957 680 3985
rect 710 3957 728 3985
rect 970 3957 988 3985
rect 1018 3957 1037 3985
rect 1242 3957 1260 3985
rect 1290 3957 1308 3985
rect 1550 3957 1568 3985
rect 1598 3957 1617 3985
rect 1822 3957 1840 3985
rect 1870 3957 1888 3985
rect 2130 3957 2148 3985
rect 2178 3957 2197 3985
rect 2402 3957 2420 3985
rect 2450 3957 2468 3985
rect 2710 3957 2728 3985
rect 2758 3957 2777 3985
rect 2982 3957 3000 3985
rect 3030 3957 3048 3985
rect 3290 3957 3308 3985
rect 3338 3957 3357 3985
rect 3562 3957 3580 3985
rect 3610 3957 3628 3985
rect 3870 3957 3888 3985
rect 3918 3957 3937 3985
rect 4142 3957 4160 3985
rect 4190 3957 4208 3985
rect 4450 3957 4468 3985
rect 4498 3957 4517 3985
rect 4722 3957 4740 3985
rect 4770 3957 4788 3985
rect 5030 3957 5048 3985
rect 5078 3957 5097 3985
rect 5302 3957 5320 3985
rect 5350 3957 5368 3985
rect 5610 3957 5628 3985
rect 5658 3957 5677 3985
rect 5882 3957 5900 3985
rect 5930 3957 5948 3985
rect 6190 3957 6208 3985
rect 6238 3957 6257 3985
rect 6462 3957 6480 3985
rect 6510 3957 6528 3985
rect 6770 3957 6788 3985
rect 6818 3957 6837 3985
rect 8 3811 36 3853
rect 66 3839 91 3853
rect 190 3843 215 3853
rect 66 3811 122 3839
rect 152 3811 186 3839
tri 200 3836 207 3843 ne
rect 207 3811 215 3843
rect 245 3811 293 3853
rect 323 3843 348 3853
rect 323 3811 331 3843
rect 447 3839 472 3853
rect 352 3811 386 3839
rect 416 3811 472 3839
rect 502 3811 530 3853
rect 588 3811 616 3853
rect 646 3839 671 3853
rect 770 3843 795 3853
rect 646 3811 702 3839
rect 732 3811 766 3839
tri 780 3836 787 3843 ne
rect 787 3811 795 3843
rect 825 3811 873 3853
rect 903 3843 928 3853
rect 903 3811 911 3843
rect 1027 3839 1052 3853
rect 932 3811 966 3839
rect 996 3811 1052 3839
rect 1082 3811 1110 3853
rect 1168 3811 1196 3853
rect 1226 3839 1251 3853
rect 1350 3843 1375 3853
rect 1226 3811 1282 3839
rect 1312 3811 1346 3839
tri 1360 3836 1367 3843 ne
rect 1367 3811 1375 3843
rect 1405 3811 1453 3853
rect 1483 3843 1508 3853
rect 1483 3811 1491 3843
rect 1607 3839 1632 3853
rect 1512 3811 1546 3839
rect 1576 3811 1632 3839
rect 1662 3811 1690 3853
rect 1748 3811 1776 3853
rect 1806 3839 1831 3853
rect 1930 3843 1955 3853
rect 1806 3811 1862 3839
rect 1892 3811 1926 3839
tri 1940 3836 1947 3843 ne
rect 1947 3811 1955 3843
rect 1985 3811 2033 3853
rect 2063 3843 2088 3853
rect 2063 3811 2071 3843
rect 2187 3839 2212 3853
rect 2092 3811 2126 3839
rect 2156 3811 2212 3839
rect 2242 3811 2270 3853
rect 2328 3811 2356 3853
rect 2386 3839 2411 3853
rect 2510 3843 2535 3853
rect 2386 3811 2442 3839
rect 2472 3811 2506 3839
tri 2520 3836 2527 3843 ne
rect 2527 3811 2535 3843
rect 2565 3811 2613 3853
rect 2643 3843 2668 3853
rect 2643 3811 2651 3843
rect 2767 3839 2792 3853
rect 2672 3811 2706 3839
rect 2736 3811 2792 3839
rect 2822 3811 2850 3853
rect 2908 3811 2936 3853
rect 2966 3839 2991 3853
rect 3090 3843 3115 3853
rect 2966 3811 3022 3839
rect 3052 3811 3086 3839
tri 3100 3836 3107 3843 ne
rect 3107 3811 3115 3843
rect 3145 3811 3193 3853
rect 3223 3843 3248 3853
rect 3223 3811 3231 3843
rect 3347 3839 3372 3853
rect 3252 3811 3286 3839
rect 3316 3811 3372 3839
rect 3402 3811 3430 3853
rect 3488 3811 3516 3853
rect 3546 3839 3571 3853
rect 3670 3843 3695 3853
rect 3546 3811 3602 3839
rect 3632 3811 3666 3839
tri 3680 3836 3687 3843 ne
rect 3687 3811 3695 3843
rect 3725 3811 3773 3853
rect 3803 3843 3828 3853
rect 3803 3811 3811 3843
rect 3927 3839 3952 3853
rect 3832 3811 3866 3839
rect 3896 3811 3952 3839
rect 3982 3811 4010 3853
rect 4068 3811 4096 3853
rect 4126 3839 4151 3853
rect 4250 3843 4275 3853
rect 4126 3811 4182 3839
rect 4212 3811 4246 3839
tri 4260 3836 4267 3843 ne
rect 4267 3811 4275 3843
rect 4305 3811 4353 3853
rect 4383 3843 4408 3853
rect 4383 3811 4391 3843
rect 4507 3839 4532 3853
rect 4412 3811 4446 3839
rect 4476 3811 4532 3839
rect 4562 3811 4590 3853
rect 4648 3811 4676 3853
rect 4706 3839 4731 3853
rect 4830 3843 4855 3853
rect 4706 3811 4762 3839
rect 4792 3811 4826 3839
tri 4840 3836 4847 3843 ne
rect 4847 3811 4855 3843
rect 4885 3811 4933 3853
rect 4963 3843 4988 3853
rect 4963 3811 4971 3843
rect 5087 3839 5112 3853
rect 4992 3811 5026 3839
rect 5056 3811 5112 3839
rect 5142 3811 5170 3853
rect 5228 3811 5256 3853
rect 5286 3839 5311 3853
rect 5410 3843 5435 3853
rect 5286 3811 5342 3839
rect 5372 3811 5406 3839
tri 5420 3836 5427 3843 ne
rect 5427 3811 5435 3843
rect 5465 3811 5513 3853
rect 5543 3843 5568 3853
rect 5543 3811 5551 3843
rect 5667 3839 5692 3853
rect 5572 3811 5606 3839
rect 5636 3811 5692 3839
rect 5722 3811 5750 3853
rect 5808 3811 5836 3853
rect 5866 3839 5891 3853
rect 5990 3843 6015 3853
rect 5866 3811 5922 3839
rect 5952 3811 5986 3839
tri 6000 3836 6007 3843 ne
rect 6007 3811 6015 3843
rect 6045 3811 6093 3853
rect 6123 3843 6148 3853
rect 6123 3811 6131 3843
rect 6247 3839 6272 3853
rect 6152 3811 6186 3839
rect 6216 3811 6272 3839
rect 6302 3811 6330 3853
rect 6388 3811 6416 3853
rect 6446 3839 6471 3853
rect 6570 3843 6595 3853
rect 6446 3811 6502 3839
rect 6532 3811 6566 3839
tri 6580 3836 6587 3843 ne
rect 6587 3811 6595 3843
rect 6625 3811 6673 3853
rect 6703 3843 6728 3853
rect 6703 3811 6711 3843
rect 6827 3839 6852 3853
rect 6732 3811 6766 3839
rect 6796 3811 6852 3839
rect 6882 3811 6910 3853
rect 159 3787 186 3811
rect 253 3789 285 3811
rect 253 3787 255 3789
rect 283 3787 285 3789
rect 352 3787 379 3811
rect 159 3773 253 3787
rect 285 3773 379 3787
rect 739 3787 766 3811
rect 833 3789 865 3811
rect 833 3787 835 3789
rect 863 3787 865 3789
rect 932 3787 959 3811
rect 739 3773 833 3787
rect 865 3773 959 3787
rect 1319 3787 1346 3811
rect 1413 3789 1445 3811
rect 1413 3787 1415 3789
rect 1443 3787 1445 3789
rect 1512 3787 1539 3811
rect 1319 3773 1413 3787
rect 1445 3773 1539 3787
rect 1899 3787 1926 3811
rect 1993 3789 2025 3811
rect 1993 3787 1995 3789
rect 2023 3787 2025 3789
rect 2092 3787 2119 3811
rect 1899 3773 1993 3787
rect 2025 3773 2119 3787
rect 2479 3787 2506 3811
rect 2573 3789 2605 3811
rect 2573 3787 2575 3789
rect 2603 3787 2605 3789
rect 2672 3787 2699 3811
rect 2479 3773 2573 3787
rect 2605 3773 2699 3787
rect 3059 3787 3086 3811
rect 3153 3789 3185 3811
rect 3153 3787 3155 3789
rect 3183 3787 3185 3789
rect 3252 3787 3279 3811
rect 3059 3773 3153 3787
rect 3185 3773 3279 3787
rect 3639 3787 3666 3811
rect 3733 3789 3765 3811
rect 3733 3787 3735 3789
rect 3763 3787 3765 3789
rect 3832 3787 3859 3811
rect 3639 3773 3733 3787
rect 3765 3773 3859 3787
rect 4219 3787 4246 3811
rect 4313 3789 4345 3811
rect 4313 3787 4315 3789
rect 4343 3787 4345 3789
rect 4412 3787 4439 3811
rect 4219 3773 4313 3787
rect 4345 3773 4439 3787
rect 4799 3787 4826 3811
rect 4893 3789 4925 3811
rect 4893 3787 4895 3789
rect 4923 3787 4925 3789
rect 4992 3787 5019 3811
rect 4799 3773 4893 3787
rect 4925 3773 5019 3787
rect 5379 3787 5406 3811
rect 5473 3789 5505 3811
rect 5473 3787 5475 3789
rect 5503 3787 5505 3789
rect 5572 3787 5599 3811
rect 5379 3773 5473 3787
rect 5505 3773 5599 3787
rect 5959 3787 5986 3811
rect 6053 3789 6085 3811
rect 6053 3787 6055 3789
rect 6083 3787 6085 3789
rect 6152 3787 6179 3811
rect 5959 3773 6053 3787
rect 6085 3773 6179 3787
rect 6539 3787 6566 3811
rect 6633 3789 6665 3811
rect 6633 3787 6635 3789
rect 6663 3787 6665 3789
rect 6732 3787 6759 3811
rect 6539 3773 6633 3787
rect 6665 3773 6759 3787
rect 82 3687 100 3715
rect 130 3687 148 3715
rect 390 3687 408 3715
rect 438 3687 457 3715
rect 662 3687 680 3715
rect 710 3687 728 3715
rect 970 3687 988 3715
rect 1018 3687 1037 3715
rect 1242 3687 1260 3715
rect 1290 3687 1308 3715
rect 1550 3687 1568 3715
rect 1598 3687 1617 3715
rect 1822 3687 1840 3715
rect 1870 3687 1888 3715
rect 2130 3687 2148 3715
rect 2178 3687 2197 3715
rect 2402 3687 2420 3715
rect 2450 3687 2468 3715
rect 2710 3687 2728 3715
rect 2758 3687 2777 3715
rect 2982 3687 3000 3715
rect 3030 3687 3048 3715
rect 3290 3687 3308 3715
rect 3338 3687 3357 3715
rect 3562 3687 3580 3715
rect 3610 3687 3628 3715
rect 3870 3687 3888 3715
rect 3918 3687 3937 3715
rect 4142 3687 4160 3715
rect 4190 3687 4208 3715
rect 4450 3687 4468 3715
rect 4498 3687 4517 3715
rect 4722 3687 4740 3715
rect 4770 3687 4788 3715
rect 5030 3687 5048 3715
rect 5078 3687 5097 3715
rect 5302 3687 5320 3715
rect 5350 3687 5368 3715
rect 5610 3687 5628 3715
rect 5658 3687 5677 3715
rect 5882 3687 5900 3715
rect 5930 3687 5948 3715
rect 6190 3687 6208 3715
rect 6238 3687 6257 3715
rect 6462 3687 6480 3715
rect 6510 3687 6528 3715
rect 6770 3687 6788 3715
rect 6818 3687 6837 3715
rect 8 3541 36 3583
rect 66 3569 91 3583
rect 190 3573 215 3583
rect 66 3541 122 3569
rect 152 3541 186 3569
tri 200 3566 207 3573 ne
rect 207 3541 215 3573
rect 245 3541 293 3583
rect 323 3573 348 3583
rect 323 3541 331 3573
rect 447 3569 472 3583
rect 352 3541 386 3569
rect 416 3541 472 3569
rect 502 3541 530 3583
rect 588 3541 616 3583
rect 646 3569 671 3583
rect 770 3573 795 3583
rect 646 3541 702 3569
rect 732 3541 766 3569
tri 780 3566 787 3573 ne
rect 787 3541 795 3573
rect 825 3541 873 3583
rect 903 3573 928 3583
rect 903 3541 911 3573
rect 1027 3569 1052 3583
rect 932 3541 966 3569
rect 996 3541 1052 3569
rect 1082 3541 1110 3583
rect 1168 3541 1196 3583
rect 1226 3569 1251 3583
rect 1350 3573 1375 3583
rect 1226 3541 1282 3569
rect 1312 3541 1346 3569
tri 1360 3566 1367 3573 ne
rect 1367 3541 1375 3573
rect 1405 3541 1453 3583
rect 1483 3573 1508 3583
rect 1483 3541 1491 3573
rect 1607 3569 1632 3583
rect 1512 3541 1546 3569
rect 1576 3541 1632 3569
rect 1662 3541 1690 3583
rect 1748 3541 1776 3583
rect 1806 3569 1831 3583
rect 1930 3573 1955 3583
rect 1806 3541 1862 3569
rect 1892 3541 1926 3569
tri 1940 3566 1947 3573 ne
rect 1947 3541 1955 3573
rect 1985 3541 2033 3583
rect 2063 3573 2088 3583
rect 2063 3541 2071 3573
rect 2187 3569 2212 3583
rect 2092 3541 2126 3569
rect 2156 3541 2212 3569
rect 2242 3541 2270 3583
rect 2328 3541 2356 3583
rect 2386 3569 2411 3583
rect 2510 3573 2535 3583
rect 2386 3541 2442 3569
rect 2472 3541 2506 3569
tri 2520 3566 2527 3573 ne
rect 2527 3541 2535 3573
rect 2565 3541 2613 3583
rect 2643 3573 2668 3583
rect 2643 3541 2651 3573
rect 2767 3569 2792 3583
rect 2672 3541 2706 3569
rect 2736 3541 2792 3569
rect 2822 3541 2850 3583
rect 2908 3541 2936 3583
rect 2966 3569 2991 3583
rect 3090 3573 3115 3583
rect 2966 3541 3022 3569
rect 3052 3541 3086 3569
tri 3100 3566 3107 3573 ne
rect 3107 3541 3115 3573
rect 3145 3541 3193 3583
rect 3223 3573 3248 3583
rect 3223 3541 3231 3573
rect 3347 3569 3372 3583
rect 3252 3541 3286 3569
rect 3316 3541 3372 3569
rect 3402 3541 3430 3583
rect 3488 3541 3516 3583
rect 3546 3569 3571 3583
rect 3670 3573 3695 3583
rect 3546 3541 3602 3569
rect 3632 3541 3666 3569
tri 3680 3566 3687 3573 ne
rect 3687 3541 3695 3573
rect 3725 3541 3773 3583
rect 3803 3573 3828 3583
rect 3803 3541 3811 3573
rect 3927 3569 3952 3583
rect 3832 3541 3866 3569
rect 3896 3541 3952 3569
rect 3982 3541 4010 3583
rect 4068 3541 4096 3583
rect 4126 3569 4151 3583
rect 4250 3573 4275 3583
rect 4126 3541 4182 3569
rect 4212 3541 4246 3569
tri 4260 3566 4267 3573 ne
rect 4267 3541 4275 3573
rect 4305 3541 4353 3583
rect 4383 3573 4408 3583
rect 4383 3541 4391 3573
rect 4507 3569 4532 3583
rect 4412 3541 4446 3569
rect 4476 3541 4532 3569
rect 4562 3541 4590 3583
rect 4648 3541 4676 3583
rect 4706 3569 4731 3583
rect 4830 3573 4855 3583
rect 4706 3541 4762 3569
rect 4792 3541 4826 3569
tri 4840 3566 4847 3573 ne
rect 4847 3541 4855 3573
rect 4885 3541 4933 3583
rect 4963 3573 4988 3583
rect 4963 3541 4971 3573
rect 5087 3569 5112 3583
rect 4992 3541 5026 3569
rect 5056 3541 5112 3569
rect 5142 3541 5170 3583
rect 5228 3541 5256 3583
rect 5286 3569 5311 3583
rect 5410 3573 5435 3583
rect 5286 3541 5342 3569
rect 5372 3541 5406 3569
tri 5420 3566 5427 3573 ne
rect 5427 3541 5435 3573
rect 5465 3541 5513 3583
rect 5543 3573 5568 3583
rect 5543 3541 5551 3573
rect 5667 3569 5692 3583
rect 5572 3541 5606 3569
rect 5636 3541 5692 3569
rect 5722 3541 5750 3583
rect 5808 3541 5836 3583
rect 5866 3569 5891 3583
rect 5990 3573 6015 3583
rect 5866 3541 5922 3569
rect 5952 3541 5986 3569
tri 6000 3566 6007 3573 ne
rect 6007 3541 6015 3573
rect 6045 3541 6093 3583
rect 6123 3573 6148 3583
rect 6123 3541 6131 3573
rect 6247 3569 6272 3583
rect 6152 3541 6186 3569
rect 6216 3541 6272 3569
rect 6302 3541 6330 3583
rect 6388 3541 6416 3583
rect 6446 3569 6471 3583
rect 6570 3573 6595 3583
rect 6446 3541 6502 3569
rect 6532 3541 6566 3569
tri 6580 3566 6587 3573 ne
rect 6587 3541 6595 3573
rect 6625 3541 6673 3583
rect 6703 3573 6728 3583
rect 6703 3541 6711 3573
rect 6827 3569 6852 3583
rect 6732 3541 6766 3569
rect 6796 3541 6852 3569
rect 6882 3541 6910 3583
rect 159 3517 186 3541
rect 253 3519 285 3541
rect 253 3517 255 3519
rect 283 3517 285 3519
rect 352 3517 379 3541
rect 159 3503 253 3517
rect 285 3503 379 3517
rect 739 3517 766 3541
rect 833 3519 865 3541
rect 833 3517 835 3519
rect 863 3517 865 3519
rect 932 3517 959 3541
rect 739 3503 833 3517
rect 865 3503 959 3517
rect 1319 3517 1346 3541
rect 1413 3519 1445 3541
rect 1413 3517 1415 3519
rect 1443 3517 1445 3519
rect 1512 3517 1539 3541
rect 1319 3503 1413 3517
rect 1445 3503 1539 3517
rect 1899 3517 1926 3541
rect 1993 3519 2025 3541
rect 1993 3517 1995 3519
rect 2023 3517 2025 3519
rect 2092 3517 2119 3541
rect 1899 3503 1993 3517
rect 2025 3503 2119 3517
rect 2479 3517 2506 3541
rect 2573 3519 2605 3541
rect 2573 3517 2575 3519
rect 2603 3517 2605 3519
rect 2672 3517 2699 3541
rect 2479 3503 2573 3517
rect 2605 3503 2699 3517
rect 3059 3517 3086 3541
rect 3153 3519 3185 3541
rect 3153 3517 3155 3519
rect 3183 3517 3185 3519
rect 3252 3517 3279 3541
rect 3059 3503 3153 3517
rect 3185 3503 3279 3517
rect 3639 3517 3666 3541
rect 3733 3519 3765 3541
rect 3733 3517 3735 3519
rect 3763 3517 3765 3519
rect 3832 3517 3859 3541
rect 3639 3503 3733 3517
rect 3765 3503 3859 3517
rect 4219 3517 4246 3541
rect 4313 3519 4345 3541
rect 4313 3517 4315 3519
rect 4343 3517 4345 3519
rect 4412 3517 4439 3541
rect 4219 3503 4313 3517
rect 4345 3503 4439 3517
rect 4799 3517 4826 3541
rect 4893 3519 4925 3541
rect 4893 3517 4895 3519
rect 4923 3517 4925 3519
rect 4992 3517 5019 3541
rect 4799 3503 4893 3517
rect 4925 3503 5019 3517
rect 5379 3517 5406 3541
rect 5473 3519 5505 3541
rect 5473 3517 5475 3519
rect 5503 3517 5505 3519
rect 5572 3517 5599 3541
rect 5379 3503 5473 3517
rect 5505 3503 5599 3517
rect 5959 3517 5986 3541
rect 6053 3519 6085 3541
rect 6053 3517 6055 3519
rect 6083 3517 6085 3519
rect 6152 3517 6179 3541
rect 5959 3503 6053 3517
rect 6085 3503 6179 3517
rect 6539 3517 6566 3541
rect 6633 3519 6665 3541
rect 6633 3517 6635 3519
rect 6663 3517 6665 3519
rect 6732 3517 6759 3541
rect 6539 3503 6633 3517
rect 6665 3503 6759 3517
rect 82 3417 100 3445
rect 130 3417 148 3445
rect 390 3417 408 3445
rect 438 3417 457 3445
rect 662 3417 680 3445
rect 710 3417 728 3445
rect 970 3417 988 3445
rect 1018 3417 1037 3445
rect 1242 3417 1260 3445
rect 1290 3417 1308 3445
rect 1550 3417 1568 3445
rect 1598 3417 1617 3445
rect 1822 3417 1840 3445
rect 1870 3417 1888 3445
rect 2130 3417 2148 3445
rect 2178 3417 2197 3445
rect 2402 3417 2420 3445
rect 2450 3417 2468 3445
rect 2710 3417 2728 3445
rect 2758 3417 2777 3445
rect 2982 3417 3000 3445
rect 3030 3417 3048 3445
rect 3290 3417 3308 3445
rect 3338 3417 3357 3445
rect 3562 3417 3580 3445
rect 3610 3417 3628 3445
rect 3870 3417 3888 3445
rect 3918 3417 3937 3445
rect 4142 3417 4160 3445
rect 4190 3417 4208 3445
rect 4450 3417 4468 3445
rect 4498 3417 4517 3445
rect 4722 3417 4740 3445
rect 4770 3417 4788 3445
rect 5030 3417 5048 3445
rect 5078 3417 5097 3445
rect 5302 3417 5320 3445
rect 5350 3417 5368 3445
rect 5610 3417 5628 3445
rect 5658 3417 5677 3445
rect 5882 3417 5900 3445
rect 5930 3417 5948 3445
rect 6190 3417 6208 3445
rect 6238 3417 6257 3445
rect 6462 3417 6480 3445
rect 6510 3417 6528 3445
rect 6770 3417 6788 3445
rect 6818 3417 6837 3445
rect 8 3271 36 3313
rect 66 3299 91 3313
rect 190 3303 215 3313
rect 66 3271 122 3299
rect 152 3271 186 3299
tri 200 3296 207 3303 ne
rect 207 3271 215 3303
rect 245 3271 293 3313
rect 323 3303 348 3313
rect 323 3271 331 3303
rect 447 3299 472 3313
rect 352 3271 386 3299
rect 416 3271 472 3299
rect 502 3271 530 3313
rect 588 3271 616 3313
rect 646 3299 671 3313
rect 770 3303 795 3313
rect 646 3271 702 3299
rect 732 3271 766 3299
tri 780 3296 787 3303 ne
rect 787 3271 795 3303
rect 825 3271 873 3313
rect 903 3303 928 3313
rect 903 3271 911 3303
rect 1027 3299 1052 3313
rect 932 3271 966 3299
rect 996 3271 1052 3299
rect 1082 3271 1110 3313
rect 1168 3271 1196 3313
rect 1226 3299 1251 3313
rect 1350 3303 1375 3313
rect 1226 3271 1282 3299
rect 1312 3271 1346 3299
tri 1360 3296 1367 3303 ne
rect 1367 3271 1375 3303
rect 1405 3271 1453 3313
rect 1483 3303 1508 3313
rect 1483 3271 1491 3303
rect 1607 3299 1632 3313
rect 1512 3271 1546 3299
rect 1576 3271 1632 3299
rect 1662 3271 1690 3313
rect 1748 3271 1776 3313
rect 1806 3299 1831 3313
rect 1930 3303 1955 3313
rect 1806 3271 1862 3299
rect 1892 3271 1926 3299
tri 1940 3296 1947 3303 ne
rect 1947 3271 1955 3303
rect 1985 3271 2033 3313
rect 2063 3303 2088 3313
rect 2063 3271 2071 3303
rect 2187 3299 2212 3313
rect 2092 3271 2126 3299
rect 2156 3271 2212 3299
rect 2242 3271 2270 3313
rect 2328 3271 2356 3313
rect 2386 3299 2411 3313
rect 2510 3303 2535 3313
rect 2386 3271 2442 3299
rect 2472 3271 2506 3299
tri 2520 3296 2527 3303 ne
rect 2527 3271 2535 3303
rect 2565 3271 2613 3313
rect 2643 3303 2668 3313
rect 2643 3271 2651 3303
rect 2767 3299 2792 3313
rect 2672 3271 2706 3299
rect 2736 3271 2792 3299
rect 2822 3271 2850 3313
rect 2908 3271 2936 3313
rect 2966 3299 2991 3313
rect 3090 3303 3115 3313
rect 2966 3271 3022 3299
rect 3052 3271 3086 3299
tri 3100 3296 3107 3303 ne
rect 3107 3271 3115 3303
rect 3145 3271 3193 3313
rect 3223 3303 3248 3313
rect 3223 3271 3231 3303
rect 3347 3299 3372 3313
rect 3252 3271 3286 3299
rect 3316 3271 3372 3299
rect 3402 3271 3430 3313
rect 3488 3271 3516 3313
rect 3546 3299 3571 3313
rect 3670 3303 3695 3313
rect 3546 3271 3602 3299
rect 3632 3271 3666 3299
tri 3680 3296 3687 3303 ne
rect 3687 3271 3695 3303
rect 3725 3271 3773 3313
rect 3803 3303 3828 3313
rect 3803 3271 3811 3303
rect 3927 3299 3952 3313
rect 3832 3271 3866 3299
rect 3896 3271 3952 3299
rect 3982 3271 4010 3313
rect 4068 3271 4096 3313
rect 4126 3299 4151 3313
rect 4250 3303 4275 3313
rect 4126 3271 4182 3299
rect 4212 3271 4246 3299
tri 4260 3296 4267 3303 ne
rect 4267 3271 4275 3303
rect 4305 3271 4353 3313
rect 4383 3303 4408 3313
rect 4383 3271 4391 3303
rect 4507 3299 4532 3313
rect 4412 3271 4446 3299
rect 4476 3271 4532 3299
rect 4562 3271 4590 3313
rect 4648 3271 4676 3313
rect 4706 3299 4731 3313
rect 4830 3303 4855 3313
rect 4706 3271 4762 3299
rect 4792 3271 4826 3299
tri 4840 3296 4847 3303 ne
rect 4847 3271 4855 3303
rect 4885 3271 4933 3313
rect 4963 3303 4988 3313
rect 4963 3271 4971 3303
rect 5087 3299 5112 3313
rect 4992 3271 5026 3299
rect 5056 3271 5112 3299
rect 5142 3271 5170 3313
rect 5228 3271 5256 3313
rect 5286 3299 5311 3313
rect 5410 3303 5435 3313
rect 5286 3271 5342 3299
rect 5372 3271 5406 3299
tri 5420 3296 5427 3303 ne
rect 5427 3271 5435 3303
rect 5465 3271 5513 3313
rect 5543 3303 5568 3313
rect 5543 3271 5551 3303
rect 5667 3299 5692 3313
rect 5572 3271 5606 3299
rect 5636 3271 5692 3299
rect 5722 3271 5750 3313
rect 5808 3271 5836 3313
rect 5866 3299 5891 3313
rect 5990 3303 6015 3313
rect 5866 3271 5922 3299
rect 5952 3271 5986 3299
tri 6000 3296 6007 3303 ne
rect 6007 3271 6015 3303
rect 6045 3271 6093 3313
rect 6123 3303 6148 3313
rect 6123 3271 6131 3303
rect 6247 3299 6272 3313
rect 6152 3271 6186 3299
rect 6216 3271 6272 3299
rect 6302 3271 6330 3313
rect 6388 3271 6416 3313
rect 6446 3299 6471 3313
rect 6570 3303 6595 3313
rect 6446 3271 6502 3299
rect 6532 3271 6566 3299
tri 6580 3296 6587 3303 ne
rect 6587 3271 6595 3303
rect 6625 3271 6673 3313
rect 6703 3303 6728 3313
rect 6703 3271 6711 3303
rect 6827 3299 6852 3313
rect 6732 3271 6766 3299
rect 6796 3271 6852 3299
rect 6882 3271 6910 3313
rect 159 3247 186 3271
rect 253 3249 285 3271
rect 253 3247 255 3249
rect 283 3247 285 3249
rect 352 3247 379 3271
rect 159 3233 253 3247
rect 285 3233 379 3247
rect 739 3247 766 3271
rect 833 3249 865 3271
rect 833 3247 835 3249
rect 863 3247 865 3249
rect 932 3247 959 3271
rect 739 3233 833 3247
rect 865 3233 959 3247
rect 1319 3247 1346 3271
rect 1413 3249 1445 3271
rect 1413 3247 1415 3249
rect 1443 3247 1445 3249
rect 1512 3247 1539 3271
rect 1319 3233 1413 3247
rect 1445 3233 1539 3247
rect 1899 3247 1926 3271
rect 1993 3249 2025 3271
rect 1993 3247 1995 3249
rect 2023 3247 2025 3249
rect 2092 3247 2119 3271
rect 1899 3233 1993 3247
rect 2025 3233 2119 3247
rect 2479 3247 2506 3271
rect 2573 3249 2605 3271
rect 2573 3247 2575 3249
rect 2603 3247 2605 3249
rect 2672 3247 2699 3271
rect 2479 3233 2573 3247
rect 2605 3233 2699 3247
rect 3059 3247 3086 3271
rect 3153 3249 3185 3271
rect 3153 3247 3155 3249
rect 3183 3247 3185 3249
rect 3252 3247 3279 3271
rect 3059 3233 3153 3247
rect 3185 3233 3279 3247
rect 3639 3247 3666 3271
rect 3733 3249 3765 3271
rect 3733 3247 3735 3249
rect 3763 3247 3765 3249
rect 3832 3247 3859 3271
rect 3639 3233 3733 3247
rect 3765 3233 3859 3247
rect 4219 3247 4246 3271
rect 4313 3249 4345 3271
rect 4313 3247 4315 3249
rect 4343 3247 4345 3249
rect 4412 3247 4439 3271
rect 4219 3233 4313 3247
rect 4345 3233 4439 3247
rect 4799 3247 4826 3271
rect 4893 3249 4925 3271
rect 4893 3247 4895 3249
rect 4923 3247 4925 3249
rect 4992 3247 5019 3271
rect 4799 3233 4893 3247
rect 4925 3233 5019 3247
rect 5379 3247 5406 3271
rect 5473 3249 5505 3271
rect 5473 3247 5475 3249
rect 5503 3247 5505 3249
rect 5572 3247 5599 3271
rect 5379 3233 5473 3247
rect 5505 3233 5599 3247
rect 5959 3247 5986 3271
rect 6053 3249 6085 3271
rect 6053 3247 6055 3249
rect 6083 3247 6085 3249
rect 6152 3247 6179 3271
rect 5959 3233 6053 3247
rect 6085 3233 6179 3247
rect 6539 3247 6566 3271
rect 6633 3249 6665 3271
rect 6633 3247 6635 3249
rect 6663 3247 6665 3249
rect 6732 3247 6759 3271
rect 6539 3233 6633 3247
rect 6665 3233 6759 3247
rect 82 3147 100 3175
rect 130 3147 148 3175
rect 390 3147 408 3175
rect 438 3147 457 3175
rect 662 3147 680 3175
rect 710 3147 728 3175
rect 970 3147 988 3175
rect 1018 3147 1037 3175
rect 1242 3147 1260 3175
rect 1290 3147 1308 3175
rect 1550 3147 1568 3175
rect 1598 3147 1617 3175
rect 1822 3147 1840 3175
rect 1870 3147 1888 3175
rect 2130 3147 2148 3175
rect 2178 3147 2197 3175
rect 2402 3147 2420 3175
rect 2450 3147 2468 3175
rect 2710 3147 2728 3175
rect 2758 3147 2777 3175
rect 2982 3147 3000 3175
rect 3030 3147 3048 3175
rect 3290 3147 3308 3175
rect 3338 3147 3357 3175
rect 3562 3147 3580 3175
rect 3610 3147 3628 3175
rect 3870 3147 3888 3175
rect 3918 3147 3937 3175
rect 4142 3147 4160 3175
rect 4190 3147 4208 3175
rect 4450 3147 4468 3175
rect 4498 3147 4517 3175
rect 4722 3147 4740 3175
rect 4770 3147 4788 3175
rect 5030 3147 5048 3175
rect 5078 3147 5097 3175
rect 5302 3147 5320 3175
rect 5350 3147 5368 3175
rect 5610 3147 5628 3175
rect 5658 3147 5677 3175
rect 5882 3147 5900 3175
rect 5930 3147 5948 3175
rect 6190 3147 6208 3175
rect 6238 3147 6257 3175
rect 6462 3147 6480 3175
rect 6510 3147 6528 3175
rect 6770 3147 6788 3175
rect 6818 3147 6837 3175
rect 8 3001 36 3043
rect 66 3029 91 3043
rect 190 3033 215 3043
rect 66 3001 122 3029
rect 152 3001 186 3029
tri 200 3026 207 3033 ne
rect 207 3001 215 3033
rect 245 3001 293 3043
rect 323 3033 348 3043
rect 323 3001 331 3033
rect 447 3029 472 3043
rect 352 3001 386 3029
rect 416 3001 472 3029
rect 502 3001 530 3043
rect 588 3001 616 3043
rect 646 3029 671 3043
rect 770 3033 795 3043
rect 646 3001 702 3029
rect 732 3001 766 3029
tri 780 3026 787 3033 ne
rect 787 3001 795 3033
rect 825 3001 873 3043
rect 903 3033 928 3043
rect 903 3001 911 3033
rect 1027 3029 1052 3043
rect 932 3001 966 3029
rect 996 3001 1052 3029
rect 1082 3001 1110 3043
rect 1168 3001 1196 3043
rect 1226 3029 1251 3043
rect 1350 3033 1375 3043
rect 1226 3001 1282 3029
rect 1312 3001 1346 3029
tri 1360 3026 1367 3033 ne
rect 1367 3001 1375 3033
rect 1405 3001 1453 3043
rect 1483 3033 1508 3043
rect 1483 3001 1491 3033
rect 1607 3029 1632 3043
rect 1512 3001 1546 3029
rect 1576 3001 1632 3029
rect 1662 3001 1690 3043
rect 1748 3001 1776 3043
rect 1806 3029 1831 3043
rect 1930 3033 1955 3043
rect 1806 3001 1862 3029
rect 1892 3001 1926 3029
tri 1940 3026 1947 3033 ne
rect 1947 3001 1955 3033
rect 1985 3001 2033 3043
rect 2063 3033 2088 3043
rect 2063 3001 2071 3033
rect 2187 3029 2212 3043
rect 2092 3001 2126 3029
rect 2156 3001 2212 3029
rect 2242 3001 2270 3043
rect 2328 3001 2356 3043
rect 2386 3029 2411 3043
rect 2510 3033 2535 3043
rect 2386 3001 2442 3029
rect 2472 3001 2506 3029
tri 2520 3026 2527 3033 ne
rect 2527 3001 2535 3033
rect 2565 3001 2613 3043
rect 2643 3033 2668 3043
rect 2643 3001 2651 3033
rect 2767 3029 2792 3043
rect 2672 3001 2706 3029
rect 2736 3001 2792 3029
rect 2822 3001 2850 3043
rect 2908 3001 2936 3043
rect 2966 3029 2991 3043
rect 3090 3033 3115 3043
rect 2966 3001 3022 3029
rect 3052 3001 3086 3029
tri 3100 3026 3107 3033 ne
rect 3107 3001 3115 3033
rect 3145 3001 3193 3043
rect 3223 3033 3248 3043
rect 3223 3001 3231 3033
rect 3347 3029 3372 3043
rect 3252 3001 3286 3029
rect 3316 3001 3372 3029
rect 3402 3001 3430 3043
rect 3488 3001 3516 3043
rect 3546 3029 3571 3043
rect 3670 3033 3695 3043
rect 3546 3001 3602 3029
rect 3632 3001 3666 3029
tri 3680 3026 3687 3033 ne
rect 3687 3001 3695 3033
rect 3725 3001 3773 3043
rect 3803 3033 3828 3043
rect 3803 3001 3811 3033
rect 3927 3029 3952 3043
rect 3832 3001 3866 3029
rect 3896 3001 3952 3029
rect 3982 3001 4010 3043
rect 4068 3001 4096 3043
rect 4126 3029 4151 3043
rect 4250 3033 4275 3043
rect 4126 3001 4182 3029
rect 4212 3001 4246 3029
tri 4260 3026 4267 3033 ne
rect 4267 3001 4275 3033
rect 4305 3001 4353 3043
rect 4383 3033 4408 3043
rect 4383 3001 4391 3033
rect 4507 3029 4532 3043
rect 4412 3001 4446 3029
rect 4476 3001 4532 3029
rect 4562 3001 4590 3043
rect 4648 3001 4676 3043
rect 4706 3029 4731 3043
rect 4830 3033 4855 3043
rect 4706 3001 4762 3029
rect 4792 3001 4826 3029
tri 4840 3026 4847 3033 ne
rect 4847 3001 4855 3033
rect 4885 3001 4933 3043
rect 4963 3033 4988 3043
rect 4963 3001 4971 3033
rect 5087 3029 5112 3043
rect 4992 3001 5026 3029
rect 5056 3001 5112 3029
rect 5142 3001 5170 3043
rect 5228 3001 5256 3043
rect 5286 3029 5311 3043
rect 5410 3033 5435 3043
rect 5286 3001 5342 3029
rect 5372 3001 5406 3029
tri 5420 3026 5427 3033 ne
rect 5427 3001 5435 3033
rect 5465 3001 5513 3043
rect 5543 3033 5568 3043
rect 5543 3001 5551 3033
rect 5667 3029 5692 3043
rect 5572 3001 5606 3029
rect 5636 3001 5692 3029
rect 5722 3001 5750 3043
rect 5808 3001 5836 3043
rect 5866 3029 5891 3043
rect 5990 3033 6015 3043
rect 5866 3001 5922 3029
rect 5952 3001 5986 3029
tri 6000 3026 6007 3033 ne
rect 6007 3001 6015 3033
rect 6045 3001 6093 3043
rect 6123 3033 6148 3043
rect 6123 3001 6131 3033
rect 6247 3029 6272 3043
rect 6152 3001 6186 3029
rect 6216 3001 6272 3029
rect 6302 3001 6330 3043
rect 6388 3001 6416 3043
rect 6446 3029 6471 3043
rect 6570 3033 6595 3043
rect 6446 3001 6502 3029
rect 6532 3001 6566 3029
tri 6580 3026 6587 3033 ne
rect 6587 3001 6595 3033
rect 6625 3001 6673 3043
rect 6703 3033 6728 3043
rect 6703 3001 6711 3033
rect 6827 3029 6852 3043
rect 6732 3001 6766 3029
rect 6796 3001 6852 3029
rect 6882 3001 6910 3043
rect 159 2977 186 3001
rect 253 2979 285 3001
rect 253 2977 255 2979
rect 283 2977 285 2979
rect 352 2977 379 3001
rect 159 2963 253 2977
rect 285 2963 379 2977
rect 739 2977 766 3001
rect 833 2979 865 3001
rect 833 2977 835 2979
rect 863 2977 865 2979
rect 932 2977 959 3001
rect 739 2963 833 2977
rect 865 2963 959 2977
rect 1319 2977 1346 3001
rect 1413 2979 1445 3001
rect 1413 2977 1415 2979
rect 1443 2977 1445 2979
rect 1512 2977 1539 3001
rect 1319 2963 1413 2977
rect 1445 2963 1539 2977
rect 1899 2977 1926 3001
rect 1993 2979 2025 3001
rect 1993 2977 1995 2979
rect 2023 2977 2025 2979
rect 2092 2977 2119 3001
rect 1899 2963 1993 2977
rect 2025 2963 2119 2977
rect 2479 2977 2506 3001
rect 2573 2979 2605 3001
rect 2573 2977 2575 2979
rect 2603 2977 2605 2979
rect 2672 2977 2699 3001
rect 2479 2963 2573 2977
rect 2605 2963 2699 2977
rect 3059 2977 3086 3001
rect 3153 2979 3185 3001
rect 3153 2977 3155 2979
rect 3183 2977 3185 2979
rect 3252 2977 3279 3001
rect 3059 2963 3153 2977
rect 3185 2963 3279 2977
rect 3639 2977 3666 3001
rect 3733 2979 3765 3001
rect 3733 2977 3735 2979
rect 3763 2977 3765 2979
rect 3832 2977 3859 3001
rect 3639 2963 3733 2977
rect 3765 2963 3859 2977
rect 4219 2977 4246 3001
rect 4313 2979 4345 3001
rect 4313 2977 4315 2979
rect 4343 2977 4345 2979
rect 4412 2977 4439 3001
rect 4219 2963 4313 2977
rect 4345 2963 4439 2977
rect 4799 2977 4826 3001
rect 4893 2979 4925 3001
rect 4893 2977 4895 2979
rect 4923 2977 4925 2979
rect 4992 2977 5019 3001
rect 4799 2963 4893 2977
rect 4925 2963 5019 2977
rect 5379 2977 5406 3001
rect 5473 2979 5505 3001
rect 5473 2977 5475 2979
rect 5503 2977 5505 2979
rect 5572 2977 5599 3001
rect 5379 2963 5473 2977
rect 5505 2963 5599 2977
rect 5959 2977 5986 3001
rect 6053 2979 6085 3001
rect 6053 2977 6055 2979
rect 6083 2977 6085 2979
rect 6152 2977 6179 3001
rect 5959 2963 6053 2977
rect 6085 2963 6179 2977
rect 6539 2977 6566 3001
rect 6633 2979 6665 3001
rect 6633 2977 6635 2979
rect 6663 2977 6665 2979
rect 6732 2977 6759 3001
rect 6539 2963 6633 2977
rect 6665 2963 6759 2977
rect 82 2877 100 2905
rect 130 2877 148 2905
rect 390 2877 408 2905
rect 438 2877 457 2905
rect 662 2877 680 2905
rect 710 2877 728 2905
rect 970 2877 988 2905
rect 1018 2877 1037 2905
rect 1242 2877 1260 2905
rect 1290 2877 1308 2905
rect 1550 2877 1568 2905
rect 1598 2877 1617 2905
rect 1822 2877 1840 2905
rect 1870 2877 1888 2905
rect 2130 2877 2148 2905
rect 2178 2877 2197 2905
rect 2402 2877 2420 2905
rect 2450 2877 2468 2905
rect 2710 2877 2728 2905
rect 2758 2877 2777 2905
rect 2982 2877 3000 2905
rect 3030 2877 3048 2905
rect 3290 2877 3308 2905
rect 3338 2877 3357 2905
rect 3562 2877 3580 2905
rect 3610 2877 3628 2905
rect 3870 2877 3888 2905
rect 3918 2877 3937 2905
rect 4142 2877 4160 2905
rect 4190 2877 4208 2905
rect 4450 2877 4468 2905
rect 4498 2877 4517 2905
rect 4722 2877 4740 2905
rect 4770 2877 4788 2905
rect 5030 2877 5048 2905
rect 5078 2877 5097 2905
rect 5302 2877 5320 2905
rect 5350 2877 5368 2905
rect 5610 2877 5628 2905
rect 5658 2877 5677 2905
rect 5882 2877 5900 2905
rect 5930 2877 5948 2905
rect 6190 2877 6208 2905
rect 6238 2877 6257 2905
rect 6462 2877 6480 2905
rect 6510 2877 6528 2905
rect 6770 2877 6788 2905
rect 6818 2877 6837 2905
rect 8 2731 36 2773
rect 66 2759 91 2773
rect 190 2763 215 2773
rect 66 2731 122 2759
rect 152 2731 186 2759
tri 200 2756 207 2763 ne
rect 207 2731 215 2763
rect 245 2731 293 2773
rect 323 2763 348 2773
rect 323 2731 331 2763
rect 447 2759 472 2773
rect 352 2731 386 2759
rect 416 2731 472 2759
rect 502 2731 530 2773
rect 588 2731 616 2773
rect 646 2759 671 2773
rect 770 2763 795 2773
rect 646 2731 702 2759
rect 732 2731 766 2759
tri 780 2756 787 2763 ne
rect 787 2731 795 2763
rect 825 2731 873 2773
rect 903 2763 928 2773
rect 903 2731 911 2763
rect 1027 2759 1052 2773
rect 932 2731 966 2759
rect 996 2731 1052 2759
rect 1082 2731 1110 2773
rect 1168 2731 1196 2773
rect 1226 2759 1251 2773
rect 1350 2763 1375 2773
rect 1226 2731 1282 2759
rect 1312 2731 1346 2759
tri 1360 2756 1367 2763 ne
rect 1367 2731 1375 2763
rect 1405 2731 1453 2773
rect 1483 2763 1508 2773
rect 1483 2731 1491 2763
rect 1607 2759 1632 2773
rect 1512 2731 1546 2759
rect 1576 2731 1632 2759
rect 1662 2731 1690 2773
rect 1748 2731 1776 2773
rect 1806 2759 1831 2773
rect 1930 2763 1955 2773
rect 1806 2731 1862 2759
rect 1892 2731 1926 2759
tri 1940 2756 1947 2763 ne
rect 1947 2731 1955 2763
rect 1985 2731 2033 2773
rect 2063 2763 2088 2773
rect 2063 2731 2071 2763
rect 2187 2759 2212 2773
rect 2092 2731 2126 2759
rect 2156 2731 2212 2759
rect 2242 2731 2270 2773
rect 2328 2731 2356 2773
rect 2386 2759 2411 2773
rect 2510 2763 2535 2773
rect 2386 2731 2442 2759
rect 2472 2731 2506 2759
tri 2520 2756 2527 2763 ne
rect 2527 2731 2535 2763
rect 2565 2731 2613 2773
rect 2643 2763 2668 2773
rect 2643 2731 2651 2763
rect 2767 2759 2792 2773
rect 2672 2731 2706 2759
rect 2736 2731 2792 2759
rect 2822 2731 2850 2773
rect 2908 2731 2936 2773
rect 2966 2759 2991 2773
rect 3090 2763 3115 2773
rect 2966 2731 3022 2759
rect 3052 2731 3086 2759
tri 3100 2756 3107 2763 ne
rect 3107 2731 3115 2763
rect 3145 2731 3193 2773
rect 3223 2763 3248 2773
rect 3223 2731 3231 2763
rect 3347 2759 3372 2773
rect 3252 2731 3286 2759
rect 3316 2731 3372 2759
rect 3402 2731 3430 2773
rect 3488 2731 3516 2773
rect 3546 2759 3571 2773
rect 3670 2763 3695 2773
rect 3546 2731 3602 2759
rect 3632 2731 3666 2759
tri 3680 2756 3687 2763 ne
rect 3687 2731 3695 2763
rect 3725 2731 3773 2773
rect 3803 2763 3828 2773
rect 3803 2731 3811 2763
rect 3927 2759 3952 2773
rect 3832 2731 3866 2759
rect 3896 2731 3952 2759
rect 3982 2731 4010 2773
rect 4068 2731 4096 2773
rect 4126 2759 4151 2773
rect 4250 2763 4275 2773
rect 4126 2731 4182 2759
rect 4212 2731 4246 2759
tri 4260 2756 4267 2763 ne
rect 4267 2731 4275 2763
rect 4305 2731 4353 2773
rect 4383 2763 4408 2773
rect 4383 2731 4391 2763
rect 4507 2759 4532 2773
rect 4412 2731 4446 2759
rect 4476 2731 4532 2759
rect 4562 2731 4590 2773
rect 4648 2731 4676 2773
rect 4706 2759 4731 2773
rect 4830 2763 4855 2773
rect 4706 2731 4762 2759
rect 4792 2731 4826 2759
tri 4840 2756 4847 2763 ne
rect 4847 2731 4855 2763
rect 4885 2731 4933 2773
rect 4963 2763 4988 2773
rect 4963 2731 4971 2763
rect 5087 2759 5112 2773
rect 4992 2731 5026 2759
rect 5056 2731 5112 2759
rect 5142 2731 5170 2773
rect 5228 2731 5256 2773
rect 5286 2759 5311 2773
rect 5410 2763 5435 2773
rect 5286 2731 5342 2759
rect 5372 2731 5406 2759
tri 5420 2756 5427 2763 ne
rect 5427 2731 5435 2763
rect 5465 2731 5513 2773
rect 5543 2763 5568 2773
rect 5543 2731 5551 2763
rect 5667 2759 5692 2773
rect 5572 2731 5606 2759
rect 5636 2731 5692 2759
rect 5722 2731 5750 2773
rect 5808 2731 5836 2773
rect 5866 2759 5891 2773
rect 5990 2763 6015 2773
rect 5866 2731 5922 2759
rect 5952 2731 5986 2759
tri 6000 2756 6007 2763 ne
rect 6007 2731 6015 2763
rect 6045 2731 6093 2773
rect 6123 2763 6148 2773
rect 6123 2731 6131 2763
rect 6247 2759 6272 2773
rect 6152 2731 6186 2759
rect 6216 2731 6272 2759
rect 6302 2731 6330 2773
rect 6388 2731 6416 2773
rect 6446 2759 6471 2773
rect 6570 2763 6595 2773
rect 6446 2731 6502 2759
rect 6532 2731 6566 2759
tri 6580 2756 6587 2763 ne
rect 6587 2731 6595 2763
rect 6625 2731 6673 2773
rect 6703 2763 6728 2773
rect 6703 2731 6711 2763
rect 6827 2759 6852 2773
rect 6732 2731 6766 2759
rect 6796 2731 6852 2759
rect 6882 2731 6910 2773
rect 159 2707 186 2731
rect 253 2709 285 2731
rect 253 2707 255 2709
rect 283 2707 285 2709
rect 352 2707 379 2731
rect 159 2693 253 2707
rect 285 2693 379 2707
rect 739 2707 766 2731
rect 833 2709 865 2731
rect 833 2707 835 2709
rect 863 2707 865 2709
rect 932 2707 959 2731
rect 739 2693 833 2707
rect 865 2693 959 2707
rect 1319 2707 1346 2731
rect 1413 2709 1445 2731
rect 1413 2707 1415 2709
rect 1443 2707 1445 2709
rect 1512 2707 1539 2731
rect 1319 2693 1413 2707
rect 1445 2693 1539 2707
rect 1899 2707 1926 2731
rect 1993 2709 2025 2731
rect 1993 2707 1995 2709
rect 2023 2707 2025 2709
rect 2092 2707 2119 2731
rect 1899 2693 1993 2707
rect 2025 2693 2119 2707
rect 2479 2707 2506 2731
rect 2573 2709 2605 2731
rect 2573 2707 2575 2709
rect 2603 2707 2605 2709
rect 2672 2707 2699 2731
rect 2479 2693 2573 2707
rect 2605 2693 2699 2707
rect 3059 2707 3086 2731
rect 3153 2709 3185 2731
rect 3153 2707 3155 2709
rect 3183 2707 3185 2709
rect 3252 2707 3279 2731
rect 3059 2693 3153 2707
rect 3185 2693 3279 2707
rect 3639 2707 3666 2731
rect 3733 2709 3765 2731
rect 3733 2707 3735 2709
rect 3763 2707 3765 2709
rect 3832 2707 3859 2731
rect 3639 2693 3733 2707
rect 3765 2693 3859 2707
rect 4219 2707 4246 2731
rect 4313 2709 4345 2731
rect 4313 2707 4315 2709
rect 4343 2707 4345 2709
rect 4412 2707 4439 2731
rect 4219 2693 4313 2707
rect 4345 2693 4439 2707
rect 4799 2707 4826 2731
rect 4893 2709 4925 2731
rect 4893 2707 4895 2709
rect 4923 2707 4925 2709
rect 4992 2707 5019 2731
rect 4799 2693 4893 2707
rect 4925 2693 5019 2707
rect 5379 2707 5406 2731
rect 5473 2709 5505 2731
rect 5473 2707 5475 2709
rect 5503 2707 5505 2709
rect 5572 2707 5599 2731
rect 5379 2693 5473 2707
rect 5505 2693 5599 2707
rect 5959 2707 5986 2731
rect 6053 2709 6085 2731
rect 6053 2707 6055 2709
rect 6083 2707 6085 2709
rect 6152 2707 6179 2731
rect 5959 2693 6053 2707
rect 6085 2693 6179 2707
rect 6539 2707 6566 2731
rect 6633 2709 6665 2731
rect 6633 2707 6635 2709
rect 6663 2707 6665 2709
rect 6732 2707 6759 2731
rect 6539 2693 6633 2707
rect 6665 2693 6759 2707
rect 82 2607 100 2635
rect 130 2607 148 2635
rect 390 2607 408 2635
rect 438 2607 457 2635
rect 662 2607 680 2635
rect 710 2607 728 2635
rect 970 2607 988 2635
rect 1018 2607 1037 2635
rect 1242 2607 1260 2635
rect 1290 2607 1308 2635
rect 1550 2607 1568 2635
rect 1598 2607 1617 2635
rect 1822 2607 1840 2635
rect 1870 2607 1888 2635
rect 2130 2607 2148 2635
rect 2178 2607 2197 2635
rect 2402 2607 2420 2635
rect 2450 2607 2468 2635
rect 2710 2607 2728 2635
rect 2758 2607 2777 2635
rect 2982 2607 3000 2635
rect 3030 2607 3048 2635
rect 3290 2607 3308 2635
rect 3338 2607 3357 2635
rect 3562 2607 3580 2635
rect 3610 2607 3628 2635
rect 3870 2607 3888 2635
rect 3918 2607 3937 2635
rect 4142 2607 4160 2635
rect 4190 2607 4208 2635
rect 4450 2607 4468 2635
rect 4498 2607 4517 2635
rect 4722 2607 4740 2635
rect 4770 2607 4788 2635
rect 5030 2607 5048 2635
rect 5078 2607 5097 2635
rect 5302 2607 5320 2635
rect 5350 2607 5368 2635
rect 5610 2607 5628 2635
rect 5658 2607 5677 2635
rect 5882 2607 5900 2635
rect 5930 2607 5948 2635
rect 6190 2607 6208 2635
rect 6238 2607 6257 2635
rect 6462 2607 6480 2635
rect 6510 2607 6528 2635
rect 6770 2607 6788 2635
rect 6818 2607 6837 2635
rect 8 2461 36 2503
rect 66 2489 91 2503
rect 190 2493 215 2503
rect 66 2461 122 2489
rect 152 2461 186 2489
tri 200 2486 207 2493 ne
rect 207 2461 215 2493
rect 245 2461 293 2503
rect 323 2493 348 2503
rect 323 2461 331 2493
rect 447 2489 472 2503
rect 352 2461 386 2489
rect 416 2461 472 2489
rect 502 2461 530 2503
rect 588 2461 616 2503
rect 646 2489 671 2503
rect 770 2493 795 2503
rect 646 2461 702 2489
rect 732 2461 766 2489
tri 780 2486 787 2493 ne
rect 787 2461 795 2493
rect 825 2461 873 2503
rect 903 2493 928 2503
rect 903 2461 911 2493
rect 1027 2489 1052 2503
rect 932 2461 966 2489
rect 996 2461 1052 2489
rect 1082 2461 1110 2503
rect 1168 2461 1196 2503
rect 1226 2489 1251 2503
rect 1350 2493 1375 2503
rect 1226 2461 1282 2489
rect 1312 2461 1346 2489
tri 1360 2486 1367 2493 ne
rect 1367 2461 1375 2493
rect 1405 2461 1453 2503
rect 1483 2493 1508 2503
rect 1483 2461 1491 2493
rect 1607 2489 1632 2503
rect 1512 2461 1546 2489
rect 1576 2461 1632 2489
rect 1662 2461 1690 2503
rect 1748 2461 1776 2503
rect 1806 2489 1831 2503
rect 1930 2493 1955 2503
rect 1806 2461 1862 2489
rect 1892 2461 1926 2489
tri 1940 2486 1947 2493 ne
rect 1947 2461 1955 2493
rect 1985 2461 2033 2503
rect 2063 2493 2088 2503
rect 2063 2461 2071 2493
rect 2187 2489 2212 2503
rect 2092 2461 2126 2489
rect 2156 2461 2212 2489
rect 2242 2461 2270 2503
rect 2328 2461 2356 2503
rect 2386 2489 2411 2503
rect 2510 2493 2535 2503
rect 2386 2461 2442 2489
rect 2472 2461 2506 2489
tri 2520 2486 2527 2493 ne
rect 2527 2461 2535 2493
rect 2565 2461 2613 2503
rect 2643 2493 2668 2503
rect 2643 2461 2651 2493
rect 2767 2489 2792 2503
rect 2672 2461 2706 2489
rect 2736 2461 2792 2489
rect 2822 2461 2850 2503
rect 2908 2461 2936 2503
rect 2966 2489 2991 2503
rect 3090 2493 3115 2503
rect 2966 2461 3022 2489
rect 3052 2461 3086 2489
tri 3100 2486 3107 2493 ne
rect 3107 2461 3115 2493
rect 3145 2461 3193 2503
rect 3223 2493 3248 2503
rect 3223 2461 3231 2493
rect 3347 2489 3372 2503
rect 3252 2461 3286 2489
rect 3316 2461 3372 2489
rect 3402 2461 3430 2503
rect 3488 2461 3516 2503
rect 3546 2489 3571 2503
rect 3670 2493 3695 2503
rect 3546 2461 3602 2489
rect 3632 2461 3666 2489
tri 3680 2486 3687 2493 ne
rect 3687 2461 3695 2493
rect 3725 2461 3773 2503
rect 3803 2493 3828 2503
rect 3803 2461 3811 2493
rect 3927 2489 3952 2503
rect 3832 2461 3866 2489
rect 3896 2461 3952 2489
rect 3982 2461 4010 2503
rect 4068 2461 4096 2503
rect 4126 2489 4151 2503
rect 4250 2493 4275 2503
rect 4126 2461 4182 2489
rect 4212 2461 4246 2489
tri 4260 2486 4267 2493 ne
rect 4267 2461 4275 2493
rect 4305 2461 4353 2503
rect 4383 2493 4408 2503
rect 4383 2461 4391 2493
rect 4507 2489 4532 2503
rect 4412 2461 4446 2489
rect 4476 2461 4532 2489
rect 4562 2461 4590 2503
rect 4648 2461 4676 2503
rect 4706 2489 4731 2503
rect 4830 2493 4855 2503
rect 4706 2461 4762 2489
rect 4792 2461 4826 2489
tri 4840 2486 4847 2493 ne
rect 4847 2461 4855 2493
rect 4885 2461 4933 2503
rect 4963 2493 4988 2503
rect 4963 2461 4971 2493
rect 5087 2489 5112 2503
rect 4992 2461 5026 2489
rect 5056 2461 5112 2489
rect 5142 2461 5170 2503
rect 5228 2461 5256 2503
rect 5286 2489 5311 2503
rect 5410 2493 5435 2503
rect 5286 2461 5342 2489
rect 5372 2461 5406 2489
tri 5420 2486 5427 2493 ne
rect 5427 2461 5435 2493
rect 5465 2461 5513 2503
rect 5543 2493 5568 2503
rect 5543 2461 5551 2493
rect 5667 2489 5692 2503
rect 5572 2461 5606 2489
rect 5636 2461 5692 2489
rect 5722 2461 5750 2503
rect 5808 2461 5836 2503
rect 5866 2489 5891 2503
rect 5990 2493 6015 2503
rect 5866 2461 5922 2489
rect 5952 2461 5986 2489
tri 6000 2486 6007 2493 ne
rect 6007 2461 6015 2493
rect 6045 2461 6093 2503
rect 6123 2493 6148 2503
rect 6123 2461 6131 2493
rect 6247 2489 6272 2503
rect 6152 2461 6186 2489
rect 6216 2461 6272 2489
rect 6302 2461 6330 2503
rect 6388 2461 6416 2503
rect 6446 2489 6471 2503
rect 6570 2493 6595 2503
rect 6446 2461 6502 2489
rect 6532 2461 6566 2489
tri 6580 2486 6587 2493 ne
rect 6587 2461 6595 2493
rect 6625 2461 6673 2503
rect 6703 2493 6728 2503
rect 6703 2461 6711 2493
rect 6827 2489 6852 2503
rect 6732 2461 6766 2489
rect 6796 2461 6852 2489
rect 6882 2461 6910 2503
rect 159 2437 186 2461
rect 253 2439 285 2461
rect 253 2437 255 2439
rect 283 2437 285 2439
rect 352 2437 379 2461
rect 159 2423 253 2437
rect 285 2423 379 2437
rect 739 2437 766 2461
rect 833 2439 865 2461
rect 833 2437 835 2439
rect 863 2437 865 2439
rect 932 2437 959 2461
rect 739 2423 833 2437
rect 865 2423 959 2437
rect 1319 2437 1346 2461
rect 1413 2439 1445 2461
rect 1413 2437 1415 2439
rect 1443 2437 1445 2439
rect 1512 2437 1539 2461
rect 1319 2423 1413 2437
rect 1445 2423 1539 2437
rect 1899 2437 1926 2461
rect 1993 2439 2025 2461
rect 1993 2437 1995 2439
rect 2023 2437 2025 2439
rect 2092 2437 2119 2461
rect 1899 2423 1993 2437
rect 2025 2423 2119 2437
rect 2479 2437 2506 2461
rect 2573 2439 2605 2461
rect 2573 2437 2575 2439
rect 2603 2437 2605 2439
rect 2672 2437 2699 2461
rect 2479 2423 2573 2437
rect 2605 2423 2699 2437
rect 3059 2437 3086 2461
rect 3153 2439 3185 2461
rect 3153 2437 3155 2439
rect 3183 2437 3185 2439
rect 3252 2437 3279 2461
rect 3059 2423 3153 2437
rect 3185 2423 3279 2437
rect 3639 2437 3666 2461
rect 3733 2439 3765 2461
rect 3733 2437 3735 2439
rect 3763 2437 3765 2439
rect 3832 2437 3859 2461
rect 3639 2423 3733 2437
rect 3765 2423 3859 2437
rect 4219 2437 4246 2461
rect 4313 2439 4345 2461
rect 4313 2437 4315 2439
rect 4343 2437 4345 2439
rect 4412 2437 4439 2461
rect 4219 2423 4313 2437
rect 4345 2423 4439 2437
rect 4799 2437 4826 2461
rect 4893 2439 4925 2461
rect 4893 2437 4895 2439
rect 4923 2437 4925 2439
rect 4992 2437 5019 2461
rect 4799 2423 4893 2437
rect 4925 2423 5019 2437
rect 5379 2437 5406 2461
rect 5473 2439 5505 2461
rect 5473 2437 5475 2439
rect 5503 2437 5505 2439
rect 5572 2437 5599 2461
rect 5379 2423 5473 2437
rect 5505 2423 5599 2437
rect 5959 2437 5986 2461
rect 6053 2439 6085 2461
rect 6053 2437 6055 2439
rect 6083 2437 6085 2439
rect 6152 2437 6179 2461
rect 5959 2423 6053 2437
rect 6085 2423 6179 2437
rect 6539 2437 6566 2461
rect 6633 2439 6665 2461
rect 6633 2437 6635 2439
rect 6663 2437 6665 2439
rect 6732 2437 6759 2461
rect 6539 2423 6633 2437
rect 6665 2423 6759 2437
rect 82 2337 100 2365
rect 130 2337 148 2365
rect 390 2337 408 2365
rect 438 2337 457 2365
rect 662 2337 680 2365
rect 710 2337 728 2365
rect 970 2337 988 2365
rect 1018 2337 1037 2365
rect 1242 2337 1260 2365
rect 1290 2337 1308 2365
rect 1550 2337 1568 2365
rect 1598 2337 1617 2365
rect 1822 2337 1840 2365
rect 1870 2337 1888 2365
rect 2130 2337 2148 2365
rect 2178 2337 2197 2365
rect 2402 2337 2420 2365
rect 2450 2337 2468 2365
rect 2710 2337 2728 2365
rect 2758 2337 2777 2365
rect 2982 2337 3000 2365
rect 3030 2337 3048 2365
rect 3290 2337 3308 2365
rect 3338 2337 3357 2365
rect 3562 2337 3580 2365
rect 3610 2337 3628 2365
rect 3870 2337 3888 2365
rect 3918 2337 3937 2365
rect 4142 2337 4160 2365
rect 4190 2337 4208 2365
rect 4450 2337 4468 2365
rect 4498 2337 4517 2365
rect 4722 2337 4740 2365
rect 4770 2337 4788 2365
rect 5030 2337 5048 2365
rect 5078 2337 5097 2365
rect 5302 2337 5320 2365
rect 5350 2337 5368 2365
rect 5610 2337 5628 2365
rect 5658 2337 5677 2365
rect 5882 2337 5900 2365
rect 5930 2337 5948 2365
rect 6190 2337 6208 2365
rect 6238 2337 6257 2365
rect 6462 2337 6480 2365
rect 6510 2337 6528 2365
rect 6770 2337 6788 2365
rect 6818 2337 6837 2365
rect 8 2191 36 2233
rect 66 2219 91 2233
rect 190 2223 215 2233
rect 66 2191 122 2219
rect 152 2191 186 2219
tri 200 2216 207 2223 ne
rect 207 2191 215 2223
rect 245 2191 293 2233
rect 323 2223 348 2233
rect 323 2191 331 2223
rect 447 2219 472 2233
rect 352 2191 386 2219
rect 416 2191 472 2219
rect 502 2191 530 2233
rect 588 2191 616 2233
rect 646 2219 671 2233
rect 770 2223 795 2233
rect 646 2191 702 2219
rect 732 2191 766 2219
tri 780 2216 787 2223 ne
rect 787 2191 795 2223
rect 825 2191 873 2233
rect 903 2223 928 2233
rect 903 2191 911 2223
rect 1027 2219 1052 2233
rect 932 2191 966 2219
rect 996 2191 1052 2219
rect 1082 2191 1110 2233
rect 1168 2191 1196 2233
rect 1226 2219 1251 2233
rect 1350 2223 1375 2233
rect 1226 2191 1282 2219
rect 1312 2191 1346 2219
tri 1360 2216 1367 2223 ne
rect 1367 2191 1375 2223
rect 1405 2191 1453 2233
rect 1483 2223 1508 2233
rect 1483 2191 1491 2223
rect 1607 2219 1632 2233
rect 1512 2191 1546 2219
rect 1576 2191 1632 2219
rect 1662 2191 1690 2233
rect 1748 2191 1776 2233
rect 1806 2219 1831 2233
rect 1930 2223 1955 2233
rect 1806 2191 1862 2219
rect 1892 2191 1926 2219
tri 1940 2216 1947 2223 ne
rect 1947 2191 1955 2223
rect 1985 2191 2033 2233
rect 2063 2223 2088 2233
rect 2063 2191 2071 2223
rect 2187 2219 2212 2233
rect 2092 2191 2126 2219
rect 2156 2191 2212 2219
rect 2242 2191 2270 2233
rect 2328 2191 2356 2233
rect 2386 2219 2411 2233
rect 2510 2223 2535 2233
rect 2386 2191 2442 2219
rect 2472 2191 2506 2219
tri 2520 2216 2527 2223 ne
rect 2527 2191 2535 2223
rect 2565 2191 2613 2233
rect 2643 2223 2668 2233
rect 2643 2191 2651 2223
rect 2767 2219 2792 2233
rect 2672 2191 2706 2219
rect 2736 2191 2792 2219
rect 2822 2191 2850 2233
rect 2908 2191 2936 2233
rect 2966 2219 2991 2233
rect 3090 2223 3115 2233
rect 2966 2191 3022 2219
rect 3052 2191 3086 2219
tri 3100 2216 3107 2223 ne
rect 3107 2191 3115 2223
rect 3145 2191 3193 2233
rect 3223 2223 3248 2233
rect 3223 2191 3231 2223
rect 3347 2219 3372 2233
rect 3252 2191 3286 2219
rect 3316 2191 3372 2219
rect 3402 2191 3430 2233
rect 3488 2191 3516 2233
rect 3546 2219 3571 2233
rect 3670 2223 3695 2233
rect 3546 2191 3602 2219
rect 3632 2191 3666 2219
tri 3680 2216 3687 2223 ne
rect 3687 2191 3695 2223
rect 3725 2191 3773 2233
rect 3803 2223 3828 2233
rect 3803 2191 3811 2223
rect 3927 2219 3952 2233
rect 3832 2191 3866 2219
rect 3896 2191 3952 2219
rect 3982 2191 4010 2233
rect 4068 2191 4096 2233
rect 4126 2219 4151 2233
rect 4250 2223 4275 2233
rect 4126 2191 4182 2219
rect 4212 2191 4246 2219
tri 4260 2216 4267 2223 ne
rect 4267 2191 4275 2223
rect 4305 2191 4353 2233
rect 4383 2223 4408 2233
rect 4383 2191 4391 2223
rect 4507 2219 4532 2233
rect 4412 2191 4446 2219
rect 4476 2191 4532 2219
rect 4562 2191 4590 2233
rect 4648 2191 4676 2233
rect 4706 2219 4731 2233
rect 4830 2223 4855 2233
rect 4706 2191 4762 2219
rect 4792 2191 4826 2219
tri 4840 2216 4847 2223 ne
rect 4847 2191 4855 2223
rect 4885 2191 4933 2233
rect 4963 2223 4988 2233
rect 4963 2191 4971 2223
rect 5087 2219 5112 2233
rect 4992 2191 5026 2219
rect 5056 2191 5112 2219
rect 5142 2191 5170 2233
rect 5228 2191 5256 2233
rect 5286 2219 5311 2233
rect 5410 2223 5435 2233
rect 5286 2191 5342 2219
rect 5372 2191 5406 2219
tri 5420 2216 5427 2223 ne
rect 5427 2191 5435 2223
rect 5465 2191 5513 2233
rect 5543 2223 5568 2233
rect 5543 2191 5551 2223
rect 5667 2219 5692 2233
rect 5572 2191 5606 2219
rect 5636 2191 5692 2219
rect 5722 2191 5750 2233
rect 5808 2191 5836 2233
rect 5866 2219 5891 2233
rect 5990 2223 6015 2233
rect 5866 2191 5922 2219
rect 5952 2191 5986 2219
tri 6000 2216 6007 2223 ne
rect 6007 2191 6015 2223
rect 6045 2191 6093 2233
rect 6123 2223 6148 2233
rect 6123 2191 6131 2223
rect 6247 2219 6272 2233
rect 6152 2191 6186 2219
rect 6216 2191 6272 2219
rect 6302 2191 6330 2233
rect 6388 2191 6416 2233
rect 6446 2219 6471 2233
rect 6570 2223 6595 2233
rect 6446 2191 6502 2219
rect 6532 2191 6566 2219
tri 6580 2216 6587 2223 ne
rect 6587 2191 6595 2223
rect 6625 2191 6673 2233
rect 6703 2223 6728 2233
rect 6703 2191 6711 2223
rect 6827 2219 6852 2233
rect 6732 2191 6766 2219
rect 6796 2191 6852 2219
rect 6882 2191 6910 2233
rect 159 2167 186 2191
rect 253 2169 285 2191
rect 253 2167 255 2169
rect 283 2167 285 2169
rect 352 2167 379 2191
rect 159 2153 253 2167
rect 285 2153 379 2167
rect 739 2167 766 2191
rect 833 2169 865 2191
rect 833 2167 835 2169
rect 863 2167 865 2169
rect 932 2167 959 2191
rect 739 2153 833 2167
rect 865 2153 959 2167
rect 1319 2167 1346 2191
rect 1413 2169 1445 2191
rect 1413 2167 1415 2169
rect 1443 2167 1445 2169
rect 1512 2167 1539 2191
rect 1319 2153 1413 2167
rect 1445 2153 1539 2167
rect 1899 2167 1926 2191
rect 1993 2169 2025 2191
rect 1993 2167 1995 2169
rect 2023 2167 2025 2169
rect 2092 2167 2119 2191
rect 1899 2153 1993 2167
rect 2025 2153 2119 2167
rect 2479 2167 2506 2191
rect 2573 2169 2605 2191
rect 2573 2167 2575 2169
rect 2603 2167 2605 2169
rect 2672 2167 2699 2191
rect 2479 2153 2573 2167
rect 2605 2153 2699 2167
rect 3059 2167 3086 2191
rect 3153 2169 3185 2191
rect 3153 2167 3155 2169
rect 3183 2167 3185 2169
rect 3252 2167 3279 2191
rect 3059 2153 3153 2167
rect 3185 2153 3279 2167
rect 3639 2167 3666 2191
rect 3733 2169 3765 2191
rect 3733 2167 3735 2169
rect 3763 2167 3765 2169
rect 3832 2167 3859 2191
rect 3639 2153 3733 2167
rect 3765 2153 3859 2167
rect 4219 2167 4246 2191
rect 4313 2169 4345 2191
rect 4313 2167 4315 2169
rect 4343 2167 4345 2169
rect 4412 2167 4439 2191
rect 4219 2153 4313 2167
rect 4345 2153 4439 2167
rect 4799 2167 4826 2191
rect 4893 2169 4925 2191
rect 4893 2167 4895 2169
rect 4923 2167 4925 2169
rect 4992 2167 5019 2191
rect 4799 2153 4893 2167
rect 4925 2153 5019 2167
rect 5379 2167 5406 2191
rect 5473 2169 5505 2191
rect 5473 2167 5475 2169
rect 5503 2167 5505 2169
rect 5572 2167 5599 2191
rect 5379 2153 5473 2167
rect 5505 2153 5599 2167
rect 5959 2167 5986 2191
rect 6053 2169 6085 2191
rect 6053 2167 6055 2169
rect 6083 2167 6085 2169
rect 6152 2167 6179 2191
rect 5959 2153 6053 2167
rect 6085 2153 6179 2167
rect 6539 2167 6566 2191
rect 6633 2169 6665 2191
rect 6633 2167 6635 2169
rect 6663 2167 6665 2169
rect 6732 2167 6759 2191
rect 6539 2153 6633 2167
rect 6665 2153 6759 2167
rect 82 2067 100 2095
rect 130 2067 148 2095
rect 390 2067 408 2095
rect 438 2067 457 2095
rect 662 2067 680 2095
rect 710 2067 728 2095
rect 970 2067 988 2095
rect 1018 2067 1037 2095
rect 1242 2067 1260 2095
rect 1290 2067 1308 2095
rect 1550 2067 1568 2095
rect 1598 2067 1617 2095
rect 1822 2067 1840 2095
rect 1870 2067 1888 2095
rect 2130 2067 2148 2095
rect 2178 2067 2197 2095
rect 2402 2067 2420 2095
rect 2450 2067 2468 2095
rect 2710 2067 2728 2095
rect 2758 2067 2777 2095
rect 2982 2067 3000 2095
rect 3030 2067 3048 2095
rect 3290 2067 3308 2095
rect 3338 2067 3357 2095
rect 3562 2067 3580 2095
rect 3610 2067 3628 2095
rect 3870 2067 3888 2095
rect 3918 2067 3937 2095
rect 4142 2067 4160 2095
rect 4190 2067 4208 2095
rect 4450 2067 4468 2095
rect 4498 2067 4517 2095
rect 4722 2067 4740 2095
rect 4770 2067 4788 2095
rect 5030 2067 5048 2095
rect 5078 2067 5097 2095
rect 5302 2067 5320 2095
rect 5350 2067 5368 2095
rect 5610 2067 5628 2095
rect 5658 2067 5677 2095
rect 5882 2067 5900 2095
rect 5930 2067 5948 2095
rect 6190 2067 6208 2095
rect 6238 2067 6257 2095
rect 6462 2067 6480 2095
rect 6510 2067 6528 2095
rect 6770 2067 6788 2095
rect 6818 2067 6837 2095
rect 8 1921 36 1963
rect 66 1949 91 1963
rect 190 1953 215 1963
rect 66 1921 122 1949
rect 152 1921 186 1949
tri 200 1946 207 1953 ne
rect 207 1921 215 1953
rect 245 1921 293 1963
rect 323 1953 348 1963
rect 323 1921 331 1953
rect 447 1949 472 1963
rect 352 1921 386 1949
rect 416 1921 472 1949
rect 502 1921 530 1963
rect 588 1921 616 1963
rect 646 1949 671 1963
rect 770 1953 795 1963
rect 646 1921 702 1949
rect 732 1921 766 1949
tri 780 1946 787 1953 ne
rect 787 1921 795 1953
rect 825 1921 873 1963
rect 903 1953 928 1963
rect 903 1921 911 1953
rect 1027 1949 1052 1963
rect 932 1921 966 1949
rect 996 1921 1052 1949
rect 1082 1921 1110 1963
rect 1168 1921 1196 1963
rect 1226 1949 1251 1963
rect 1350 1953 1375 1963
rect 1226 1921 1282 1949
rect 1312 1921 1346 1949
tri 1360 1946 1367 1953 ne
rect 1367 1921 1375 1953
rect 1405 1921 1453 1963
rect 1483 1953 1508 1963
rect 1483 1921 1491 1953
rect 1607 1949 1632 1963
rect 1512 1921 1546 1949
rect 1576 1921 1632 1949
rect 1662 1921 1690 1963
rect 1748 1921 1776 1963
rect 1806 1949 1831 1963
rect 1930 1953 1955 1963
rect 1806 1921 1862 1949
rect 1892 1921 1926 1949
tri 1940 1946 1947 1953 ne
rect 1947 1921 1955 1953
rect 1985 1921 2033 1963
rect 2063 1953 2088 1963
rect 2063 1921 2071 1953
rect 2187 1949 2212 1963
rect 2092 1921 2126 1949
rect 2156 1921 2212 1949
rect 2242 1921 2270 1963
rect 2328 1921 2356 1963
rect 2386 1949 2411 1963
rect 2510 1953 2535 1963
rect 2386 1921 2442 1949
rect 2472 1921 2506 1949
tri 2520 1946 2527 1953 ne
rect 2527 1921 2535 1953
rect 2565 1921 2613 1963
rect 2643 1953 2668 1963
rect 2643 1921 2651 1953
rect 2767 1949 2792 1963
rect 2672 1921 2706 1949
rect 2736 1921 2792 1949
rect 2822 1921 2850 1963
rect 2908 1921 2936 1963
rect 2966 1949 2991 1963
rect 3090 1953 3115 1963
rect 2966 1921 3022 1949
rect 3052 1921 3086 1949
tri 3100 1946 3107 1953 ne
rect 3107 1921 3115 1953
rect 3145 1921 3193 1963
rect 3223 1953 3248 1963
rect 3223 1921 3231 1953
rect 3347 1949 3372 1963
rect 3252 1921 3286 1949
rect 3316 1921 3372 1949
rect 3402 1921 3430 1963
rect 3488 1921 3516 1963
rect 3546 1949 3571 1963
rect 3670 1953 3695 1963
rect 3546 1921 3602 1949
rect 3632 1921 3666 1949
tri 3680 1946 3687 1953 ne
rect 3687 1921 3695 1953
rect 3725 1921 3773 1963
rect 3803 1953 3828 1963
rect 3803 1921 3811 1953
rect 3927 1949 3952 1963
rect 3832 1921 3866 1949
rect 3896 1921 3952 1949
rect 3982 1921 4010 1963
rect 4068 1921 4096 1963
rect 4126 1949 4151 1963
rect 4250 1953 4275 1963
rect 4126 1921 4182 1949
rect 4212 1921 4246 1949
tri 4260 1946 4267 1953 ne
rect 4267 1921 4275 1953
rect 4305 1921 4353 1963
rect 4383 1953 4408 1963
rect 4383 1921 4391 1953
rect 4507 1949 4532 1963
rect 4412 1921 4446 1949
rect 4476 1921 4532 1949
rect 4562 1921 4590 1963
rect 4648 1921 4676 1963
rect 4706 1949 4731 1963
rect 4830 1953 4855 1963
rect 4706 1921 4762 1949
rect 4792 1921 4826 1949
tri 4840 1946 4847 1953 ne
rect 4847 1921 4855 1953
rect 4885 1921 4933 1963
rect 4963 1953 4988 1963
rect 4963 1921 4971 1953
rect 5087 1949 5112 1963
rect 4992 1921 5026 1949
rect 5056 1921 5112 1949
rect 5142 1921 5170 1963
rect 5228 1921 5256 1963
rect 5286 1949 5311 1963
rect 5410 1953 5435 1963
rect 5286 1921 5342 1949
rect 5372 1921 5406 1949
tri 5420 1946 5427 1953 ne
rect 5427 1921 5435 1953
rect 5465 1921 5513 1963
rect 5543 1953 5568 1963
rect 5543 1921 5551 1953
rect 5667 1949 5692 1963
rect 5572 1921 5606 1949
rect 5636 1921 5692 1949
rect 5722 1921 5750 1963
rect 5808 1921 5836 1963
rect 5866 1949 5891 1963
rect 5990 1953 6015 1963
rect 5866 1921 5922 1949
rect 5952 1921 5986 1949
tri 6000 1946 6007 1953 ne
rect 6007 1921 6015 1953
rect 6045 1921 6093 1963
rect 6123 1953 6148 1963
rect 6123 1921 6131 1953
rect 6247 1949 6272 1963
rect 6152 1921 6186 1949
rect 6216 1921 6272 1949
rect 6302 1921 6330 1963
rect 6388 1921 6416 1963
rect 6446 1949 6471 1963
rect 6570 1953 6595 1963
rect 6446 1921 6502 1949
rect 6532 1921 6566 1949
tri 6580 1946 6587 1953 ne
rect 6587 1921 6595 1953
rect 6625 1921 6673 1963
rect 6703 1953 6728 1963
rect 6703 1921 6711 1953
rect 6827 1949 6852 1963
rect 6732 1921 6766 1949
rect 6796 1921 6852 1949
rect 6882 1921 6910 1963
rect 159 1897 186 1921
rect 253 1899 285 1921
rect 253 1897 255 1899
rect 283 1897 285 1899
rect 352 1897 379 1921
rect 159 1883 253 1897
rect 285 1883 379 1897
rect 739 1897 766 1921
rect 833 1899 865 1921
rect 833 1897 835 1899
rect 863 1897 865 1899
rect 932 1897 959 1921
rect 739 1883 833 1897
rect 865 1883 959 1897
rect 1319 1897 1346 1921
rect 1413 1899 1445 1921
rect 1413 1897 1415 1899
rect 1443 1897 1445 1899
rect 1512 1897 1539 1921
rect 1319 1883 1413 1897
rect 1445 1883 1539 1897
rect 1899 1897 1926 1921
rect 1993 1899 2025 1921
rect 1993 1897 1995 1899
rect 2023 1897 2025 1899
rect 2092 1897 2119 1921
rect 1899 1883 1993 1897
rect 2025 1883 2119 1897
rect 2479 1897 2506 1921
rect 2573 1899 2605 1921
rect 2573 1897 2575 1899
rect 2603 1897 2605 1899
rect 2672 1897 2699 1921
rect 2479 1883 2573 1897
rect 2605 1883 2699 1897
rect 3059 1897 3086 1921
rect 3153 1899 3185 1921
rect 3153 1897 3155 1899
rect 3183 1897 3185 1899
rect 3252 1897 3279 1921
rect 3059 1883 3153 1897
rect 3185 1883 3279 1897
rect 3639 1897 3666 1921
rect 3733 1899 3765 1921
rect 3733 1897 3735 1899
rect 3763 1897 3765 1899
rect 3832 1897 3859 1921
rect 3639 1883 3733 1897
rect 3765 1883 3859 1897
rect 4219 1897 4246 1921
rect 4313 1899 4345 1921
rect 4313 1897 4315 1899
rect 4343 1897 4345 1899
rect 4412 1897 4439 1921
rect 4219 1883 4313 1897
rect 4345 1883 4439 1897
rect 4799 1897 4826 1921
rect 4893 1899 4925 1921
rect 4893 1897 4895 1899
rect 4923 1897 4925 1899
rect 4992 1897 5019 1921
rect 4799 1883 4893 1897
rect 4925 1883 5019 1897
rect 5379 1897 5406 1921
rect 5473 1899 5505 1921
rect 5473 1897 5475 1899
rect 5503 1897 5505 1899
rect 5572 1897 5599 1921
rect 5379 1883 5473 1897
rect 5505 1883 5599 1897
rect 5959 1897 5986 1921
rect 6053 1899 6085 1921
rect 6053 1897 6055 1899
rect 6083 1897 6085 1899
rect 6152 1897 6179 1921
rect 5959 1883 6053 1897
rect 6085 1883 6179 1897
rect 6539 1897 6566 1921
rect 6633 1899 6665 1921
rect 6633 1897 6635 1899
rect 6663 1897 6665 1899
rect 6732 1897 6759 1921
rect 6539 1883 6633 1897
rect 6665 1883 6759 1897
rect 82 1797 100 1825
rect 130 1797 148 1825
rect 390 1797 408 1825
rect 438 1797 457 1825
rect 662 1797 680 1825
rect 710 1797 728 1825
rect 970 1797 988 1825
rect 1018 1797 1037 1825
rect 1242 1797 1260 1825
rect 1290 1797 1308 1825
rect 1550 1797 1568 1825
rect 1598 1797 1617 1825
rect 1822 1797 1840 1825
rect 1870 1797 1888 1825
rect 2130 1797 2148 1825
rect 2178 1797 2197 1825
rect 2402 1797 2420 1825
rect 2450 1797 2468 1825
rect 2710 1797 2728 1825
rect 2758 1797 2777 1825
rect 2982 1797 3000 1825
rect 3030 1797 3048 1825
rect 3290 1797 3308 1825
rect 3338 1797 3357 1825
rect 3562 1797 3580 1825
rect 3610 1797 3628 1825
rect 3870 1797 3888 1825
rect 3918 1797 3937 1825
rect 4142 1797 4160 1825
rect 4190 1797 4208 1825
rect 4450 1797 4468 1825
rect 4498 1797 4517 1825
rect 4722 1797 4740 1825
rect 4770 1797 4788 1825
rect 5030 1797 5048 1825
rect 5078 1797 5097 1825
rect 5302 1797 5320 1825
rect 5350 1797 5368 1825
rect 5610 1797 5628 1825
rect 5658 1797 5677 1825
rect 5882 1797 5900 1825
rect 5930 1797 5948 1825
rect 6190 1797 6208 1825
rect 6238 1797 6257 1825
rect 6462 1797 6480 1825
rect 6510 1797 6528 1825
rect 6770 1797 6788 1825
rect 6818 1797 6837 1825
rect 8 1651 36 1693
rect 66 1679 91 1693
rect 190 1683 215 1693
rect 66 1651 122 1679
rect 152 1651 186 1679
tri 200 1676 207 1683 ne
rect 207 1651 215 1683
rect 245 1651 293 1693
rect 323 1683 348 1693
rect 323 1651 331 1683
rect 447 1679 472 1693
rect 352 1651 386 1679
rect 416 1651 472 1679
rect 502 1651 530 1693
rect 588 1651 616 1693
rect 646 1679 671 1693
rect 770 1683 795 1693
rect 646 1651 702 1679
rect 732 1651 766 1679
tri 780 1676 787 1683 ne
rect 787 1651 795 1683
rect 825 1651 873 1693
rect 903 1683 928 1693
rect 903 1651 911 1683
rect 1027 1679 1052 1693
rect 932 1651 966 1679
rect 996 1651 1052 1679
rect 1082 1651 1110 1693
rect 1168 1651 1196 1693
rect 1226 1679 1251 1693
rect 1350 1683 1375 1693
rect 1226 1651 1282 1679
rect 1312 1651 1346 1679
tri 1360 1676 1367 1683 ne
rect 1367 1651 1375 1683
rect 1405 1651 1453 1693
rect 1483 1683 1508 1693
rect 1483 1651 1491 1683
rect 1607 1679 1632 1693
rect 1512 1651 1546 1679
rect 1576 1651 1632 1679
rect 1662 1651 1690 1693
rect 1748 1651 1776 1693
rect 1806 1679 1831 1693
rect 1930 1683 1955 1693
rect 1806 1651 1862 1679
rect 1892 1651 1926 1679
tri 1940 1676 1947 1683 ne
rect 1947 1651 1955 1683
rect 1985 1651 2033 1693
rect 2063 1683 2088 1693
rect 2063 1651 2071 1683
rect 2187 1679 2212 1693
rect 2092 1651 2126 1679
rect 2156 1651 2212 1679
rect 2242 1651 2270 1693
rect 2328 1651 2356 1693
rect 2386 1679 2411 1693
rect 2510 1683 2535 1693
rect 2386 1651 2442 1679
rect 2472 1651 2506 1679
tri 2520 1676 2527 1683 ne
rect 2527 1651 2535 1683
rect 2565 1651 2613 1693
rect 2643 1683 2668 1693
rect 2643 1651 2651 1683
rect 2767 1679 2792 1693
rect 2672 1651 2706 1679
rect 2736 1651 2792 1679
rect 2822 1651 2850 1693
rect 2908 1651 2936 1693
rect 2966 1679 2991 1693
rect 3090 1683 3115 1693
rect 2966 1651 3022 1679
rect 3052 1651 3086 1679
tri 3100 1676 3107 1683 ne
rect 3107 1651 3115 1683
rect 3145 1651 3193 1693
rect 3223 1683 3248 1693
rect 3223 1651 3231 1683
rect 3347 1679 3372 1693
rect 3252 1651 3286 1679
rect 3316 1651 3372 1679
rect 3402 1651 3430 1693
rect 3488 1651 3516 1693
rect 3546 1679 3571 1693
rect 3670 1683 3695 1693
rect 3546 1651 3602 1679
rect 3632 1651 3666 1679
tri 3680 1676 3687 1683 ne
rect 3687 1651 3695 1683
rect 3725 1651 3773 1693
rect 3803 1683 3828 1693
rect 3803 1651 3811 1683
rect 3927 1679 3952 1693
rect 3832 1651 3866 1679
rect 3896 1651 3952 1679
rect 3982 1651 4010 1693
rect 4068 1651 4096 1693
rect 4126 1679 4151 1693
rect 4250 1683 4275 1693
rect 4126 1651 4182 1679
rect 4212 1651 4246 1679
tri 4260 1676 4267 1683 ne
rect 4267 1651 4275 1683
rect 4305 1651 4353 1693
rect 4383 1683 4408 1693
rect 4383 1651 4391 1683
rect 4507 1679 4532 1693
rect 4412 1651 4446 1679
rect 4476 1651 4532 1679
rect 4562 1651 4590 1693
rect 4648 1651 4676 1693
rect 4706 1679 4731 1693
rect 4830 1683 4855 1693
rect 4706 1651 4762 1679
rect 4792 1651 4826 1679
tri 4840 1676 4847 1683 ne
rect 4847 1651 4855 1683
rect 4885 1651 4933 1693
rect 4963 1683 4988 1693
rect 4963 1651 4971 1683
rect 5087 1679 5112 1693
rect 4992 1651 5026 1679
rect 5056 1651 5112 1679
rect 5142 1651 5170 1693
rect 5228 1651 5256 1693
rect 5286 1679 5311 1693
rect 5410 1683 5435 1693
rect 5286 1651 5342 1679
rect 5372 1651 5406 1679
tri 5420 1676 5427 1683 ne
rect 5427 1651 5435 1683
rect 5465 1651 5513 1693
rect 5543 1683 5568 1693
rect 5543 1651 5551 1683
rect 5667 1679 5692 1693
rect 5572 1651 5606 1679
rect 5636 1651 5692 1679
rect 5722 1651 5750 1693
rect 5808 1651 5836 1693
rect 5866 1679 5891 1693
rect 5990 1683 6015 1693
rect 5866 1651 5922 1679
rect 5952 1651 5986 1679
tri 6000 1676 6007 1683 ne
rect 6007 1651 6015 1683
rect 6045 1651 6093 1693
rect 6123 1683 6148 1693
rect 6123 1651 6131 1683
rect 6247 1679 6272 1693
rect 6152 1651 6186 1679
rect 6216 1651 6272 1679
rect 6302 1651 6330 1693
rect 6388 1651 6416 1693
rect 6446 1679 6471 1693
rect 6570 1683 6595 1693
rect 6446 1651 6502 1679
rect 6532 1651 6566 1679
tri 6580 1676 6587 1683 ne
rect 6587 1651 6595 1683
rect 6625 1651 6673 1693
rect 6703 1683 6728 1693
rect 6703 1651 6711 1683
rect 6827 1679 6852 1693
rect 6732 1651 6766 1679
rect 6796 1651 6852 1679
rect 6882 1651 6910 1693
rect 159 1627 186 1651
rect 253 1629 285 1651
rect 253 1627 255 1629
rect 283 1627 285 1629
rect 352 1627 379 1651
rect 159 1613 253 1627
rect 285 1613 379 1627
rect 739 1627 766 1651
rect 833 1629 865 1651
rect 833 1627 835 1629
rect 863 1627 865 1629
rect 932 1627 959 1651
rect 739 1613 833 1627
rect 865 1613 959 1627
rect 1319 1627 1346 1651
rect 1413 1629 1445 1651
rect 1413 1627 1415 1629
rect 1443 1627 1445 1629
rect 1512 1627 1539 1651
rect 1319 1613 1413 1627
rect 1445 1613 1539 1627
rect 1899 1627 1926 1651
rect 1993 1629 2025 1651
rect 1993 1627 1995 1629
rect 2023 1627 2025 1629
rect 2092 1627 2119 1651
rect 1899 1613 1993 1627
rect 2025 1613 2119 1627
rect 2479 1627 2506 1651
rect 2573 1629 2605 1651
rect 2573 1627 2575 1629
rect 2603 1627 2605 1629
rect 2672 1627 2699 1651
rect 2479 1613 2573 1627
rect 2605 1613 2699 1627
rect 3059 1627 3086 1651
rect 3153 1629 3185 1651
rect 3153 1627 3155 1629
rect 3183 1627 3185 1629
rect 3252 1627 3279 1651
rect 3059 1613 3153 1627
rect 3185 1613 3279 1627
rect 3639 1627 3666 1651
rect 3733 1629 3765 1651
rect 3733 1627 3735 1629
rect 3763 1627 3765 1629
rect 3832 1627 3859 1651
rect 3639 1613 3733 1627
rect 3765 1613 3859 1627
rect 4219 1627 4246 1651
rect 4313 1629 4345 1651
rect 4313 1627 4315 1629
rect 4343 1627 4345 1629
rect 4412 1627 4439 1651
rect 4219 1613 4313 1627
rect 4345 1613 4439 1627
rect 4799 1627 4826 1651
rect 4893 1629 4925 1651
rect 4893 1627 4895 1629
rect 4923 1627 4925 1629
rect 4992 1627 5019 1651
rect 4799 1613 4893 1627
rect 4925 1613 5019 1627
rect 5379 1627 5406 1651
rect 5473 1629 5505 1651
rect 5473 1627 5475 1629
rect 5503 1627 5505 1629
rect 5572 1627 5599 1651
rect 5379 1613 5473 1627
rect 5505 1613 5599 1627
rect 5959 1627 5986 1651
rect 6053 1629 6085 1651
rect 6053 1627 6055 1629
rect 6083 1627 6085 1629
rect 6152 1627 6179 1651
rect 5959 1613 6053 1627
rect 6085 1613 6179 1627
rect 6539 1627 6566 1651
rect 6633 1629 6665 1651
rect 6633 1627 6635 1629
rect 6663 1627 6665 1629
rect 6732 1627 6759 1651
rect 6539 1613 6633 1627
rect 6665 1613 6759 1627
rect 82 1527 100 1555
rect 130 1527 148 1555
rect 390 1527 408 1555
rect 438 1527 457 1555
rect 662 1527 680 1555
rect 710 1527 728 1555
rect 970 1527 988 1555
rect 1018 1527 1037 1555
rect 1242 1527 1260 1555
rect 1290 1527 1308 1555
rect 1550 1527 1568 1555
rect 1598 1527 1617 1555
rect 1822 1527 1840 1555
rect 1870 1527 1888 1555
rect 2130 1527 2148 1555
rect 2178 1527 2197 1555
rect 2402 1527 2420 1555
rect 2450 1527 2468 1555
rect 2710 1527 2728 1555
rect 2758 1527 2777 1555
rect 2982 1527 3000 1555
rect 3030 1527 3048 1555
rect 3290 1527 3308 1555
rect 3338 1527 3357 1555
rect 3562 1527 3580 1555
rect 3610 1527 3628 1555
rect 3870 1527 3888 1555
rect 3918 1527 3937 1555
rect 4142 1527 4160 1555
rect 4190 1527 4208 1555
rect 4450 1527 4468 1555
rect 4498 1527 4517 1555
rect 4722 1527 4740 1555
rect 4770 1527 4788 1555
rect 5030 1527 5048 1555
rect 5078 1527 5097 1555
rect 5302 1527 5320 1555
rect 5350 1527 5368 1555
rect 5610 1527 5628 1555
rect 5658 1527 5677 1555
rect 5882 1527 5900 1555
rect 5930 1527 5948 1555
rect 6190 1527 6208 1555
rect 6238 1527 6257 1555
rect 6462 1527 6480 1555
rect 6510 1527 6528 1555
rect 6770 1527 6788 1555
rect 6818 1527 6837 1555
rect 8 1381 36 1423
rect 66 1409 91 1423
rect 190 1413 215 1423
rect 66 1381 122 1409
rect 152 1381 186 1409
tri 200 1406 207 1413 ne
rect 207 1381 215 1413
rect 245 1381 293 1423
rect 323 1413 348 1423
rect 323 1381 331 1413
rect 447 1409 472 1423
rect 352 1381 386 1409
rect 416 1381 472 1409
rect 502 1381 530 1423
rect 588 1381 616 1423
rect 646 1409 671 1423
rect 770 1413 795 1423
rect 646 1381 702 1409
rect 732 1381 766 1409
tri 780 1406 787 1413 ne
rect 787 1381 795 1413
rect 825 1381 873 1423
rect 903 1413 928 1423
rect 903 1381 911 1413
rect 1027 1409 1052 1423
rect 932 1381 966 1409
rect 996 1381 1052 1409
rect 1082 1381 1110 1423
rect 1168 1381 1196 1423
rect 1226 1409 1251 1423
rect 1350 1413 1375 1423
rect 1226 1381 1282 1409
rect 1312 1381 1346 1409
tri 1360 1406 1367 1413 ne
rect 1367 1381 1375 1413
rect 1405 1381 1453 1423
rect 1483 1413 1508 1423
rect 1483 1381 1491 1413
rect 1607 1409 1632 1423
rect 1512 1381 1546 1409
rect 1576 1381 1632 1409
rect 1662 1381 1690 1423
rect 1748 1381 1776 1423
rect 1806 1409 1831 1423
rect 1930 1413 1955 1423
rect 1806 1381 1862 1409
rect 1892 1381 1926 1409
tri 1940 1406 1947 1413 ne
rect 1947 1381 1955 1413
rect 1985 1381 2033 1423
rect 2063 1413 2088 1423
rect 2063 1381 2071 1413
rect 2187 1409 2212 1423
rect 2092 1381 2126 1409
rect 2156 1381 2212 1409
rect 2242 1381 2270 1423
rect 2328 1381 2356 1423
rect 2386 1409 2411 1423
rect 2510 1413 2535 1423
rect 2386 1381 2442 1409
rect 2472 1381 2506 1409
tri 2520 1406 2527 1413 ne
rect 2527 1381 2535 1413
rect 2565 1381 2613 1423
rect 2643 1413 2668 1423
rect 2643 1381 2651 1413
rect 2767 1409 2792 1423
rect 2672 1381 2706 1409
rect 2736 1381 2792 1409
rect 2822 1381 2850 1423
rect 2908 1381 2936 1423
rect 2966 1409 2991 1423
rect 3090 1413 3115 1423
rect 2966 1381 3022 1409
rect 3052 1381 3086 1409
tri 3100 1406 3107 1413 ne
rect 3107 1381 3115 1413
rect 3145 1381 3193 1423
rect 3223 1413 3248 1423
rect 3223 1381 3231 1413
rect 3347 1409 3372 1423
rect 3252 1381 3286 1409
rect 3316 1381 3372 1409
rect 3402 1381 3430 1423
rect 3488 1381 3516 1423
rect 3546 1409 3571 1423
rect 3670 1413 3695 1423
rect 3546 1381 3602 1409
rect 3632 1381 3666 1409
tri 3680 1406 3687 1413 ne
rect 3687 1381 3695 1413
rect 3725 1381 3773 1423
rect 3803 1413 3828 1423
rect 3803 1381 3811 1413
rect 3927 1409 3952 1423
rect 3832 1381 3866 1409
rect 3896 1381 3952 1409
rect 3982 1381 4010 1423
rect 4068 1381 4096 1423
rect 4126 1409 4151 1423
rect 4250 1413 4275 1423
rect 4126 1381 4182 1409
rect 4212 1381 4246 1409
tri 4260 1406 4267 1413 ne
rect 4267 1381 4275 1413
rect 4305 1381 4353 1423
rect 4383 1413 4408 1423
rect 4383 1381 4391 1413
rect 4507 1409 4532 1423
rect 4412 1381 4446 1409
rect 4476 1381 4532 1409
rect 4562 1381 4590 1423
rect 4648 1381 4676 1423
rect 4706 1409 4731 1423
rect 4830 1413 4855 1423
rect 4706 1381 4762 1409
rect 4792 1381 4826 1409
tri 4840 1406 4847 1413 ne
rect 4847 1381 4855 1413
rect 4885 1381 4933 1423
rect 4963 1413 4988 1423
rect 4963 1381 4971 1413
rect 5087 1409 5112 1423
rect 4992 1381 5026 1409
rect 5056 1381 5112 1409
rect 5142 1381 5170 1423
rect 5228 1381 5256 1423
rect 5286 1409 5311 1423
rect 5410 1413 5435 1423
rect 5286 1381 5342 1409
rect 5372 1381 5406 1409
tri 5420 1406 5427 1413 ne
rect 5427 1381 5435 1413
rect 5465 1381 5513 1423
rect 5543 1413 5568 1423
rect 5543 1381 5551 1413
rect 5667 1409 5692 1423
rect 5572 1381 5606 1409
rect 5636 1381 5692 1409
rect 5722 1381 5750 1423
rect 5808 1381 5836 1423
rect 5866 1409 5891 1423
rect 5990 1413 6015 1423
rect 5866 1381 5922 1409
rect 5952 1381 5986 1409
tri 6000 1406 6007 1413 ne
rect 6007 1381 6015 1413
rect 6045 1381 6093 1423
rect 6123 1413 6148 1423
rect 6123 1381 6131 1413
rect 6247 1409 6272 1423
rect 6152 1381 6186 1409
rect 6216 1381 6272 1409
rect 6302 1381 6330 1423
rect 6388 1381 6416 1423
rect 6446 1409 6471 1423
rect 6570 1413 6595 1423
rect 6446 1381 6502 1409
rect 6532 1381 6566 1409
tri 6580 1406 6587 1413 ne
rect 6587 1381 6595 1413
rect 6625 1381 6673 1423
rect 6703 1413 6728 1423
rect 6703 1381 6711 1413
rect 6827 1409 6852 1423
rect 6732 1381 6766 1409
rect 6796 1381 6852 1409
rect 6882 1381 6910 1423
rect 159 1357 186 1381
rect 253 1359 285 1381
rect 253 1357 255 1359
rect 283 1357 285 1359
rect 352 1357 379 1381
rect 159 1343 253 1357
rect 285 1343 379 1357
rect 739 1357 766 1381
rect 833 1359 865 1381
rect 833 1357 835 1359
rect 863 1357 865 1359
rect 932 1357 959 1381
rect 739 1343 833 1357
rect 865 1343 959 1357
rect 1319 1357 1346 1381
rect 1413 1359 1445 1381
rect 1413 1357 1415 1359
rect 1443 1357 1445 1359
rect 1512 1357 1539 1381
rect 1319 1343 1413 1357
rect 1445 1343 1539 1357
rect 1899 1357 1926 1381
rect 1993 1359 2025 1381
rect 1993 1357 1995 1359
rect 2023 1357 2025 1359
rect 2092 1357 2119 1381
rect 1899 1343 1993 1357
rect 2025 1343 2119 1357
rect 2479 1357 2506 1381
rect 2573 1359 2605 1381
rect 2573 1357 2575 1359
rect 2603 1357 2605 1359
rect 2672 1357 2699 1381
rect 2479 1343 2573 1357
rect 2605 1343 2699 1357
rect 3059 1357 3086 1381
rect 3153 1359 3185 1381
rect 3153 1357 3155 1359
rect 3183 1357 3185 1359
rect 3252 1357 3279 1381
rect 3059 1343 3153 1357
rect 3185 1343 3279 1357
rect 3639 1357 3666 1381
rect 3733 1359 3765 1381
rect 3733 1357 3735 1359
rect 3763 1357 3765 1359
rect 3832 1357 3859 1381
rect 3639 1343 3733 1357
rect 3765 1343 3859 1357
rect 4219 1357 4246 1381
rect 4313 1359 4345 1381
rect 4313 1357 4315 1359
rect 4343 1357 4345 1359
rect 4412 1357 4439 1381
rect 4219 1343 4313 1357
rect 4345 1343 4439 1357
rect 4799 1357 4826 1381
rect 4893 1359 4925 1381
rect 4893 1357 4895 1359
rect 4923 1357 4925 1359
rect 4992 1357 5019 1381
rect 4799 1343 4893 1357
rect 4925 1343 5019 1357
rect 5379 1357 5406 1381
rect 5473 1359 5505 1381
rect 5473 1357 5475 1359
rect 5503 1357 5505 1359
rect 5572 1357 5599 1381
rect 5379 1343 5473 1357
rect 5505 1343 5599 1357
rect 5959 1357 5986 1381
rect 6053 1359 6085 1381
rect 6053 1357 6055 1359
rect 6083 1357 6085 1359
rect 6152 1357 6179 1381
rect 5959 1343 6053 1357
rect 6085 1343 6179 1357
rect 6539 1357 6566 1381
rect 6633 1359 6665 1381
rect 6633 1357 6635 1359
rect 6663 1357 6665 1359
rect 6732 1357 6759 1381
rect 6539 1343 6633 1357
rect 6665 1343 6759 1357
rect 82 1257 100 1285
rect 130 1257 148 1285
rect 390 1257 408 1285
rect 438 1257 457 1285
rect 662 1257 680 1285
rect 710 1257 728 1285
rect 970 1257 988 1285
rect 1018 1257 1037 1285
rect 1242 1257 1260 1285
rect 1290 1257 1308 1285
rect 1550 1257 1568 1285
rect 1598 1257 1617 1285
rect 1822 1257 1840 1285
rect 1870 1257 1888 1285
rect 2130 1257 2148 1285
rect 2178 1257 2197 1285
rect 2402 1257 2420 1285
rect 2450 1257 2468 1285
rect 2710 1257 2728 1285
rect 2758 1257 2777 1285
rect 2982 1257 3000 1285
rect 3030 1257 3048 1285
rect 3290 1257 3308 1285
rect 3338 1257 3357 1285
rect 3562 1257 3580 1285
rect 3610 1257 3628 1285
rect 3870 1257 3888 1285
rect 3918 1257 3937 1285
rect 4142 1257 4160 1285
rect 4190 1257 4208 1285
rect 4450 1257 4468 1285
rect 4498 1257 4517 1285
rect 4722 1257 4740 1285
rect 4770 1257 4788 1285
rect 5030 1257 5048 1285
rect 5078 1257 5097 1285
rect 5302 1257 5320 1285
rect 5350 1257 5368 1285
rect 5610 1257 5628 1285
rect 5658 1257 5677 1285
rect 5882 1257 5900 1285
rect 5930 1257 5948 1285
rect 6190 1257 6208 1285
rect 6238 1257 6257 1285
rect 6462 1257 6480 1285
rect 6510 1257 6528 1285
rect 6770 1257 6788 1285
rect 6818 1257 6837 1285
rect 8 1111 36 1153
rect 66 1139 91 1153
rect 190 1143 215 1153
rect 66 1111 122 1139
rect 152 1111 186 1139
tri 200 1136 207 1143 ne
rect 207 1111 215 1143
rect 245 1111 293 1153
rect 323 1143 348 1153
rect 323 1111 331 1143
rect 447 1139 472 1153
rect 352 1111 386 1139
rect 416 1111 472 1139
rect 502 1111 530 1153
rect 588 1111 616 1153
rect 646 1139 671 1153
rect 770 1143 795 1153
rect 646 1111 702 1139
rect 732 1111 766 1139
tri 780 1136 787 1143 ne
rect 787 1111 795 1143
rect 825 1111 873 1153
rect 903 1143 928 1153
rect 903 1111 911 1143
rect 1027 1139 1052 1153
rect 932 1111 966 1139
rect 996 1111 1052 1139
rect 1082 1111 1110 1153
rect 1168 1111 1196 1153
rect 1226 1139 1251 1153
rect 1350 1143 1375 1153
rect 1226 1111 1282 1139
rect 1312 1111 1346 1139
tri 1360 1136 1367 1143 ne
rect 1367 1111 1375 1143
rect 1405 1111 1453 1153
rect 1483 1143 1508 1153
rect 1483 1111 1491 1143
rect 1607 1139 1632 1153
rect 1512 1111 1546 1139
rect 1576 1111 1632 1139
rect 1662 1111 1690 1153
rect 1748 1111 1776 1153
rect 1806 1139 1831 1153
rect 1930 1143 1955 1153
rect 1806 1111 1862 1139
rect 1892 1111 1926 1139
tri 1940 1136 1947 1143 ne
rect 1947 1111 1955 1143
rect 1985 1111 2033 1153
rect 2063 1143 2088 1153
rect 2063 1111 2071 1143
rect 2187 1139 2212 1153
rect 2092 1111 2126 1139
rect 2156 1111 2212 1139
rect 2242 1111 2270 1153
rect 2328 1111 2356 1153
rect 2386 1139 2411 1153
rect 2510 1143 2535 1153
rect 2386 1111 2442 1139
rect 2472 1111 2506 1139
tri 2520 1136 2527 1143 ne
rect 2527 1111 2535 1143
rect 2565 1111 2613 1153
rect 2643 1143 2668 1153
rect 2643 1111 2651 1143
rect 2767 1139 2792 1153
rect 2672 1111 2706 1139
rect 2736 1111 2792 1139
rect 2822 1111 2850 1153
rect 2908 1111 2936 1153
rect 2966 1139 2991 1153
rect 3090 1143 3115 1153
rect 2966 1111 3022 1139
rect 3052 1111 3086 1139
tri 3100 1136 3107 1143 ne
rect 3107 1111 3115 1143
rect 3145 1111 3193 1153
rect 3223 1143 3248 1153
rect 3223 1111 3231 1143
rect 3347 1139 3372 1153
rect 3252 1111 3286 1139
rect 3316 1111 3372 1139
rect 3402 1111 3430 1153
rect 3488 1111 3516 1153
rect 3546 1139 3571 1153
rect 3670 1143 3695 1153
rect 3546 1111 3602 1139
rect 3632 1111 3666 1139
tri 3680 1136 3687 1143 ne
rect 3687 1111 3695 1143
rect 3725 1111 3773 1153
rect 3803 1143 3828 1153
rect 3803 1111 3811 1143
rect 3927 1139 3952 1153
rect 3832 1111 3866 1139
rect 3896 1111 3952 1139
rect 3982 1111 4010 1153
rect 4068 1111 4096 1153
rect 4126 1139 4151 1153
rect 4250 1143 4275 1153
rect 4126 1111 4182 1139
rect 4212 1111 4246 1139
tri 4260 1136 4267 1143 ne
rect 4267 1111 4275 1143
rect 4305 1111 4353 1153
rect 4383 1143 4408 1153
rect 4383 1111 4391 1143
rect 4507 1139 4532 1153
rect 4412 1111 4446 1139
rect 4476 1111 4532 1139
rect 4562 1111 4590 1153
rect 4648 1111 4676 1153
rect 4706 1139 4731 1153
rect 4830 1143 4855 1153
rect 4706 1111 4762 1139
rect 4792 1111 4826 1139
tri 4840 1136 4847 1143 ne
rect 4847 1111 4855 1143
rect 4885 1111 4933 1153
rect 4963 1143 4988 1153
rect 4963 1111 4971 1143
rect 5087 1139 5112 1153
rect 4992 1111 5026 1139
rect 5056 1111 5112 1139
rect 5142 1111 5170 1153
rect 5228 1111 5256 1153
rect 5286 1139 5311 1153
rect 5410 1143 5435 1153
rect 5286 1111 5342 1139
rect 5372 1111 5406 1139
tri 5420 1136 5427 1143 ne
rect 5427 1111 5435 1143
rect 5465 1111 5513 1153
rect 5543 1143 5568 1153
rect 5543 1111 5551 1143
rect 5667 1139 5692 1153
rect 5572 1111 5606 1139
rect 5636 1111 5692 1139
rect 5722 1111 5750 1153
rect 5808 1111 5836 1153
rect 5866 1139 5891 1153
rect 5990 1143 6015 1153
rect 5866 1111 5922 1139
rect 5952 1111 5986 1139
tri 6000 1136 6007 1143 ne
rect 6007 1111 6015 1143
rect 6045 1111 6093 1153
rect 6123 1143 6148 1153
rect 6123 1111 6131 1143
rect 6247 1139 6272 1153
rect 6152 1111 6186 1139
rect 6216 1111 6272 1139
rect 6302 1111 6330 1153
rect 6388 1111 6416 1153
rect 6446 1139 6471 1153
rect 6570 1143 6595 1153
rect 6446 1111 6502 1139
rect 6532 1111 6566 1139
tri 6580 1136 6587 1143 ne
rect 6587 1111 6595 1143
rect 6625 1111 6673 1153
rect 6703 1143 6728 1153
rect 6703 1111 6711 1143
rect 6827 1139 6852 1153
rect 6732 1111 6766 1139
rect 6796 1111 6852 1139
rect 6882 1111 6910 1153
rect 159 1087 186 1111
rect 253 1089 285 1111
rect 253 1087 255 1089
rect 283 1087 285 1089
rect 352 1087 379 1111
rect 159 1073 253 1087
rect 285 1073 379 1087
rect 739 1087 766 1111
rect 833 1089 865 1111
rect 833 1087 835 1089
rect 863 1087 865 1089
rect 932 1087 959 1111
rect 739 1073 833 1087
rect 865 1073 959 1087
rect 1319 1087 1346 1111
rect 1413 1089 1445 1111
rect 1413 1087 1415 1089
rect 1443 1087 1445 1089
rect 1512 1087 1539 1111
rect 1319 1073 1413 1087
rect 1445 1073 1539 1087
rect 1899 1087 1926 1111
rect 1993 1089 2025 1111
rect 1993 1087 1995 1089
rect 2023 1087 2025 1089
rect 2092 1087 2119 1111
rect 1899 1073 1993 1087
rect 2025 1073 2119 1087
rect 2479 1087 2506 1111
rect 2573 1089 2605 1111
rect 2573 1087 2575 1089
rect 2603 1087 2605 1089
rect 2672 1087 2699 1111
rect 2479 1073 2573 1087
rect 2605 1073 2699 1087
rect 3059 1087 3086 1111
rect 3153 1089 3185 1111
rect 3153 1087 3155 1089
rect 3183 1087 3185 1089
rect 3252 1087 3279 1111
rect 3059 1073 3153 1087
rect 3185 1073 3279 1087
rect 3639 1087 3666 1111
rect 3733 1089 3765 1111
rect 3733 1087 3735 1089
rect 3763 1087 3765 1089
rect 3832 1087 3859 1111
rect 3639 1073 3733 1087
rect 3765 1073 3859 1087
rect 4219 1087 4246 1111
rect 4313 1089 4345 1111
rect 4313 1087 4315 1089
rect 4343 1087 4345 1089
rect 4412 1087 4439 1111
rect 4219 1073 4313 1087
rect 4345 1073 4439 1087
rect 4799 1087 4826 1111
rect 4893 1089 4925 1111
rect 4893 1087 4895 1089
rect 4923 1087 4925 1089
rect 4992 1087 5019 1111
rect 4799 1073 4893 1087
rect 4925 1073 5019 1087
rect 5379 1087 5406 1111
rect 5473 1089 5505 1111
rect 5473 1087 5475 1089
rect 5503 1087 5505 1089
rect 5572 1087 5599 1111
rect 5379 1073 5473 1087
rect 5505 1073 5599 1087
rect 5959 1087 5986 1111
rect 6053 1089 6085 1111
rect 6053 1087 6055 1089
rect 6083 1087 6085 1089
rect 6152 1087 6179 1111
rect 5959 1073 6053 1087
rect 6085 1073 6179 1087
rect 6539 1087 6566 1111
rect 6633 1089 6665 1111
rect 6633 1087 6635 1089
rect 6663 1087 6665 1089
rect 6732 1087 6759 1111
rect 6539 1073 6633 1087
rect 6665 1073 6759 1087
rect 82 987 100 1015
rect 130 987 148 1015
rect 390 987 408 1015
rect 438 987 457 1015
rect 662 987 680 1015
rect 710 987 728 1015
rect 970 987 988 1015
rect 1018 987 1037 1015
rect 1242 987 1260 1015
rect 1290 987 1308 1015
rect 1550 987 1568 1015
rect 1598 987 1617 1015
rect 1822 987 1840 1015
rect 1870 987 1888 1015
rect 2130 987 2148 1015
rect 2178 987 2197 1015
rect 2402 987 2420 1015
rect 2450 987 2468 1015
rect 2710 987 2728 1015
rect 2758 987 2777 1015
rect 2982 987 3000 1015
rect 3030 987 3048 1015
rect 3290 987 3308 1015
rect 3338 987 3357 1015
rect 3562 987 3580 1015
rect 3610 987 3628 1015
rect 3870 987 3888 1015
rect 3918 987 3937 1015
rect 4142 987 4160 1015
rect 4190 987 4208 1015
rect 4450 987 4468 1015
rect 4498 987 4517 1015
rect 4722 987 4740 1015
rect 4770 987 4788 1015
rect 5030 987 5048 1015
rect 5078 987 5097 1015
rect 5302 987 5320 1015
rect 5350 987 5368 1015
rect 5610 987 5628 1015
rect 5658 987 5677 1015
rect 5882 987 5900 1015
rect 5930 987 5948 1015
rect 6190 987 6208 1015
rect 6238 987 6257 1015
rect 6462 987 6480 1015
rect 6510 987 6528 1015
rect 6770 987 6788 1015
rect 6818 987 6837 1015
rect 8 841 36 883
rect 66 869 91 883
rect 190 873 215 883
rect 66 841 122 869
rect 152 841 186 869
tri 200 866 207 873 ne
rect 207 841 215 873
rect 245 841 293 883
rect 323 873 348 883
rect 323 841 331 873
rect 447 869 472 883
rect 352 841 386 869
rect 416 841 472 869
rect 502 841 530 883
rect 588 841 616 883
rect 646 869 671 883
rect 770 873 795 883
rect 646 841 702 869
rect 732 841 766 869
tri 780 866 787 873 ne
rect 787 841 795 873
rect 825 841 873 883
rect 903 873 928 883
rect 903 841 911 873
rect 1027 869 1052 883
rect 932 841 966 869
rect 996 841 1052 869
rect 1082 841 1110 883
rect 1168 841 1196 883
rect 1226 869 1251 883
rect 1350 873 1375 883
rect 1226 841 1282 869
rect 1312 841 1346 869
tri 1360 866 1367 873 ne
rect 1367 841 1375 873
rect 1405 841 1453 883
rect 1483 873 1508 883
rect 1483 841 1491 873
rect 1607 869 1632 883
rect 1512 841 1546 869
rect 1576 841 1632 869
rect 1662 841 1690 883
rect 1748 841 1776 883
rect 1806 869 1831 883
rect 1930 873 1955 883
rect 1806 841 1862 869
rect 1892 841 1926 869
tri 1940 866 1947 873 ne
rect 1947 841 1955 873
rect 1985 841 2033 883
rect 2063 873 2088 883
rect 2063 841 2071 873
rect 2187 869 2212 883
rect 2092 841 2126 869
rect 2156 841 2212 869
rect 2242 841 2270 883
rect 2328 841 2356 883
rect 2386 869 2411 883
rect 2510 873 2535 883
rect 2386 841 2442 869
rect 2472 841 2506 869
tri 2520 866 2527 873 ne
rect 2527 841 2535 873
rect 2565 841 2613 883
rect 2643 873 2668 883
rect 2643 841 2651 873
rect 2767 869 2792 883
rect 2672 841 2706 869
rect 2736 841 2792 869
rect 2822 841 2850 883
rect 2908 841 2936 883
rect 2966 869 2991 883
rect 3090 873 3115 883
rect 2966 841 3022 869
rect 3052 841 3086 869
tri 3100 866 3107 873 ne
rect 3107 841 3115 873
rect 3145 841 3193 883
rect 3223 873 3248 883
rect 3223 841 3231 873
rect 3347 869 3372 883
rect 3252 841 3286 869
rect 3316 841 3372 869
rect 3402 841 3430 883
rect 3488 841 3516 883
rect 3546 869 3571 883
rect 3670 873 3695 883
rect 3546 841 3602 869
rect 3632 841 3666 869
tri 3680 866 3687 873 ne
rect 3687 841 3695 873
rect 3725 841 3773 883
rect 3803 873 3828 883
rect 3803 841 3811 873
rect 3927 869 3952 883
rect 3832 841 3866 869
rect 3896 841 3952 869
rect 3982 841 4010 883
rect 4068 841 4096 883
rect 4126 869 4151 883
rect 4250 873 4275 883
rect 4126 841 4182 869
rect 4212 841 4246 869
tri 4260 866 4267 873 ne
rect 4267 841 4275 873
rect 4305 841 4353 883
rect 4383 873 4408 883
rect 4383 841 4391 873
rect 4507 869 4532 883
rect 4412 841 4446 869
rect 4476 841 4532 869
rect 4562 841 4590 883
rect 4648 841 4676 883
rect 4706 869 4731 883
rect 4830 873 4855 883
rect 4706 841 4762 869
rect 4792 841 4826 869
tri 4840 866 4847 873 ne
rect 4847 841 4855 873
rect 4885 841 4933 883
rect 4963 873 4988 883
rect 4963 841 4971 873
rect 5087 869 5112 883
rect 4992 841 5026 869
rect 5056 841 5112 869
rect 5142 841 5170 883
rect 5228 841 5256 883
rect 5286 869 5311 883
rect 5410 873 5435 883
rect 5286 841 5342 869
rect 5372 841 5406 869
tri 5420 866 5427 873 ne
rect 5427 841 5435 873
rect 5465 841 5513 883
rect 5543 873 5568 883
rect 5543 841 5551 873
rect 5667 869 5692 883
rect 5572 841 5606 869
rect 5636 841 5692 869
rect 5722 841 5750 883
rect 5808 841 5836 883
rect 5866 869 5891 883
rect 5990 873 6015 883
rect 5866 841 5922 869
rect 5952 841 5986 869
tri 6000 866 6007 873 ne
rect 6007 841 6015 873
rect 6045 841 6093 883
rect 6123 873 6148 883
rect 6123 841 6131 873
rect 6247 869 6272 883
rect 6152 841 6186 869
rect 6216 841 6272 869
rect 6302 841 6330 883
rect 6388 841 6416 883
rect 6446 869 6471 883
rect 6570 873 6595 883
rect 6446 841 6502 869
rect 6532 841 6566 869
tri 6580 866 6587 873 ne
rect 6587 841 6595 873
rect 6625 841 6673 883
rect 6703 873 6728 883
rect 6703 841 6711 873
rect 6827 869 6852 883
rect 6732 841 6766 869
rect 6796 841 6852 869
rect 6882 841 6910 883
rect 159 817 186 841
rect 253 819 285 841
rect 253 817 255 819
rect 283 817 285 819
rect 352 817 379 841
rect 159 803 253 817
rect 285 803 379 817
rect 739 817 766 841
rect 833 819 865 841
rect 833 817 835 819
rect 863 817 865 819
rect 932 817 959 841
rect 739 803 833 817
rect 865 803 959 817
rect 1319 817 1346 841
rect 1413 819 1445 841
rect 1413 817 1415 819
rect 1443 817 1445 819
rect 1512 817 1539 841
rect 1319 803 1413 817
rect 1445 803 1539 817
rect 1899 817 1926 841
rect 1993 819 2025 841
rect 1993 817 1995 819
rect 2023 817 2025 819
rect 2092 817 2119 841
rect 1899 803 1993 817
rect 2025 803 2119 817
rect 2479 817 2506 841
rect 2573 819 2605 841
rect 2573 817 2575 819
rect 2603 817 2605 819
rect 2672 817 2699 841
rect 2479 803 2573 817
rect 2605 803 2699 817
rect 3059 817 3086 841
rect 3153 819 3185 841
rect 3153 817 3155 819
rect 3183 817 3185 819
rect 3252 817 3279 841
rect 3059 803 3153 817
rect 3185 803 3279 817
rect 3639 817 3666 841
rect 3733 819 3765 841
rect 3733 817 3735 819
rect 3763 817 3765 819
rect 3832 817 3859 841
rect 3639 803 3733 817
rect 3765 803 3859 817
rect 4219 817 4246 841
rect 4313 819 4345 841
rect 4313 817 4315 819
rect 4343 817 4345 819
rect 4412 817 4439 841
rect 4219 803 4313 817
rect 4345 803 4439 817
rect 4799 817 4826 841
rect 4893 819 4925 841
rect 4893 817 4895 819
rect 4923 817 4925 819
rect 4992 817 5019 841
rect 4799 803 4893 817
rect 4925 803 5019 817
rect 5379 817 5406 841
rect 5473 819 5505 841
rect 5473 817 5475 819
rect 5503 817 5505 819
rect 5572 817 5599 841
rect 5379 803 5473 817
rect 5505 803 5599 817
rect 5959 817 5986 841
rect 6053 819 6085 841
rect 6053 817 6055 819
rect 6083 817 6085 819
rect 6152 817 6179 841
rect 5959 803 6053 817
rect 6085 803 6179 817
rect 6539 817 6566 841
rect 6633 819 6665 841
rect 6633 817 6635 819
rect 6663 817 6665 819
rect 6732 817 6759 841
rect 6539 803 6633 817
rect 6665 803 6759 817
rect 82 717 100 745
rect 130 717 148 745
rect 390 717 408 745
rect 438 717 457 745
rect 662 717 680 745
rect 710 717 728 745
rect 970 717 988 745
rect 1018 717 1037 745
rect 1242 717 1260 745
rect 1290 717 1308 745
rect 1550 717 1568 745
rect 1598 717 1617 745
rect 1822 717 1840 745
rect 1870 717 1888 745
rect 2130 717 2148 745
rect 2178 717 2197 745
rect 2402 717 2420 745
rect 2450 717 2468 745
rect 2710 717 2728 745
rect 2758 717 2777 745
rect 2982 717 3000 745
rect 3030 717 3048 745
rect 3290 717 3308 745
rect 3338 717 3357 745
rect 3562 717 3580 745
rect 3610 717 3628 745
rect 3870 717 3888 745
rect 3918 717 3937 745
rect 4142 717 4160 745
rect 4190 717 4208 745
rect 4450 717 4468 745
rect 4498 717 4517 745
rect 4722 717 4740 745
rect 4770 717 4788 745
rect 5030 717 5048 745
rect 5078 717 5097 745
rect 5302 717 5320 745
rect 5350 717 5368 745
rect 5610 717 5628 745
rect 5658 717 5677 745
rect 5882 717 5900 745
rect 5930 717 5948 745
rect 6190 717 6208 745
rect 6238 717 6257 745
rect 6462 717 6480 745
rect 6510 717 6528 745
rect 6770 717 6788 745
rect 6818 717 6837 745
rect 8 571 36 613
rect 66 599 91 613
rect 190 603 215 613
rect 66 571 122 599
rect 152 571 186 599
tri 200 596 207 603 ne
rect 207 571 215 603
rect 245 571 293 613
rect 323 603 348 613
rect 323 571 331 603
rect 447 599 472 613
rect 352 571 386 599
rect 416 571 472 599
rect 502 571 530 613
rect 588 571 616 613
rect 646 599 671 613
rect 770 603 795 613
rect 646 571 702 599
rect 732 571 766 599
tri 780 596 787 603 ne
rect 787 571 795 603
rect 825 571 873 613
rect 903 603 928 613
rect 903 571 911 603
rect 1027 599 1052 613
rect 932 571 966 599
rect 996 571 1052 599
rect 1082 571 1110 613
rect 1168 571 1196 613
rect 1226 599 1251 613
rect 1350 603 1375 613
rect 1226 571 1282 599
rect 1312 571 1346 599
tri 1360 596 1367 603 ne
rect 1367 571 1375 603
rect 1405 571 1453 613
rect 1483 603 1508 613
rect 1483 571 1491 603
rect 1607 599 1632 613
rect 1512 571 1546 599
rect 1576 571 1632 599
rect 1662 571 1690 613
rect 1748 571 1776 613
rect 1806 599 1831 613
rect 1930 603 1955 613
rect 1806 571 1862 599
rect 1892 571 1926 599
tri 1940 596 1947 603 ne
rect 1947 571 1955 603
rect 1985 571 2033 613
rect 2063 603 2088 613
rect 2063 571 2071 603
rect 2187 599 2212 613
rect 2092 571 2126 599
rect 2156 571 2212 599
rect 2242 571 2270 613
rect 2328 571 2356 613
rect 2386 599 2411 613
rect 2510 603 2535 613
rect 2386 571 2442 599
rect 2472 571 2506 599
tri 2520 596 2527 603 ne
rect 2527 571 2535 603
rect 2565 571 2613 613
rect 2643 603 2668 613
rect 2643 571 2651 603
rect 2767 599 2792 613
rect 2672 571 2706 599
rect 2736 571 2792 599
rect 2822 571 2850 613
rect 2908 571 2936 613
rect 2966 599 2991 613
rect 3090 603 3115 613
rect 2966 571 3022 599
rect 3052 571 3086 599
tri 3100 596 3107 603 ne
rect 3107 571 3115 603
rect 3145 571 3193 613
rect 3223 603 3248 613
rect 3223 571 3231 603
rect 3347 599 3372 613
rect 3252 571 3286 599
rect 3316 571 3372 599
rect 3402 571 3430 613
rect 3488 571 3516 613
rect 3546 599 3571 613
rect 3670 603 3695 613
rect 3546 571 3602 599
rect 3632 571 3666 599
tri 3680 596 3687 603 ne
rect 3687 571 3695 603
rect 3725 571 3773 613
rect 3803 603 3828 613
rect 3803 571 3811 603
rect 3927 599 3952 613
rect 3832 571 3866 599
rect 3896 571 3952 599
rect 3982 571 4010 613
rect 4068 571 4096 613
rect 4126 599 4151 613
rect 4250 603 4275 613
rect 4126 571 4182 599
rect 4212 571 4246 599
tri 4260 596 4267 603 ne
rect 4267 571 4275 603
rect 4305 571 4353 613
rect 4383 603 4408 613
rect 4383 571 4391 603
rect 4507 599 4532 613
rect 4412 571 4446 599
rect 4476 571 4532 599
rect 4562 571 4590 613
rect 4648 571 4676 613
rect 4706 599 4731 613
rect 4830 603 4855 613
rect 4706 571 4762 599
rect 4792 571 4826 599
tri 4840 596 4847 603 ne
rect 4847 571 4855 603
rect 4885 571 4933 613
rect 4963 603 4988 613
rect 4963 571 4971 603
rect 5087 599 5112 613
rect 4992 571 5026 599
rect 5056 571 5112 599
rect 5142 571 5170 613
rect 5228 571 5256 613
rect 5286 599 5311 613
rect 5410 603 5435 613
rect 5286 571 5342 599
rect 5372 571 5406 599
tri 5420 596 5427 603 ne
rect 5427 571 5435 603
rect 5465 571 5513 613
rect 5543 603 5568 613
rect 5543 571 5551 603
rect 5667 599 5692 613
rect 5572 571 5606 599
rect 5636 571 5692 599
rect 5722 571 5750 613
rect 5808 571 5836 613
rect 5866 599 5891 613
rect 5990 603 6015 613
rect 5866 571 5922 599
rect 5952 571 5986 599
tri 6000 596 6007 603 ne
rect 6007 571 6015 603
rect 6045 571 6093 613
rect 6123 603 6148 613
rect 6123 571 6131 603
rect 6247 599 6272 613
rect 6152 571 6186 599
rect 6216 571 6272 599
rect 6302 571 6330 613
rect 6388 571 6416 613
rect 6446 599 6471 613
rect 6570 603 6595 613
rect 6446 571 6502 599
rect 6532 571 6566 599
tri 6580 596 6587 603 ne
rect 6587 571 6595 603
rect 6625 571 6673 613
rect 6703 603 6728 613
rect 6703 571 6711 603
rect 6827 599 6852 613
rect 6732 571 6766 599
rect 6796 571 6852 599
rect 6882 571 6910 613
rect 159 547 186 571
rect 253 549 285 571
rect 253 547 255 549
rect 283 547 285 549
rect 352 547 379 571
rect 159 533 253 547
rect 285 533 379 547
rect 739 547 766 571
rect 833 549 865 571
rect 833 547 835 549
rect 863 547 865 549
rect 932 547 959 571
rect 739 533 833 547
rect 865 533 959 547
rect 1319 547 1346 571
rect 1413 549 1445 571
rect 1413 547 1415 549
rect 1443 547 1445 549
rect 1512 547 1539 571
rect 1319 533 1413 547
rect 1445 533 1539 547
rect 1899 547 1926 571
rect 1993 549 2025 571
rect 1993 547 1995 549
rect 2023 547 2025 549
rect 2092 547 2119 571
rect 1899 533 1993 547
rect 2025 533 2119 547
rect 2479 547 2506 571
rect 2573 549 2605 571
rect 2573 547 2575 549
rect 2603 547 2605 549
rect 2672 547 2699 571
rect 2479 533 2573 547
rect 2605 533 2699 547
rect 3059 547 3086 571
rect 3153 549 3185 571
rect 3153 547 3155 549
rect 3183 547 3185 549
rect 3252 547 3279 571
rect 3059 533 3153 547
rect 3185 533 3279 547
rect 3639 547 3666 571
rect 3733 549 3765 571
rect 3733 547 3735 549
rect 3763 547 3765 549
rect 3832 547 3859 571
rect 3639 533 3733 547
rect 3765 533 3859 547
rect 4219 547 4246 571
rect 4313 549 4345 571
rect 4313 547 4315 549
rect 4343 547 4345 549
rect 4412 547 4439 571
rect 4219 533 4313 547
rect 4345 533 4439 547
rect 4799 547 4826 571
rect 4893 549 4925 571
rect 4893 547 4895 549
rect 4923 547 4925 549
rect 4992 547 5019 571
rect 4799 533 4893 547
rect 4925 533 5019 547
rect 5379 547 5406 571
rect 5473 549 5505 571
rect 5473 547 5475 549
rect 5503 547 5505 549
rect 5572 547 5599 571
rect 5379 533 5473 547
rect 5505 533 5599 547
rect 5959 547 5986 571
rect 6053 549 6085 571
rect 6053 547 6055 549
rect 6083 547 6085 549
rect 6152 547 6179 571
rect 5959 533 6053 547
rect 6085 533 6179 547
rect 6539 547 6566 571
rect 6633 549 6665 571
rect 6633 547 6635 549
rect 6663 547 6665 549
rect 6732 547 6759 571
rect 6539 533 6633 547
rect 6665 533 6759 547
rect 82 447 100 475
rect 130 447 148 475
rect 390 447 408 475
rect 438 447 457 475
rect 662 447 680 475
rect 710 447 728 475
rect 970 447 988 475
rect 1018 447 1037 475
rect 1242 447 1260 475
rect 1290 447 1308 475
rect 1550 447 1568 475
rect 1598 447 1617 475
rect 1822 447 1840 475
rect 1870 447 1888 475
rect 2130 447 2148 475
rect 2178 447 2197 475
rect 2402 447 2420 475
rect 2450 447 2468 475
rect 2710 447 2728 475
rect 2758 447 2777 475
rect 2982 447 3000 475
rect 3030 447 3048 475
rect 3290 447 3308 475
rect 3338 447 3357 475
rect 3562 447 3580 475
rect 3610 447 3628 475
rect 3870 447 3888 475
rect 3918 447 3937 475
rect 4142 447 4160 475
rect 4190 447 4208 475
rect 4450 447 4468 475
rect 4498 447 4517 475
rect 4722 447 4740 475
rect 4770 447 4788 475
rect 5030 447 5048 475
rect 5078 447 5097 475
rect 5302 447 5320 475
rect 5350 447 5368 475
rect 5610 447 5628 475
rect 5658 447 5677 475
rect 5882 447 5900 475
rect 5930 447 5948 475
rect 6190 447 6208 475
rect 6238 447 6257 475
rect 6462 447 6480 475
rect 6510 447 6528 475
rect 6770 447 6788 475
rect 6818 447 6837 475
rect 8 301 36 343
rect 66 329 91 343
rect 190 333 215 343
rect 66 301 122 329
rect 152 301 186 329
tri 200 326 207 333 ne
rect 207 301 215 333
rect 245 301 293 343
rect 323 333 348 343
rect 323 301 331 333
rect 447 329 472 343
rect 352 301 386 329
rect 416 301 472 329
rect 502 301 530 343
rect 588 301 616 343
rect 646 329 671 343
rect 770 333 795 343
rect 646 301 702 329
rect 732 301 766 329
tri 780 326 787 333 ne
rect 787 301 795 333
rect 825 301 873 343
rect 903 333 928 343
rect 903 301 911 333
rect 1027 329 1052 343
rect 932 301 966 329
rect 996 301 1052 329
rect 1082 301 1110 343
rect 1168 301 1196 343
rect 1226 329 1251 343
rect 1350 333 1375 343
rect 1226 301 1282 329
rect 1312 301 1346 329
tri 1360 326 1367 333 ne
rect 1367 301 1375 333
rect 1405 301 1453 343
rect 1483 333 1508 343
rect 1483 301 1491 333
rect 1607 329 1632 343
rect 1512 301 1546 329
rect 1576 301 1632 329
rect 1662 301 1690 343
rect 1748 301 1776 343
rect 1806 329 1831 343
rect 1930 333 1955 343
rect 1806 301 1862 329
rect 1892 301 1926 329
tri 1940 326 1947 333 ne
rect 1947 301 1955 333
rect 1985 301 2033 343
rect 2063 333 2088 343
rect 2063 301 2071 333
rect 2187 329 2212 343
rect 2092 301 2126 329
rect 2156 301 2212 329
rect 2242 301 2270 343
rect 2328 301 2356 343
rect 2386 329 2411 343
rect 2510 333 2535 343
rect 2386 301 2442 329
rect 2472 301 2506 329
tri 2520 326 2527 333 ne
rect 2527 301 2535 333
rect 2565 301 2613 343
rect 2643 333 2668 343
rect 2643 301 2651 333
rect 2767 329 2792 343
rect 2672 301 2706 329
rect 2736 301 2792 329
rect 2822 301 2850 343
rect 2908 301 2936 343
rect 2966 329 2991 343
rect 3090 333 3115 343
rect 2966 301 3022 329
rect 3052 301 3086 329
tri 3100 326 3107 333 ne
rect 3107 301 3115 333
rect 3145 301 3193 343
rect 3223 333 3248 343
rect 3223 301 3231 333
rect 3347 329 3372 343
rect 3252 301 3286 329
rect 3316 301 3372 329
rect 3402 301 3430 343
rect 3488 301 3516 343
rect 3546 329 3571 343
rect 3670 333 3695 343
rect 3546 301 3602 329
rect 3632 301 3666 329
tri 3680 326 3687 333 ne
rect 3687 301 3695 333
rect 3725 301 3773 343
rect 3803 333 3828 343
rect 3803 301 3811 333
rect 3927 329 3952 343
rect 3832 301 3866 329
rect 3896 301 3952 329
rect 3982 301 4010 343
rect 4068 301 4096 343
rect 4126 329 4151 343
rect 4250 333 4275 343
rect 4126 301 4182 329
rect 4212 301 4246 329
tri 4260 326 4267 333 ne
rect 4267 301 4275 333
rect 4305 301 4353 343
rect 4383 333 4408 343
rect 4383 301 4391 333
rect 4507 329 4532 343
rect 4412 301 4446 329
rect 4476 301 4532 329
rect 4562 301 4590 343
rect 4648 301 4676 343
rect 4706 329 4731 343
rect 4830 333 4855 343
rect 4706 301 4762 329
rect 4792 301 4826 329
tri 4840 326 4847 333 ne
rect 4847 301 4855 333
rect 4885 301 4933 343
rect 4963 333 4988 343
rect 4963 301 4971 333
rect 5087 329 5112 343
rect 4992 301 5026 329
rect 5056 301 5112 329
rect 5142 301 5170 343
rect 5228 301 5256 343
rect 5286 329 5311 343
rect 5410 333 5435 343
rect 5286 301 5342 329
rect 5372 301 5406 329
tri 5420 326 5427 333 ne
rect 5427 301 5435 333
rect 5465 301 5513 343
rect 5543 333 5568 343
rect 5543 301 5551 333
rect 5667 329 5692 343
rect 5572 301 5606 329
rect 5636 301 5692 329
rect 5722 301 5750 343
rect 5808 301 5836 343
rect 5866 329 5891 343
rect 5990 333 6015 343
rect 5866 301 5922 329
rect 5952 301 5986 329
tri 6000 326 6007 333 ne
rect 6007 301 6015 333
rect 6045 301 6093 343
rect 6123 333 6148 343
rect 6123 301 6131 333
rect 6247 329 6272 343
rect 6152 301 6186 329
rect 6216 301 6272 329
rect 6302 301 6330 343
rect 6388 301 6416 343
rect 6446 329 6471 343
rect 6570 333 6595 343
rect 6446 301 6502 329
rect 6532 301 6566 329
tri 6580 326 6587 333 ne
rect 6587 301 6595 333
rect 6625 301 6673 343
rect 6703 333 6728 343
rect 6703 301 6711 333
rect 6827 329 6852 343
rect 6732 301 6766 329
rect 6796 301 6852 329
rect 6882 301 6910 343
rect 159 277 186 301
rect 253 279 285 301
rect 253 277 255 279
rect 283 277 285 279
rect 352 277 379 301
rect 159 263 253 277
rect 285 263 379 277
rect 739 277 766 301
rect 833 279 865 301
rect 833 277 835 279
rect 863 277 865 279
rect 932 277 959 301
rect 739 263 833 277
rect 865 263 959 277
rect 1319 277 1346 301
rect 1413 279 1445 301
rect 1413 277 1415 279
rect 1443 277 1445 279
rect 1512 277 1539 301
rect 1319 263 1413 277
rect 1445 263 1539 277
rect 1899 277 1926 301
rect 1993 279 2025 301
rect 1993 277 1995 279
rect 2023 277 2025 279
rect 2092 277 2119 301
rect 1899 263 1993 277
rect 2025 263 2119 277
rect 2479 277 2506 301
rect 2573 279 2605 301
rect 2573 277 2575 279
rect 2603 277 2605 279
rect 2672 277 2699 301
rect 2479 263 2573 277
rect 2605 263 2699 277
rect 3059 277 3086 301
rect 3153 279 3185 301
rect 3153 277 3155 279
rect 3183 277 3185 279
rect 3252 277 3279 301
rect 3059 263 3153 277
rect 3185 263 3279 277
rect 3639 277 3666 301
rect 3733 279 3765 301
rect 3733 277 3735 279
rect 3763 277 3765 279
rect 3832 277 3859 301
rect 3639 263 3733 277
rect 3765 263 3859 277
rect 4219 277 4246 301
rect 4313 279 4345 301
rect 4313 277 4315 279
rect 4343 277 4345 279
rect 4412 277 4439 301
rect 4219 263 4313 277
rect 4345 263 4439 277
rect 4799 277 4826 301
rect 4893 279 4925 301
rect 4893 277 4895 279
rect 4923 277 4925 279
rect 4992 277 5019 301
rect 4799 263 4893 277
rect 4925 263 5019 277
rect 5379 277 5406 301
rect 5473 279 5505 301
rect 5473 277 5475 279
rect 5503 277 5505 279
rect 5572 277 5599 301
rect 5379 263 5473 277
rect 5505 263 5599 277
rect 5959 277 5986 301
rect 6053 279 6085 301
rect 6053 277 6055 279
rect 6083 277 6085 279
rect 6152 277 6179 301
rect 5959 263 6053 277
rect 6085 263 6179 277
rect 6539 277 6566 301
rect 6633 279 6665 301
rect 6633 277 6635 279
rect 6663 277 6665 279
rect 6732 277 6759 301
rect 6539 263 6633 277
rect 6665 263 6759 277
rect 82 177 100 205
rect 130 177 148 205
rect 390 177 408 205
rect 438 177 457 205
rect 662 177 680 205
rect 710 177 728 205
rect 970 177 988 205
rect 1018 177 1037 205
rect 1242 177 1260 205
rect 1290 177 1308 205
rect 1550 177 1568 205
rect 1598 177 1617 205
rect 1822 177 1840 205
rect 1870 177 1888 205
rect 2130 177 2148 205
rect 2178 177 2197 205
rect 2402 177 2420 205
rect 2450 177 2468 205
rect 2710 177 2728 205
rect 2758 177 2777 205
rect 2982 177 3000 205
rect 3030 177 3048 205
rect 3290 177 3308 205
rect 3338 177 3357 205
rect 3562 177 3580 205
rect 3610 177 3628 205
rect 3870 177 3888 205
rect 3918 177 3937 205
rect 4142 177 4160 205
rect 4190 177 4208 205
rect 4450 177 4468 205
rect 4498 177 4517 205
rect 4722 177 4740 205
rect 4770 177 4788 205
rect 5030 177 5048 205
rect 5078 177 5097 205
rect 5302 177 5320 205
rect 5350 177 5368 205
rect 5610 177 5628 205
rect 5658 177 5677 205
rect 5882 177 5900 205
rect 5930 177 5948 205
rect 6190 177 6208 205
rect 6238 177 6257 205
rect 6462 177 6480 205
rect 6510 177 6528 205
rect 6770 177 6788 205
rect 6818 177 6837 205
rect 8 31 36 73
rect 66 59 91 73
rect 190 63 215 73
rect 66 31 122 59
rect 152 31 186 59
tri 200 56 207 63 ne
rect 207 31 215 63
rect 245 31 293 73
rect 323 63 348 73
rect 323 31 331 63
rect 447 59 472 73
rect 352 31 386 59
rect 416 31 472 59
rect 502 31 530 73
rect 588 31 616 73
rect 646 59 671 73
rect 770 63 795 73
rect 646 31 702 59
rect 732 31 766 59
tri 780 56 787 63 ne
rect 787 31 795 63
rect 825 31 873 73
rect 903 63 928 73
rect 903 31 911 63
rect 1027 59 1052 73
rect 932 31 966 59
rect 996 31 1052 59
rect 1082 31 1110 73
rect 1168 31 1196 73
rect 1226 59 1251 73
rect 1350 63 1375 73
rect 1226 31 1282 59
rect 1312 31 1346 59
tri 1360 56 1367 63 ne
rect 1367 31 1375 63
rect 1405 31 1453 73
rect 1483 63 1508 73
rect 1483 31 1491 63
rect 1607 59 1632 73
rect 1512 31 1546 59
rect 1576 31 1632 59
rect 1662 31 1690 73
rect 1748 31 1776 73
rect 1806 59 1831 73
rect 1930 63 1955 73
rect 1806 31 1862 59
rect 1892 31 1926 59
tri 1940 56 1947 63 ne
rect 1947 31 1955 63
rect 1985 31 2033 73
rect 2063 63 2088 73
rect 2063 31 2071 63
rect 2187 59 2212 73
rect 2092 31 2126 59
rect 2156 31 2212 59
rect 2242 31 2270 73
rect 2328 31 2356 73
rect 2386 59 2411 73
rect 2510 63 2535 73
rect 2386 31 2442 59
rect 2472 31 2506 59
tri 2520 56 2527 63 ne
rect 2527 31 2535 63
rect 2565 31 2613 73
rect 2643 63 2668 73
rect 2643 31 2651 63
rect 2767 59 2792 73
rect 2672 31 2706 59
rect 2736 31 2792 59
rect 2822 31 2850 73
rect 2908 31 2936 73
rect 2966 59 2991 73
rect 3090 63 3115 73
rect 2966 31 3022 59
rect 3052 31 3086 59
tri 3100 56 3107 63 ne
rect 3107 31 3115 63
rect 3145 31 3193 73
rect 3223 63 3248 73
rect 3223 31 3231 63
rect 3347 59 3372 73
rect 3252 31 3286 59
rect 3316 31 3372 59
rect 3402 31 3430 73
rect 3488 31 3516 73
rect 3546 59 3571 73
rect 3670 63 3695 73
rect 3546 31 3602 59
rect 3632 31 3666 59
tri 3680 56 3687 63 ne
rect 3687 31 3695 63
rect 3725 31 3773 73
rect 3803 63 3828 73
rect 3803 31 3811 63
rect 3927 59 3952 73
rect 3832 31 3866 59
rect 3896 31 3952 59
rect 3982 31 4010 73
rect 4068 31 4096 73
rect 4126 59 4151 73
rect 4250 63 4275 73
rect 4126 31 4182 59
rect 4212 31 4246 59
tri 4260 56 4267 63 ne
rect 4267 31 4275 63
rect 4305 31 4353 73
rect 4383 63 4408 73
rect 4383 31 4391 63
rect 4507 59 4532 73
rect 4412 31 4446 59
rect 4476 31 4532 59
rect 4562 31 4590 73
rect 4648 31 4676 73
rect 4706 59 4731 73
rect 4830 63 4855 73
rect 4706 31 4762 59
rect 4792 31 4826 59
tri 4840 56 4847 63 ne
rect 4847 31 4855 63
rect 4885 31 4933 73
rect 4963 63 4988 73
rect 4963 31 4971 63
rect 5087 59 5112 73
rect 4992 31 5026 59
rect 5056 31 5112 59
rect 5142 31 5170 73
rect 5228 31 5256 73
rect 5286 59 5311 73
rect 5410 63 5435 73
rect 5286 31 5342 59
rect 5372 31 5406 59
tri 5420 56 5427 63 ne
rect 5427 31 5435 63
rect 5465 31 5513 73
rect 5543 63 5568 73
rect 5543 31 5551 63
rect 5667 59 5692 73
rect 5572 31 5606 59
rect 5636 31 5692 59
rect 5722 31 5750 73
rect 5808 31 5836 73
rect 5866 59 5891 73
rect 5990 63 6015 73
rect 5866 31 5922 59
rect 5952 31 5986 59
tri 6000 56 6007 63 ne
rect 6007 31 6015 63
rect 6045 31 6093 73
rect 6123 63 6148 73
rect 6123 31 6131 63
rect 6247 59 6272 73
rect 6152 31 6186 59
rect 6216 31 6272 59
rect 6302 31 6330 73
rect 6388 31 6416 73
rect 6446 59 6471 73
rect 6570 63 6595 73
rect 6446 31 6502 59
rect 6532 31 6566 59
tri 6580 56 6587 63 ne
rect 6587 31 6595 63
rect 6625 31 6673 73
rect 6703 63 6728 73
rect 6703 31 6711 63
rect 6827 59 6852 73
rect 6732 31 6766 59
rect 6796 31 6852 59
rect 6882 31 6910 73
rect 159 7 186 31
rect 253 9 285 31
rect 253 7 255 9
rect 283 7 285 9
rect 352 7 379 31
rect 159 -7 253 7
rect 285 -7 379 7
rect 739 7 766 31
rect 833 9 865 31
rect 833 7 835 9
rect 863 7 865 9
rect 932 7 959 31
rect 739 -7 833 7
rect 865 -7 959 7
rect 1319 7 1346 31
rect 1413 9 1445 31
rect 1413 7 1415 9
rect 1443 7 1445 9
rect 1512 7 1539 31
rect 1319 -7 1413 7
rect 1445 -7 1539 7
rect 1899 7 1926 31
rect 1993 9 2025 31
rect 1993 7 1995 9
rect 2023 7 2025 9
rect 2092 7 2119 31
rect 1899 -7 1993 7
rect 2025 -7 2119 7
rect 2479 7 2506 31
rect 2573 9 2605 31
rect 2573 7 2575 9
rect 2603 7 2605 9
rect 2672 7 2699 31
rect 2479 -7 2573 7
rect 2605 -7 2699 7
rect 3059 7 3086 31
rect 3153 9 3185 31
rect 3153 7 3155 9
rect 3183 7 3185 9
rect 3252 7 3279 31
rect 3059 -7 3153 7
rect 3185 -7 3279 7
rect 3639 7 3666 31
rect 3733 9 3765 31
rect 3733 7 3735 9
rect 3763 7 3765 9
rect 3832 7 3859 31
rect 3639 -7 3733 7
rect 3765 -7 3859 7
rect 4219 7 4246 31
rect 4313 9 4345 31
rect 4313 7 4315 9
rect 4343 7 4345 9
rect 4412 7 4439 31
rect 4219 -7 4313 7
rect 4345 -7 4439 7
rect 4799 7 4826 31
rect 4893 9 4925 31
rect 4893 7 4895 9
rect 4923 7 4925 9
rect 4992 7 5019 31
rect 4799 -7 4893 7
rect 4925 -7 5019 7
rect 5379 7 5406 31
rect 5473 9 5505 31
rect 5473 7 5475 9
rect 5503 7 5505 9
rect 5572 7 5599 31
rect 5379 -7 5473 7
rect 5505 -7 5599 7
rect 5959 7 5986 31
rect 6053 9 6085 31
rect 6053 7 6055 9
rect 6083 7 6085 9
rect 6152 7 6179 31
rect 5959 -7 6053 7
rect 6085 -7 6179 7
rect 6539 7 6566 31
rect 6633 9 6665 31
rect 6633 7 6635 9
rect 6663 7 6665 9
rect 6732 7 6759 31
rect 6539 -7 6633 7
rect 6665 -7 6759 7
<< pdiff >>
rect 253 4267 255 4269
rect 283 4267 285 4269
rect 253 4245 285 4267
rect 206 4217 215 4245
rect 245 4217 293 4245
rect 323 4217 332 4245
tri 332 4217 344 4229 sw
rect 833 4267 835 4269
rect 863 4267 865 4269
rect 833 4245 865 4267
rect 786 4217 795 4245
rect 825 4217 873 4245
rect 903 4217 912 4245
tri 912 4217 924 4229 sw
rect 1413 4267 1415 4269
rect 1443 4267 1445 4269
rect 1413 4245 1445 4267
rect 1366 4217 1375 4245
rect 1405 4217 1453 4245
rect 1483 4217 1492 4245
tri 1492 4217 1504 4229 sw
rect 1993 4267 1995 4269
rect 2023 4267 2025 4269
rect 1993 4245 2025 4267
rect 1946 4217 1955 4245
rect 1985 4217 2033 4245
rect 2063 4217 2072 4245
tri 2072 4217 2084 4229 sw
rect 2573 4267 2575 4269
rect 2603 4267 2605 4269
rect 2573 4245 2605 4267
rect 2526 4217 2535 4245
rect 2565 4217 2613 4245
rect 2643 4217 2652 4245
tri 2652 4217 2664 4229 sw
rect 3153 4267 3155 4269
rect 3183 4267 3185 4269
rect 3153 4245 3185 4267
rect 3106 4217 3115 4245
rect 3145 4217 3193 4245
rect 3223 4217 3232 4245
tri 3232 4217 3244 4229 sw
rect 3733 4267 3735 4269
rect 3763 4267 3765 4269
rect 3733 4245 3765 4267
rect 3686 4217 3695 4245
rect 3725 4217 3773 4245
rect 3803 4217 3812 4245
tri 3812 4217 3824 4229 sw
rect 4313 4267 4315 4269
rect 4343 4267 4345 4269
rect 4313 4245 4345 4267
rect 4266 4217 4275 4245
rect 4305 4217 4353 4245
rect 4383 4217 4392 4245
tri 4392 4217 4404 4229 sw
rect 4893 4267 4895 4269
rect 4923 4267 4925 4269
rect 4893 4245 4925 4267
rect 4846 4217 4855 4245
rect 4885 4217 4933 4245
rect 4963 4217 4972 4245
tri 4972 4217 4984 4229 sw
rect 5473 4267 5475 4269
rect 5503 4267 5505 4269
rect 5473 4245 5505 4267
rect 5426 4217 5435 4245
rect 5465 4217 5513 4245
rect 5543 4217 5552 4245
tri 5552 4217 5564 4229 sw
rect 6053 4267 6055 4269
rect 6083 4267 6085 4269
rect 6053 4245 6085 4267
rect 6006 4217 6015 4245
rect 6045 4217 6093 4245
rect 6123 4217 6132 4245
tri 6132 4217 6144 4229 sw
rect 6633 4267 6635 4269
rect 6663 4267 6665 4269
rect 6633 4245 6665 4267
rect 6586 4217 6595 4245
rect 6625 4217 6673 4245
rect 6703 4217 6712 4245
tri 6712 4217 6724 4229 sw
rect 253 3997 255 3999
rect 283 3997 285 3999
rect 253 3975 285 3997
rect 206 3947 215 3975
rect 245 3947 293 3975
rect 323 3947 332 3975
tri 332 3947 344 3959 sw
rect 833 3997 835 3999
rect 863 3997 865 3999
rect 833 3975 865 3997
rect 786 3947 795 3975
rect 825 3947 873 3975
rect 903 3947 912 3975
tri 912 3947 924 3959 sw
rect 1413 3997 1415 3999
rect 1443 3997 1445 3999
rect 1413 3975 1445 3997
rect 1366 3947 1375 3975
rect 1405 3947 1453 3975
rect 1483 3947 1492 3975
tri 1492 3947 1504 3959 sw
rect 1993 3997 1995 3999
rect 2023 3997 2025 3999
rect 1993 3975 2025 3997
rect 1946 3947 1955 3975
rect 1985 3947 2033 3975
rect 2063 3947 2072 3975
tri 2072 3947 2084 3959 sw
rect 2573 3997 2575 3999
rect 2603 3997 2605 3999
rect 2573 3975 2605 3997
rect 2526 3947 2535 3975
rect 2565 3947 2613 3975
rect 2643 3947 2652 3975
tri 2652 3947 2664 3959 sw
rect 3153 3997 3155 3999
rect 3183 3997 3185 3999
rect 3153 3975 3185 3997
rect 3106 3947 3115 3975
rect 3145 3947 3193 3975
rect 3223 3947 3232 3975
tri 3232 3947 3244 3959 sw
rect 3733 3997 3735 3999
rect 3763 3997 3765 3999
rect 3733 3975 3765 3997
rect 3686 3947 3695 3975
rect 3725 3947 3773 3975
rect 3803 3947 3812 3975
tri 3812 3947 3824 3959 sw
rect 4313 3997 4315 3999
rect 4343 3997 4345 3999
rect 4313 3975 4345 3997
rect 4266 3947 4275 3975
rect 4305 3947 4353 3975
rect 4383 3947 4392 3975
tri 4392 3947 4404 3959 sw
rect 4893 3997 4895 3999
rect 4923 3997 4925 3999
rect 4893 3975 4925 3997
rect 4846 3947 4855 3975
rect 4885 3947 4933 3975
rect 4963 3947 4972 3975
tri 4972 3947 4984 3959 sw
rect 5473 3997 5475 3999
rect 5503 3997 5505 3999
rect 5473 3975 5505 3997
rect 5426 3947 5435 3975
rect 5465 3947 5513 3975
rect 5543 3947 5552 3975
tri 5552 3947 5564 3959 sw
rect 6053 3997 6055 3999
rect 6083 3997 6085 3999
rect 6053 3975 6085 3997
rect 6006 3947 6015 3975
rect 6045 3947 6093 3975
rect 6123 3947 6132 3975
tri 6132 3947 6144 3959 sw
rect 6633 3997 6635 3999
rect 6663 3997 6665 3999
rect 6633 3975 6665 3997
rect 6586 3947 6595 3975
rect 6625 3947 6673 3975
rect 6703 3947 6712 3975
tri 6712 3947 6724 3959 sw
rect 253 3727 255 3729
rect 283 3727 285 3729
rect 253 3705 285 3727
rect 206 3677 215 3705
rect 245 3677 293 3705
rect 323 3677 332 3705
tri 332 3677 344 3689 sw
rect 833 3727 835 3729
rect 863 3727 865 3729
rect 833 3705 865 3727
rect 786 3677 795 3705
rect 825 3677 873 3705
rect 903 3677 912 3705
tri 912 3677 924 3689 sw
rect 1413 3727 1415 3729
rect 1443 3727 1445 3729
rect 1413 3705 1445 3727
rect 1366 3677 1375 3705
rect 1405 3677 1453 3705
rect 1483 3677 1492 3705
tri 1492 3677 1504 3689 sw
rect 1993 3727 1995 3729
rect 2023 3727 2025 3729
rect 1993 3705 2025 3727
rect 1946 3677 1955 3705
rect 1985 3677 2033 3705
rect 2063 3677 2072 3705
tri 2072 3677 2084 3689 sw
rect 2573 3727 2575 3729
rect 2603 3727 2605 3729
rect 2573 3705 2605 3727
rect 2526 3677 2535 3705
rect 2565 3677 2613 3705
rect 2643 3677 2652 3705
tri 2652 3677 2664 3689 sw
rect 3153 3727 3155 3729
rect 3183 3727 3185 3729
rect 3153 3705 3185 3727
rect 3106 3677 3115 3705
rect 3145 3677 3193 3705
rect 3223 3677 3232 3705
tri 3232 3677 3244 3689 sw
rect 3733 3727 3735 3729
rect 3763 3727 3765 3729
rect 3733 3705 3765 3727
rect 3686 3677 3695 3705
rect 3725 3677 3773 3705
rect 3803 3677 3812 3705
tri 3812 3677 3824 3689 sw
rect 4313 3727 4315 3729
rect 4343 3727 4345 3729
rect 4313 3705 4345 3727
rect 4266 3677 4275 3705
rect 4305 3677 4353 3705
rect 4383 3677 4392 3705
tri 4392 3677 4404 3689 sw
rect 4893 3727 4895 3729
rect 4923 3727 4925 3729
rect 4893 3705 4925 3727
rect 4846 3677 4855 3705
rect 4885 3677 4933 3705
rect 4963 3677 4972 3705
tri 4972 3677 4984 3689 sw
rect 5473 3727 5475 3729
rect 5503 3727 5505 3729
rect 5473 3705 5505 3727
rect 5426 3677 5435 3705
rect 5465 3677 5513 3705
rect 5543 3677 5552 3705
tri 5552 3677 5564 3689 sw
rect 6053 3727 6055 3729
rect 6083 3727 6085 3729
rect 6053 3705 6085 3727
rect 6006 3677 6015 3705
rect 6045 3677 6093 3705
rect 6123 3677 6132 3705
tri 6132 3677 6144 3689 sw
rect 6633 3727 6635 3729
rect 6663 3727 6665 3729
rect 6633 3705 6665 3727
rect 6586 3677 6595 3705
rect 6625 3677 6673 3705
rect 6703 3677 6712 3705
tri 6712 3677 6724 3689 sw
rect 253 3457 255 3459
rect 283 3457 285 3459
rect 253 3435 285 3457
rect 206 3407 215 3435
rect 245 3407 293 3435
rect 323 3407 332 3435
tri 332 3407 344 3419 sw
rect 833 3457 835 3459
rect 863 3457 865 3459
rect 833 3435 865 3457
rect 786 3407 795 3435
rect 825 3407 873 3435
rect 903 3407 912 3435
tri 912 3407 924 3419 sw
rect 1413 3457 1415 3459
rect 1443 3457 1445 3459
rect 1413 3435 1445 3457
rect 1366 3407 1375 3435
rect 1405 3407 1453 3435
rect 1483 3407 1492 3435
tri 1492 3407 1504 3419 sw
rect 1993 3457 1995 3459
rect 2023 3457 2025 3459
rect 1993 3435 2025 3457
rect 1946 3407 1955 3435
rect 1985 3407 2033 3435
rect 2063 3407 2072 3435
tri 2072 3407 2084 3419 sw
rect 2573 3457 2575 3459
rect 2603 3457 2605 3459
rect 2573 3435 2605 3457
rect 2526 3407 2535 3435
rect 2565 3407 2613 3435
rect 2643 3407 2652 3435
tri 2652 3407 2664 3419 sw
rect 3153 3457 3155 3459
rect 3183 3457 3185 3459
rect 3153 3435 3185 3457
rect 3106 3407 3115 3435
rect 3145 3407 3193 3435
rect 3223 3407 3232 3435
tri 3232 3407 3244 3419 sw
rect 3733 3457 3735 3459
rect 3763 3457 3765 3459
rect 3733 3435 3765 3457
rect 3686 3407 3695 3435
rect 3725 3407 3773 3435
rect 3803 3407 3812 3435
tri 3812 3407 3824 3419 sw
rect 4313 3457 4315 3459
rect 4343 3457 4345 3459
rect 4313 3435 4345 3457
rect 4266 3407 4275 3435
rect 4305 3407 4353 3435
rect 4383 3407 4392 3435
tri 4392 3407 4404 3419 sw
rect 4893 3457 4895 3459
rect 4923 3457 4925 3459
rect 4893 3435 4925 3457
rect 4846 3407 4855 3435
rect 4885 3407 4933 3435
rect 4963 3407 4972 3435
tri 4972 3407 4984 3419 sw
rect 5473 3457 5475 3459
rect 5503 3457 5505 3459
rect 5473 3435 5505 3457
rect 5426 3407 5435 3435
rect 5465 3407 5513 3435
rect 5543 3407 5552 3435
tri 5552 3407 5564 3419 sw
rect 6053 3457 6055 3459
rect 6083 3457 6085 3459
rect 6053 3435 6085 3457
rect 6006 3407 6015 3435
rect 6045 3407 6093 3435
rect 6123 3407 6132 3435
tri 6132 3407 6144 3419 sw
rect 6633 3457 6635 3459
rect 6663 3457 6665 3459
rect 6633 3435 6665 3457
rect 6586 3407 6595 3435
rect 6625 3407 6673 3435
rect 6703 3407 6712 3435
tri 6712 3407 6724 3419 sw
rect 253 3187 255 3189
rect 283 3187 285 3189
rect 253 3165 285 3187
rect 206 3137 215 3165
rect 245 3137 293 3165
rect 323 3137 332 3165
tri 332 3137 344 3149 sw
rect 833 3187 835 3189
rect 863 3187 865 3189
rect 833 3165 865 3187
rect 786 3137 795 3165
rect 825 3137 873 3165
rect 903 3137 912 3165
tri 912 3137 924 3149 sw
rect 1413 3187 1415 3189
rect 1443 3187 1445 3189
rect 1413 3165 1445 3187
rect 1366 3137 1375 3165
rect 1405 3137 1453 3165
rect 1483 3137 1492 3165
tri 1492 3137 1504 3149 sw
rect 1993 3187 1995 3189
rect 2023 3187 2025 3189
rect 1993 3165 2025 3187
rect 1946 3137 1955 3165
rect 1985 3137 2033 3165
rect 2063 3137 2072 3165
tri 2072 3137 2084 3149 sw
rect 2573 3187 2575 3189
rect 2603 3187 2605 3189
rect 2573 3165 2605 3187
rect 2526 3137 2535 3165
rect 2565 3137 2613 3165
rect 2643 3137 2652 3165
tri 2652 3137 2664 3149 sw
rect 3153 3187 3155 3189
rect 3183 3187 3185 3189
rect 3153 3165 3185 3187
rect 3106 3137 3115 3165
rect 3145 3137 3193 3165
rect 3223 3137 3232 3165
tri 3232 3137 3244 3149 sw
rect 3733 3187 3735 3189
rect 3763 3187 3765 3189
rect 3733 3165 3765 3187
rect 3686 3137 3695 3165
rect 3725 3137 3773 3165
rect 3803 3137 3812 3165
tri 3812 3137 3824 3149 sw
rect 4313 3187 4315 3189
rect 4343 3187 4345 3189
rect 4313 3165 4345 3187
rect 4266 3137 4275 3165
rect 4305 3137 4353 3165
rect 4383 3137 4392 3165
tri 4392 3137 4404 3149 sw
rect 4893 3187 4895 3189
rect 4923 3187 4925 3189
rect 4893 3165 4925 3187
rect 4846 3137 4855 3165
rect 4885 3137 4933 3165
rect 4963 3137 4972 3165
tri 4972 3137 4984 3149 sw
rect 5473 3187 5475 3189
rect 5503 3187 5505 3189
rect 5473 3165 5505 3187
rect 5426 3137 5435 3165
rect 5465 3137 5513 3165
rect 5543 3137 5552 3165
tri 5552 3137 5564 3149 sw
rect 6053 3187 6055 3189
rect 6083 3187 6085 3189
rect 6053 3165 6085 3187
rect 6006 3137 6015 3165
rect 6045 3137 6093 3165
rect 6123 3137 6132 3165
tri 6132 3137 6144 3149 sw
rect 6633 3187 6635 3189
rect 6663 3187 6665 3189
rect 6633 3165 6665 3187
rect 6586 3137 6595 3165
rect 6625 3137 6673 3165
rect 6703 3137 6712 3165
tri 6712 3137 6724 3149 sw
rect 253 2917 255 2919
rect 283 2917 285 2919
rect 253 2895 285 2917
rect 206 2867 215 2895
rect 245 2867 293 2895
rect 323 2867 332 2895
tri 332 2867 344 2879 sw
rect 833 2917 835 2919
rect 863 2917 865 2919
rect 833 2895 865 2917
rect 786 2867 795 2895
rect 825 2867 873 2895
rect 903 2867 912 2895
tri 912 2867 924 2879 sw
rect 1413 2917 1415 2919
rect 1443 2917 1445 2919
rect 1413 2895 1445 2917
rect 1366 2867 1375 2895
rect 1405 2867 1453 2895
rect 1483 2867 1492 2895
tri 1492 2867 1504 2879 sw
rect 1993 2917 1995 2919
rect 2023 2917 2025 2919
rect 1993 2895 2025 2917
rect 1946 2867 1955 2895
rect 1985 2867 2033 2895
rect 2063 2867 2072 2895
tri 2072 2867 2084 2879 sw
rect 2573 2917 2575 2919
rect 2603 2917 2605 2919
rect 2573 2895 2605 2917
rect 2526 2867 2535 2895
rect 2565 2867 2613 2895
rect 2643 2867 2652 2895
tri 2652 2867 2664 2879 sw
rect 3153 2917 3155 2919
rect 3183 2917 3185 2919
rect 3153 2895 3185 2917
rect 3106 2867 3115 2895
rect 3145 2867 3193 2895
rect 3223 2867 3232 2895
tri 3232 2867 3244 2879 sw
rect 3733 2917 3735 2919
rect 3763 2917 3765 2919
rect 3733 2895 3765 2917
rect 3686 2867 3695 2895
rect 3725 2867 3773 2895
rect 3803 2867 3812 2895
tri 3812 2867 3824 2879 sw
rect 4313 2917 4315 2919
rect 4343 2917 4345 2919
rect 4313 2895 4345 2917
rect 4266 2867 4275 2895
rect 4305 2867 4353 2895
rect 4383 2867 4392 2895
tri 4392 2867 4404 2879 sw
rect 4893 2917 4895 2919
rect 4923 2917 4925 2919
rect 4893 2895 4925 2917
rect 4846 2867 4855 2895
rect 4885 2867 4933 2895
rect 4963 2867 4972 2895
tri 4972 2867 4984 2879 sw
rect 5473 2917 5475 2919
rect 5503 2917 5505 2919
rect 5473 2895 5505 2917
rect 5426 2867 5435 2895
rect 5465 2867 5513 2895
rect 5543 2867 5552 2895
tri 5552 2867 5564 2879 sw
rect 6053 2917 6055 2919
rect 6083 2917 6085 2919
rect 6053 2895 6085 2917
rect 6006 2867 6015 2895
rect 6045 2867 6093 2895
rect 6123 2867 6132 2895
tri 6132 2867 6144 2879 sw
rect 6633 2917 6635 2919
rect 6663 2917 6665 2919
rect 6633 2895 6665 2917
rect 6586 2867 6595 2895
rect 6625 2867 6673 2895
rect 6703 2867 6712 2895
tri 6712 2867 6724 2879 sw
rect 253 2647 255 2649
rect 283 2647 285 2649
rect 253 2625 285 2647
rect 206 2597 215 2625
rect 245 2597 293 2625
rect 323 2597 332 2625
tri 332 2597 344 2609 sw
rect 833 2647 835 2649
rect 863 2647 865 2649
rect 833 2625 865 2647
rect 786 2597 795 2625
rect 825 2597 873 2625
rect 903 2597 912 2625
tri 912 2597 924 2609 sw
rect 1413 2647 1415 2649
rect 1443 2647 1445 2649
rect 1413 2625 1445 2647
rect 1366 2597 1375 2625
rect 1405 2597 1453 2625
rect 1483 2597 1492 2625
tri 1492 2597 1504 2609 sw
rect 1993 2647 1995 2649
rect 2023 2647 2025 2649
rect 1993 2625 2025 2647
rect 1946 2597 1955 2625
rect 1985 2597 2033 2625
rect 2063 2597 2072 2625
tri 2072 2597 2084 2609 sw
rect 2573 2647 2575 2649
rect 2603 2647 2605 2649
rect 2573 2625 2605 2647
rect 2526 2597 2535 2625
rect 2565 2597 2613 2625
rect 2643 2597 2652 2625
tri 2652 2597 2664 2609 sw
rect 3153 2647 3155 2649
rect 3183 2647 3185 2649
rect 3153 2625 3185 2647
rect 3106 2597 3115 2625
rect 3145 2597 3193 2625
rect 3223 2597 3232 2625
tri 3232 2597 3244 2609 sw
rect 3733 2647 3735 2649
rect 3763 2647 3765 2649
rect 3733 2625 3765 2647
rect 3686 2597 3695 2625
rect 3725 2597 3773 2625
rect 3803 2597 3812 2625
tri 3812 2597 3824 2609 sw
rect 4313 2647 4315 2649
rect 4343 2647 4345 2649
rect 4313 2625 4345 2647
rect 4266 2597 4275 2625
rect 4305 2597 4353 2625
rect 4383 2597 4392 2625
tri 4392 2597 4404 2609 sw
rect 4893 2647 4895 2649
rect 4923 2647 4925 2649
rect 4893 2625 4925 2647
rect 4846 2597 4855 2625
rect 4885 2597 4933 2625
rect 4963 2597 4972 2625
tri 4972 2597 4984 2609 sw
rect 5473 2647 5475 2649
rect 5503 2647 5505 2649
rect 5473 2625 5505 2647
rect 5426 2597 5435 2625
rect 5465 2597 5513 2625
rect 5543 2597 5552 2625
tri 5552 2597 5564 2609 sw
rect 6053 2647 6055 2649
rect 6083 2647 6085 2649
rect 6053 2625 6085 2647
rect 6006 2597 6015 2625
rect 6045 2597 6093 2625
rect 6123 2597 6132 2625
tri 6132 2597 6144 2609 sw
rect 6633 2647 6635 2649
rect 6663 2647 6665 2649
rect 6633 2625 6665 2647
rect 6586 2597 6595 2625
rect 6625 2597 6673 2625
rect 6703 2597 6712 2625
tri 6712 2597 6724 2609 sw
rect 253 2377 255 2379
rect 283 2377 285 2379
rect 253 2355 285 2377
rect 206 2327 215 2355
rect 245 2327 293 2355
rect 323 2327 332 2355
tri 332 2327 344 2339 sw
rect 833 2377 835 2379
rect 863 2377 865 2379
rect 833 2355 865 2377
rect 786 2327 795 2355
rect 825 2327 873 2355
rect 903 2327 912 2355
tri 912 2327 924 2339 sw
rect 1413 2377 1415 2379
rect 1443 2377 1445 2379
rect 1413 2355 1445 2377
rect 1366 2327 1375 2355
rect 1405 2327 1453 2355
rect 1483 2327 1492 2355
tri 1492 2327 1504 2339 sw
rect 1993 2377 1995 2379
rect 2023 2377 2025 2379
rect 1993 2355 2025 2377
rect 1946 2327 1955 2355
rect 1985 2327 2033 2355
rect 2063 2327 2072 2355
tri 2072 2327 2084 2339 sw
rect 2573 2377 2575 2379
rect 2603 2377 2605 2379
rect 2573 2355 2605 2377
rect 2526 2327 2535 2355
rect 2565 2327 2613 2355
rect 2643 2327 2652 2355
tri 2652 2327 2664 2339 sw
rect 3153 2377 3155 2379
rect 3183 2377 3185 2379
rect 3153 2355 3185 2377
rect 3106 2327 3115 2355
rect 3145 2327 3193 2355
rect 3223 2327 3232 2355
tri 3232 2327 3244 2339 sw
rect 3733 2377 3735 2379
rect 3763 2377 3765 2379
rect 3733 2355 3765 2377
rect 3686 2327 3695 2355
rect 3725 2327 3773 2355
rect 3803 2327 3812 2355
tri 3812 2327 3824 2339 sw
rect 4313 2377 4315 2379
rect 4343 2377 4345 2379
rect 4313 2355 4345 2377
rect 4266 2327 4275 2355
rect 4305 2327 4353 2355
rect 4383 2327 4392 2355
tri 4392 2327 4404 2339 sw
rect 4893 2377 4895 2379
rect 4923 2377 4925 2379
rect 4893 2355 4925 2377
rect 4846 2327 4855 2355
rect 4885 2327 4933 2355
rect 4963 2327 4972 2355
tri 4972 2327 4984 2339 sw
rect 5473 2377 5475 2379
rect 5503 2377 5505 2379
rect 5473 2355 5505 2377
rect 5426 2327 5435 2355
rect 5465 2327 5513 2355
rect 5543 2327 5552 2355
tri 5552 2327 5564 2339 sw
rect 6053 2377 6055 2379
rect 6083 2377 6085 2379
rect 6053 2355 6085 2377
rect 6006 2327 6015 2355
rect 6045 2327 6093 2355
rect 6123 2327 6132 2355
tri 6132 2327 6144 2339 sw
rect 6633 2377 6635 2379
rect 6663 2377 6665 2379
rect 6633 2355 6665 2377
rect 6586 2327 6595 2355
rect 6625 2327 6673 2355
rect 6703 2327 6712 2355
tri 6712 2327 6724 2339 sw
rect 253 2107 255 2109
rect 283 2107 285 2109
rect 253 2085 285 2107
rect 206 2057 215 2085
rect 245 2057 293 2085
rect 323 2057 332 2085
tri 332 2057 344 2069 sw
rect 833 2107 835 2109
rect 863 2107 865 2109
rect 833 2085 865 2107
rect 786 2057 795 2085
rect 825 2057 873 2085
rect 903 2057 912 2085
tri 912 2057 924 2069 sw
rect 1413 2107 1415 2109
rect 1443 2107 1445 2109
rect 1413 2085 1445 2107
rect 1366 2057 1375 2085
rect 1405 2057 1453 2085
rect 1483 2057 1492 2085
tri 1492 2057 1504 2069 sw
rect 1993 2107 1995 2109
rect 2023 2107 2025 2109
rect 1993 2085 2025 2107
rect 1946 2057 1955 2085
rect 1985 2057 2033 2085
rect 2063 2057 2072 2085
tri 2072 2057 2084 2069 sw
rect 2573 2107 2575 2109
rect 2603 2107 2605 2109
rect 2573 2085 2605 2107
rect 2526 2057 2535 2085
rect 2565 2057 2613 2085
rect 2643 2057 2652 2085
tri 2652 2057 2664 2069 sw
rect 3153 2107 3155 2109
rect 3183 2107 3185 2109
rect 3153 2085 3185 2107
rect 3106 2057 3115 2085
rect 3145 2057 3193 2085
rect 3223 2057 3232 2085
tri 3232 2057 3244 2069 sw
rect 3733 2107 3735 2109
rect 3763 2107 3765 2109
rect 3733 2085 3765 2107
rect 3686 2057 3695 2085
rect 3725 2057 3773 2085
rect 3803 2057 3812 2085
tri 3812 2057 3824 2069 sw
rect 4313 2107 4315 2109
rect 4343 2107 4345 2109
rect 4313 2085 4345 2107
rect 4266 2057 4275 2085
rect 4305 2057 4353 2085
rect 4383 2057 4392 2085
tri 4392 2057 4404 2069 sw
rect 4893 2107 4895 2109
rect 4923 2107 4925 2109
rect 4893 2085 4925 2107
rect 4846 2057 4855 2085
rect 4885 2057 4933 2085
rect 4963 2057 4972 2085
tri 4972 2057 4984 2069 sw
rect 5473 2107 5475 2109
rect 5503 2107 5505 2109
rect 5473 2085 5505 2107
rect 5426 2057 5435 2085
rect 5465 2057 5513 2085
rect 5543 2057 5552 2085
tri 5552 2057 5564 2069 sw
rect 6053 2107 6055 2109
rect 6083 2107 6085 2109
rect 6053 2085 6085 2107
rect 6006 2057 6015 2085
rect 6045 2057 6093 2085
rect 6123 2057 6132 2085
tri 6132 2057 6144 2069 sw
rect 6633 2107 6635 2109
rect 6663 2107 6665 2109
rect 6633 2085 6665 2107
rect 6586 2057 6595 2085
rect 6625 2057 6673 2085
rect 6703 2057 6712 2085
tri 6712 2057 6724 2069 sw
rect 253 1837 255 1839
rect 283 1837 285 1839
rect 253 1815 285 1837
rect 206 1787 215 1815
rect 245 1787 293 1815
rect 323 1787 332 1815
tri 332 1787 344 1799 sw
rect 833 1837 835 1839
rect 863 1837 865 1839
rect 833 1815 865 1837
rect 786 1787 795 1815
rect 825 1787 873 1815
rect 903 1787 912 1815
tri 912 1787 924 1799 sw
rect 1413 1837 1415 1839
rect 1443 1837 1445 1839
rect 1413 1815 1445 1837
rect 1366 1787 1375 1815
rect 1405 1787 1453 1815
rect 1483 1787 1492 1815
tri 1492 1787 1504 1799 sw
rect 1993 1837 1995 1839
rect 2023 1837 2025 1839
rect 1993 1815 2025 1837
rect 1946 1787 1955 1815
rect 1985 1787 2033 1815
rect 2063 1787 2072 1815
tri 2072 1787 2084 1799 sw
rect 2573 1837 2575 1839
rect 2603 1837 2605 1839
rect 2573 1815 2605 1837
rect 2526 1787 2535 1815
rect 2565 1787 2613 1815
rect 2643 1787 2652 1815
tri 2652 1787 2664 1799 sw
rect 3153 1837 3155 1839
rect 3183 1837 3185 1839
rect 3153 1815 3185 1837
rect 3106 1787 3115 1815
rect 3145 1787 3193 1815
rect 3223 1787 3232 1815
tri 3232 1787 3244 1799 sw
rect 3733 1837 3735 1839
rect 3763 1837 3765 1839
rect 3733 1815 3765 1837
rect 3686 1787 3695 1815
rect 3725 1787 3773 1815
rect 3803 1787 3812 1815
tri 3812 1787 3824 1799 sw
rect 4313 1837 4315 1839
rect 4343 1837 4345 1839
rect 4313 1815 4345 1837
rect 4266 1787 4275 1815
rect 4305 1787 4353 1815
rect 4383 1787 4392 1815
tri 4392 1787 4404 1799 sw
rect 4893 1837 4895 1839
rect 4923 1837 4925 1839
rect 4893 1815 4925 1837
rect 4846 1787 4855 1815
rect 4885 1787 4933 1815
rect 4963 1787 4972 1815
tri 4972 1787 4984 1799 sw
rect 5473 1837 5475 1839
rect 5503 1837 5505 1839
rect 5473 1815 5505 1837
rect 5426 1787 5435 1815
rect 5465 1787 5513 1815
rect 5543 1787 5552 1815
tri 5552 1787 5564 1799 sw
rect 6053 1837 6055 1839
rect 6083 1837 6085 1839
rect 6053 1815 6085 1837
rect 6006 1787 6015 1815
rect 6045 1787 6093 1815
rect 6123 1787 6132 1815
tri 6132 1787 6144 1799 sw
rect 6633 1837 6635 1839
rect 6663 1837 6665 1839
rect 6633 1815 6665 1837
rect 6586 1787 6595 1815
rect 6625 1787 6673 1815
rect 6703 1787 6712 1815
tri 6712 1787 6724 1799 sw
rect 253 1567 255 1569
rect 283 1567 285 1569
rect 253 1545 285 1567
rect 206 1517 215 1545
rect 245 1517 293 1545
rect 323 1517 332 1545
tri 332 1517 344 1529 sw
rect 833 1567 835 1569
rect 863 1567 865 1569
rect 833 1545 865 1567
rect 786 1517 795 1545
rect 825 1517 873 1545
rect 903 1517 912 1545
tri 912 1517 924 1529 sw
rect 1413 1567 1415 1569
rect 1443 1567 1445 1569
rect 1413 1545 1445 1567
rect 1366 1517 1375 1545
rect 1405 1517 1453 1545
rect 1483 1517 1492 1545
tri 1492 1517 1504 1529 sw
rect 1993 1567 1995 1569
rect 2023 1567 2025 1569
rect 1993 1545 2025 1567
rect 1946 1517 1955 1545
rect 1985 1517 2033 1545
rect 2063 1517 2072 1545
tri 2072 1517 2084 1529 sw
rect 2573 1567 2575 1569
rect 2603 1567 2605 1569
rect 2573 1545 2605 1567
rect 2526 1517 2535 1545
rect 2565 1517 2613 1545
rect 2643 1517 2652 1545
tri 2652 1517 2664 1529 sw
rect 3153 1567 3155 1569
rect 3183 1567 3185 1569
rect 3153 1545 3185 1567
rect 3106 1517 3115 1545
rect 3145 1517 3193 1545
rect 3223 1517 3232 1545
tri 3232 1517 3244 1529 sw
rect 3733 1567 3735 1569
rect 3763 1567 3765 1569
rect 3733 1545 3765 1567
rect 3686 1517 3695 1545
rect 3725 1517 3773 1545
rect 3803 1517 3812 1545
tri 3812 1517 3824 1529 sw
rect 4313 1567 4315 1569
rect 4343 1567 4345 1569
rect 4313 1545 4345 1567
rect 4266 1517 4275 1545
rect 4305 1517 4353 1545
rect 4383 1517 4392 1545
tri 4392 1517 4404 1529 sw
rect 4893 1567 4895 1569
rect 4923 1567 4925 1569
rect 4893 1545 4925 1567
rect 4846 1517 4855 1545
rect 4885 1517 4933 1545
rect 4963 1517 4972 1545
tri 4972 1517 4984 1529 sw
rect 5473 1567 5475 1569
rect 5503 1567 5505 1569
rect 5473 1545 5505 1567
rect 5426 1517 5435 1545
rect 5465 1517 5513 1545
rect 5543 1517 5552 1545
tri 5552 1517 5564 1529 sw
rect 6053 1567 6055 1569
rect 6083 1567 6085 1569
rect 6053 1545 6085 1567
rect 6006 1517 6015 1545
rect 6045 1517 6093 1545
rect 6123 1517 6132 1545
tri 6132 1517 6144 1529 sw
rect 6633 1567 6635 1569
rect 6663 1567 6665 1569
rect 6633 1545 6665 1567
rect 6586 1517 6595 1545
rect 6625 1517 6673 1545
rect 6703 1517 6712 1545
tri 6712 1517 6724 1529 sw
rect 253 1297 255 1299
rect 283 1297 285 1299
rect 253 1275 285 1297
rect 206 1247 215 1275
rect 245 1247 293 1275
rect 323 1247 332 1275
tri 332 1247 344 1259 sw
rect 833 1297 835 1299
rect 863 1297 865 1299
rect 833 1275 865 1297
rect 786 1247 795 1275
rect 825 1247 873 1275
rect 903 1247 912 1275
tri 912 1247 924 1259 sw
rect 1413 1297 1415 1299
rect 1443 1297 1445 1299
rect 1413 1275 1445 1297
rect 1366 1247 1375 1275
rect 1405 1247 1453 1275
rect 1483 1247 1492 1275
tri 1492 1247 1504 1259 sw
rect 1993 1297 1995 1299
rect 2023 1297 2025 1299
rect 1993 1275 2025 1297
rect 1946 1247 1955 1275
rect 1985 1247 2033 1275
rect 2063 1247 2072 1275
tri 2072 1247 2084 1259 sw
rect 2573 1297 2575 1299
rect 2603 1297 2605 1299
rect 2573 1275 2605 1297
rect 2526 1247 2535 1275
rect 2565 1247 2613 1275
rect 2643 1247 2652 1275
tri 2652 1247 2664 1259 sw
rect 3153 1297 3155 1299
rect 3183 1297 3185 1299
rect 3153 1275 3185 1297
rect 3106 1247 3115 1275
rect 3145 1247 3193 1275
rect 3223 1247 3232 1275
tri 3232 1247 3244 1259 sw
rect 3733 1297 3735 1299
rect 3763 1297 3765 1299
rect 3733 1275 3765 1297
rect 3686 1247 3695 1275
rect 3725 1247 3773 1275
rect 3803 1247 3812 1275
tri 3812 1247 3824 1259 sw
rect 4313 1297 4315 1299
rect 4343 1297 4345 1299
rect 4313 1275 4345 1297
rect 4266 1247 4275 1275
rect 4305 1247 4353 1275
rect 4383 1247 4392 1275
tri 4392 1247 4404 1259 sw
rect 4893 1297 4895 1299
rect 4923 1297 4925 1299
rect 4893 1275 4925 1297
rect 4846 1247 4855 1275
rect 4885 1247 4933 1275
rect 4963 1247 4972 1275
tri 4972 1247 4984 1259 sw
rect 5473 1297 5475 1299
rect 5503 1297 5505 1299
rect 5473 1275 5505 1297
rect 5426 1247 5435 1275
rect 5465 1247 5513 1275
rect 5543 1247 5552 1275
tri 5552 1247 5564 1259 sw
rect 6053 1297 6055 1299
rect 6083 1297 6085 1299
rect 6053 1275 6085 1297
rect 6006 1247 6015 1275
rect 6045 1247 6093 1275
rect 6123 1247 6132 1275
tri 6132 1247 6144 1259 sw
rect 6633 1297 6635 1299
rect 6663 1297 6665 1299
rect 6633 1275 6665 1297
rect 6586 1247 6595 1275
rect 6625 1247 6673 1275
rect 6703 1247 6712 1275
tri 6712 1247 6724 1259 sw
rect 253 1027 255 1029
rect 283 1027 285 1029
rect 253 1005 285 1027
rect 206 977 215 1005
rect 245 977 293 1005
rect 323 977 332 1005
tri 332 977 344 989 sw
rect 833 1027 835 1029
rect 863 1027 865 1029
rect 833 1005 865 1027
rect 786 977 795 1005
rect 825 977 873 1005
rect 903 977 912 1005
tri 912 977 924 989 sw
rect 1413 1027 1415 1029
rect 1443 1027 1445 1029
rect 1413 1005 1445 1027
rect 1366 977 1375 1005
rect 1405 977 1453 1005
rect 1483 977 1492 1005
tri 1492 977 1504 989 sw
rect 1993 1027 1995 1029
rect 2023 1027 2025 1029
rect 1993 1005 2025 1027
rect 1946 977 1955 1005
rect 1985 977 2033 1005
rect 2063 977 2072 1005
tri 2072 977 2084 989 sw
rect 2573 1027 2575 1029
rect 2603 1027 2605 1029
rect 2573 1005 2605 1027
rect 2526 977 2535 1005
rect 2565 977 2613 1005
rect 2643 977 2652 1005
tri 2652 977 2664 989 sw
rect 3153 1027 3155 1029
rect 3183 1027 3185 1029
rect 3153 1005 3185 1027
rect 3106 977 3115 1005
rect 3145 977 3193 1005
rect 3223 977 3232 1005
tri 3232 977 3244 989 sw
rect 3733 1027 3735 1029
rect 3763 1027 3765 1029
rect 3733 1005 3765 1027
rect 3686 977 3695 1005
rect 3725 977 3773 1005
rect 3803 977 3812 1005
tri 3812 977 3824 989 sw
rect 4313 1027 4315 1029
rect 4343 1027 4345 1029
rect 4313 1005 4345 1027
rect 4266 977 4275 1005
rect 4305 977 4353 1005
rect 4383 977 4392 1005
tri 4392 977 4404 989 sw
rect 4893 1027 4895 1029
rect 4923 1027 4925 1029
rect 4893 1005 4925 1027
rect 4846 977 4855 1005
rect 4885 977 4933 1005
rect 4963 977 4972 1005
tri 4972 977 4984 989 sw
rect 5473 1027 5475 1029
rect 5503 1027 5505 1029
rect 5473 1005 5505 1027
rect 5426 977 5435 1005
rect 5465 977 5513 1005
rect 5543 977 5552 1005
tri 5552 977 5564 989 sw
rect 6053 1027 6055 1029
rect 6083 1027 6085 1029
rect 6053 1005 6085 1027
rect 6006 977 6015 1005
rect 6045 977 6093 1005
rect 6123 977 6132 1005
tri 6132 977 6144 989 sw
rect 6633 1027 6635 1029
rect 6663 1027 6665 1029
rect 6633 1005 6665 1027
rect 6586 977 6595 1005
rect 6625 977 6673 1005
rect 6703 977 6712 1005
tri 6712 977 6724 989 sw
rect 253 757 255 759
rect 283 757 285 759
rect 253 735 285 757
rect 206 707 215 735
rect 245 707 293 735
rect 323 707 332 735
tri 332 707 344 719 sw
rect 833 757 835 759
rect 863 757 865 759
rect 833 735 865 757
rect 786 707 795 735
rect 825 707 873 735
rect 903 707 912 735
tri 912 707 924 719 sw
rect 1413 757 1415 759
rect 1443 757 1445 759
rect 1413 735 1445 757
rect 1366 707 1375 735
rect 1405 707 1453 735
rect 1483 707 1492 735
tri 1492 707 1504 719 sw
rect 1993 757 1995 759
rect 2023 757 2025 759
rect 1993 735 2025 757
rect 1946 707 1955 735
rect 1985 707 2033 735
rect 2063 707 2072 735
tri 2072 707 2084 719 sw
rect 2573 757 2575 759
rect 2603 757 2605 759
rect 2573 735 2605 757
rect 2526 707 2535 735
rect 2565 707 2613 735
rect 2643 707 2652 735
tri 2652 707 2664 719 sw
rect 3153 757 3155 759
rect 3183 757 3185 759
rect 3153 735 3185 757
rect 3106 707 3115 735
rect 3145 707 3193 735
rect 3223 707 3232 735
tri 3232 707 3244 719 sw
rect 3733 757 3735 759
rect 3763 757 3765 759
rect 3733 735 3765 757
rect 3686 707 3695 735
rect 3725 707 3773 735
rect 3803 707 3812 735
tri 3812 707 3824 719 sw
rect 4313 757 4315 759
rect 4343 757 4345 759
rect 4313 735 4345 757
rect 4266 707 4275 735
rect 4305 707 4353 735
rect 4383 707 4392 735
tri 4392 707 4404 719 sw
rect 4893 757 4895 759
rect 4923 757 4925 759
rect 4893 735 4925 757
rect 4846 707 4855 735
rect 4885 707 4933 735
rect 4963 707 4972 735
tri 4972 707 4984 719 sw
rect 5473 757 5475 759
rect 5503 757 5505 759
rect 5473 735 5505 757
rect 5426 707 5435 735
rect 5465 707 5513 735
rect 5543 707 5552 735
tri 5552 707 5564 719 sw
rect 6053 757 6055 759
rect 6083 757 6085 759
rect 6053 735 6085 757
rect 6006 707 6015 735
rect 6045 707 6093 735
rect 6123 707 6132 735
tri 6132 707 6144 719 sw
rect 6633 757 6635 759
rect 6663 757 6665 759
rect 6633 735 6665 757
rect 6586 707 6595 735
rect 6625 707 6673 735
rect 6703 707 6712 735
tri 6712 707 6724 719 sw
rect 253 487 255 489
rect 283 487 285 489
rect 253 465 285 487
rect 206 437 215 465
rect 245 437 293 465
rect 323 437 332 465
tri 332 437 344 449 sw
rect 833 487 835 489
rect 863 487 865 489
rect 833 465 865 487
rect 786 437 795 465
rect 825 437 873 465
rect 903 437 912 465
tri 912 437 924 449 sw
rect 1413 487 1415 489
rect 1443 487 1445 489
rect 1413 465 1445 487
rect 1366 437 1375 465
rect 1405 437 1453 465
rect 1483 437 1492 465
tri 1492 437 1504 449 sw
rect 1993 487 1995 489
rect 2023 487 2025 489
rect 1993 465 2025 487
rect 1946 437 1955 465
rect 1985 437 2033 465
rect 2063 437 2072 465
tri 2072 437 2084 449 sw
rect 2573 487 2575 489
rect 2603 487 2605 489
rect 2573 465 2605 487
rect 2526 437 2535 465
rect 2565 437 2613 465
rect 2643 437 2652 465
tri 2652 437 2664 449 sw
rect 3153 487 3155 489
rect 3183 487 3185 489
rect 3153 465 3185 487
rect 3106 437 3115 465
rect 3145 437 3193 465
rect 3223 437 3232 465
tri 3232 437 3244 449 sw
rect 3733 487 3735 489
rect 3763 487 3765 489
rect 3733 465 3765 487
rect 3686 437 3695 465
rect 3725 437 3773 465
rect 3803 437 3812 465
tri 3812 437 3824 449 sw
rect 4313 487 4315 489
rect 4343 487 4345 489
rect 4313 465 4345 487
rect 4266 437 4275 465
rect 4305 437 4353 465
rect 4383 437 4392 465
tri 4392 437 4404 449 sw
rect 4893 487 4895 489
rect 4923 487 4925 489
rect 4893 465 4925 487
rect 4846 437 4855 465
rect 4885 437 4933 465
rect 4963 437 4972 465
tri 4972 437 4984 449 sw
rect 5473 487 5475 489
rect 5503 487 5505 489
rect 5473 465 5505 487
rect 5426 437 5435 465
rect 5465 437 5513 465
rect 5543 437 5552 465
tri 5552 437 5564 449 sw
rect 6053 487 6055 489
rect 6083 487 6085 489
rect 6053 465 6085 487
rect 6006 437 6015 465
rect 6045 437 6093 465
rect 6123 437 6132 465
tri 6132 437 6144 449 sw
rect 6633 487 6635 489
rect 6663 487 6665 489
rect 6633 465 6665 487
rect 6586 437 6595 465
rect 6625 437 6673 465
rect 6703 437 6712 465
tri 6712 437 6724 449 sw
rect 253 217 255 219
rect 283 217 285 219
rect 253 195 285 217
rect 206 167 215 195
rect 245 167 293 195
rect 323 167 332 195
tri 332 167 344 179 sw
rect 833 217 835 219
rect 863 217 865 219
rect 833 195 865 217
rect 786 167 795 195
rect 825 167 873 195
rect 903 167 912 195
tri 912 167 924 179 sw
rect 1413 217 1415 219
rect 1443 217 1445 219
rect 1413 195 1445 217
rect 1366 167 1375 195
rect 1405 167 1453 195
rect 1483 167 1492 195
tri 1492 167 1504 179 sw
rect 1993 217 1995 219
rect 2023 217 2025 219
rect 1993 195 2025 217
rect 1946 167 1955 195
rect 1985 167 2033 195
rect 2063 167 2072 195
tri 2072 167 2084 179 sw
rect 2573 217 2575 219
rect 2603 217 2605 219
rect 2573 195 2605 217
rect 2526 167 2535 195
rect 2565 167 2613 195
rect 2643 167 2652 195
tri 2652 167 2664 179 sw
rect 3153 217 3155 219
rect 3183 217 3185 219
rect 3153 195 3185 217
rect 3106 167 3115 195
rect 3145 167 3193 195
rect 3223 167 3232 195
tri 3232 167 3244 179 sw
rect 3733 217 3735 219
rect 3763 217 3765 219
rect 3733 195 3765 217
rect 3686 167 3695 195
rect 3725 167 3773 195
rect 3803 167 3812 195
tri 3812 167 3824 179 sw
rect 4313 217 4315 219
rect 4343 217 4345 219
rect 4313 195 4345 217
rect 4266 167 4275 195
rect 4305 167 4353 195
rect 4383 167 4392 195
tri 4392 167 4404 179 sw
rect 4893 217 4895 219
rect 4923 217 4925 219
rect 4893 195 4925 217
rect 4846 167 4855 195
rect 4885 167 4933 195
rect 4963 167 4972 195
tri 4972 167 4984 179 sw
rect 5473 217 5475 219
rect 5503 217 5505 219
rect 5473 195 5505 217
rect 5426 167 5435 195
rect 5465 167 5513 195
rect 5543 167 5552 195
tri 5552 167 5564 179 sw
rect 6053 217 6055 219
rect 6083 217 6085 219
rect 6053 195 6085 217
rect 6006 167 6015 195
rect 6045 167 6093 195
rect 6123 167 6132 195
tri 6132 167 6144 179 sw
rect 6633 217 6635 219
rect 6663 217 6665 219
rect 6633 195 6665 217
rect 6586 167 6595 195
rect 6625 167 6673 195
rect 6703 167 6712 195
tri 6712 167 6724 179 sw
<< ndiffc >>
rect 67 4227 82 4255
rect 148 4227 163 4255
rect 375 4227 390 4255
rect 457 4227 472 4256
rect 647 4227 662 4255
rect 728 4227 743 4255
rect 955 4227 970 4255
rect 1037 4227 1052 4256
rect 1227 4227 1242 4255
rect 1308 4227 1323 4255
rect 1535 4227 1550 4255
rect 1617 4227 1632 4256
rect 1807 4227 1822 4255
rect 1888 4227 1903 4255
rect 2115 4227 2130 4255
rect 2197 4227 2212 4256
rect 2387 4227 2402 4255
rect 2468 4227 2483 4255
rect 2695 4227 2710 4255
rect 2777 4227 2792 4256
rect 2967 4227 2982 4255
rect 3048 4227 3063 4255
rect 3275 4227 3290 4255
rect 3357 4227 3372 4256
rect 3547 4227 3562 4255
rect 3628 4227 3643 4255
rect 3855 4227 3870 4255
rect 3937 4227 3952 4256
rect 4127 4227 4142 4255
rect 4208 4227 4223 4255
rect 4435 4227 4450 4255
rect 4517 4227 4532 4256
rect 4707 4227 4722 4255
rect 4788 4227 4803 4255
rect 5015 4227 5030 4255
rect 5097 4227 5112 4256
rect 5287 4227 5302 4255
rect 5368 4227 5383 4255
rect 5595 4227 5610 4255
rect 5677 4227 5692 4256
rect 5867 4227 5882 4255
rect 5948 4227 5963 4255
rect 6175 4227 6190 4255
rect 6257 4227 6272 4256
rect 6447 4227 6462 4255
rect 6528 4227 6543 4255
rect 6755 4227 6770 4255
rect 6837 4227 6852 4256
rect -7 4081 8 4123
rect 190 4106 200 4113
tri 200 4106 207 4113 sw
rect 190 4081 207 4106
rect 331 4081 348 4113
rect 530 4081 545 4123
rect 573 4081 588 4123
rect 770 4106 780 4113
tri 780 4106 787 4113 sw
rect 770 4081 787 4106
rect 911 4081 928 4113
rect 1110 4081 1125 4123
rect 1153 4081 1168 4123
rect 1350 4106 1360 4113
tri 1360 4106 1367 4113 sw
rect 1350 4081 1367 4106
rect 1491 4081 1508 4113
rect 1690 4081 1705 4123
rect 1733 4081 1748 4123
rect 1930 4106 1940 4113
tri 1940 4106 1947 4113 sw
rect 1930 4081 1947 4106
rect 2071 4081 2088 4113
rect 2270 4081 2285 4123
rect 2313 4081 2328 4123
rect 2510 4106 2520 4113
tri 2520 4106 2527 4113 sw
rect 2510 4081 2527 4106
rect 2651 4081 2668 4113
rect 2850 4081 2865 4123
rect 2893 4081 2908 4123
rect 3090 4106 3100 4113
tri 3100 4106 3107 4113 sw
rect 3090 4081 3107 4106
rect 3231 4081 3248 4113
rect 3430 4081 3445 4123
rect 3473 4081 3488 4123
rect 3670 4106 3680 4113
tri 3680 4106 3687 4113 sw
rect 3670 4081 3687 4106
rect 3811 4081 3828 4113
rect 4010 4081 4025 4123
rect 4053 4081 4068 4123
rect 4250 4106 4260 4113
tri 4260 4106 4267 4113 sw
rect 4250 4081 4267 4106
rect 4391 4081 4408 4113
rect 4590 4081 4605 4123
rect 4633 4081 4648 4123
rect 4830 4106 4840 4113
tri 4840 4106 4847 4113 sw
rect 4830 4081 4847 4106
rect 4971 4081 4988 4113
rect 5170 4081 5185 4123
rect 5213 4081 5228 4123
rect 5410 4106 5420 4113
tri 5420 4106 5427 4113 sw
rect 5410 4081 5427 4106
rect 5551 4081 5568 4113
rect 5750 4081 5765 4123
rect 5793 4081 5808 4123
rect 5990 4106 6000 4113
tri 6000 4106 6007 4113 sw
rect 5990 4081 6007 4106
rect 6131 4081 6148 4113
rect 6330 4081 6345 4123
rect 6373 4081 6388 4123
rect 6570 4106 6580 4113
tri 6580 4106 6587 4113 sw
rect 6570 4081 6587 4106
rect 6711 4081 6728 4113
rect 6910 4081 6925 4123
rect 253 4043 285 4057
rect 833 4043 865 4057
rect 1413 4043 1445 4057
rect 1993 4043 2025 4057
rect 2573 4043 2605 4057
rect 3153 4043 3185 4057
rect 3733 4043 3765 4057
rect 4313 4043 4345 4057
rect 4893 4043 4925 4057
rect 5473 4043 5505 4057
rect 6053 4043 6085 4057
rect 6633 4043 6665 4057
rect 67 3957 82 3985
rect 148 3957 163 3985
rect 375 3957 390 3985
rect 457 3957 472 3986
rect 647 3957 662 3985
rect 728 3957 743 3985
rect 955 3957 970 3985
rect 1037 3957 1052 3986
rect 1227 3957 1242 3985
rect 1308 3957 1323 3985
rect 1535 3957 1550 3985
rect 1617 3957 1632 3986
rect 1807 3957 1822 3985
rect 1888 3957 1903 3985
rect 2115 3957 2130 3985
rect 2197 3957 2212 3986
rect 2387 3957 2402 3985
rect 2468 3957 2483 3985
rect 2695 3957 2710 3985
rect 2777 3957 2792 3986
rect 2967 3957 2982 3985
rect 3048 3957 3063 3985
rect 3275 3957 3290 3985
rect 3357 3957 3372 3986
rect 3547 3957 3562 3985
rect 3628 3957 3643 3985
rect 3855 3957 3870 3985
rect 3937 3957 3952 3986
rect 4127 3957 4142 3985
rect 4208 3957 4223 3985
rect 4435 3957 4450 3985
rect 4517 3957 4532 3986
rect 4707 3957 4722 3985
rect 4788 3957 4803 3985
rect 5015 3957 5030 3985
rect 5097 3957 5112 3986
rect 5287 3957 5302 3985
rect 5368 3957 5383 3985
rect 5595 3957 5610 3985
rect 5677 3957 5692 3986
rect 5867 3957 5882 3985
rect 5948 3957 5963 3985
rect 6175 3957 6190 3985
rect 6257 3957 6272 3986
rect 6447 3957 6462 3985
rect 6528 3957 6543 3985
rect 6755 3957 6770 3985
rect 6837 3957 6852 3986
rect -7 3811 8 3853
rect 190 3836 200 3843
tri 200 3836 207 3843 sw
rect 190 3811 207 3836
rect 331 3811 348 3843
rect 530 3811 545 3853
rect 573 3811 588 3853
rect 770 3836 780 3843
tri 780 3836 787 3843 sw
rect 770 3811 787 3836
rect 911 3811 928 3843
rect 1110 3811 1125 3853
rect 1153 3811 1168 3853
rect 1350 3836 1360 3843
tri 1360 3836 1367 3843 sw
rect 1350 3811 1367 3836
rect 1491 3811 1508 3843
rect 1690 3811 1705 3853
rect 1733 3811 1748 3853
rect 1930 3836 1940 3843
tri 1940 3836 1947 3843 sw
rect 1930 3811 1947 3836
rect 2071 3811 2088 3843
rect 2270 3811 2285 3853
rect 2313 3811 2328 3853
rect 2510 3836 2520 3843
tri 2520 3836 2527 3843 sw
rect 2510 3811 2527 3836
rect 2651 3811 2668 3843
rect 2850 3811 2865 3853
rect 2893 3811 2908 3853
rect 3090 3836 3100 3843
tri 3100 3836 3107 3843 sw
rect 3090 3811 3107 3836
rect 3231 3811 3248 3843
rect 3430 3811 3445 3853
rect 3473 3811 3488 3853
rect 3670 3836 3680 3843
tri 3680 3836 3687 3843 sw
rect 3670 3811 3687 3836
rect 3811 3811 3828 3843
rect 4010 3811 4025 3853
rect 4053 3811 4068 3853
rect 4250 3836 4260 3843
tri 4260 3836 4267 3843 sw
rect 4250 3811 4267 3836
rect 4391 3811 4408 3843
rect 4590 3811 4605 3853
rect 4633 3811 4648 3853
rect 4830 3836 4840 3843
tri 4840 3836 4847 3843 sw
rect 4830 3811 4847 3836
rect 4971 3811 4988 3843
rect 5170 3811 5185 3853
rect 5213 3811 5228 3853
rect 5410 3836 5420 3843
tri 5420 3836 5427 3843 sw
rect 5410 3811 5427 3836
rect 5551 3811 5568 3843
rect 5750 3811 5765 3853
rect 5793 3811 5808 3853
rect 5990 3836 6000 3843
tri 6000 3836 6007 3843 sw
rect 5990 3811 6007 3836
rect 6131 3811 6148 3843
rect 6330 3811 6345 3853
rect 6373 3811 6388 3853
rect 6570 3836 6580 3843
tri 6580 3836 6587 3843 sw
rect 6570 3811 6587 3836
rect 6711 3811 6728 3843
rect 6910 3811 6925 3853
rect 253 3773 285 3787
rect 833 3773 865 3787
rect 1413 3773 1445 3787
rect 1993 3773 2025 3787
rect 2573 3773 2605 3787
rect 3153 3773 3185 3787
rect 3733 3773 3765 3787
rect 4313 3773 4345 3787
rect 4893 3773 4925 3787
rect 5473 3773 5505 3787
rect 6053 3773 6085 3787
rect 6633 3773 6665 3787
rect 67 3687 82 3715
rect 148 3687 163 3715
rect 375 3687 390 3715
rect 457 3687 472 3716
rect 647 3687 662 3715
rect 728 3687 743 3715
rect 955 3687 970 3715
rect 1037 3687 1052 3716
rect 1227 3687 1242 3715
rect 1308 3687 1323 3715
rect 1535 3687 1550 3715
rect 1617 3687 1632 3716
rect 1807 3687 1822 3715
rect 1888 3687 1903 3715
rect 2115 3687 2130 3715
rect 2197 3687 2212 3716
rect 2387 3687 2402 3715
rect 2468 3687 2483 3715
rect 2695 3687 2710 3715
rect 2777 3687 2792 3716
rect 2967 3687 2982 3715
rect 3048 3687 3063 3715
rect 3275 3687 3290 3715
rect 3357 3687 3372 3716
rect 3547 3687 3562 3715
rect 3628 3687 3643 3715
rect 3855 3687 3870 3715
rect 3937 3687 3952 3716
rect 4127 3687 4142 3715
rect 4208 3687 4223 3715
rect 4435 3687 4450 3715
rect 4517 3687 4532 3716
rect 4707 3687 4722 3715
rect 4788 3687 4803 3715
rect 5015 3687 5030 3715
rect 5097 3687 5112 3716
rect 5287 3687 5302 3715
rect 5368 3687 5383 3715
rect 5595 3687 5610 3715
rect 5677 3687 5692 3716
rect 5867 3687 5882 3715
rect 5948 3687 5963 3715
rect 6175 3687 6190 3715
rect 6257 3687 6272 3716
rect 6447 3687 6462 3715
rect 6528 3687 6543 3715
rect 6755 3687 6770 3715
rect 6837 3687 6852 3716
rect -7 3541 8 3583
rect 190 3566 200 3573
tri 200 3566 207 3573 sw
rect 190 3541 207 3566
rect 331 3541 348 3573
rect 530 3541 545 3583
rect 573 3541 588 3583
rect 770 3566 780 3573
tri 780 3566 787 3573 sw
rect 770 3541 787 3566
rect 911 3541 928 3573
rect 1110 3541 1125 3583
rect 1153 3541 1168 3583
rect 1350 3566 1360 3573
tri 1360 3566 1367 3573 sw
rect 1350 3541 1367 3566
rect 1491 3541 1508 3573
rect 1690 3541 1705 3583
rect 1733 3541 1748 3583
rect 1930 3566 1940 3573
tri 1940 3566 1947 3573 sw
rect 1930 3541 1947 3566
rect 2071 3541 2088 3573
rect 2270 3541 2285 3583
rect 2313 3541 2328 3583
rect 2510 3566 2520 3573
tri 2520 3566 2527 3573 sw
rect 2510 3541 2527 3566
rect 2651 3541 2668 3573
rect 2850 3541 2865 3583
rect 2893 3541 2908 3583
rect 3090 3566 3100 3573
tri 3100 3566 3107 3573 sw
rect 3090 3541 3107 3566
rect 3231 3541 3248 3573
rect 3430 3541 3445 3583
rect 3473 3541 3488 3583
rect 3670 3566 3680 3573
tri 3680 3566 3687 3573 sw
rect 3670 3541 3687 3566
rect 3811 3541 3828 3573
rect 4010 3541 4025 3583
rect 4053 3541 4068 3583
rect 4250 3566 4260 3573
tri 4260 3566 4267 3573 sw
rect 4250 3541 4267 3566
rect 4391 3541 4408 3573
rect 4590 3541 4605 3583
rect 4633 3541 4648 3583
rect 4830 3566 4840 3573
tri 4840 3566 4847 3573 sw
rect 4830 3541 4847 3566
rect 4971 3541 4988 3573
rect 5170 3541 5185 3583
rect 5213 3541 5228 3583
rect 5410 3566 5420 3573
tri 5420 3566 5427 3573 sw
rect 5410 3541 5427 3566
rect 5551 3541 5568 3573
rect 5750 3541 5765 3583
rect 5793 3541 5808 3583
rect 5990 3566 6000 3573
tri 6000 3566 6007 3573 sw
rect 5990 3541 6007 3566
rect 6131 3541 6148 3573
rect 6330 3541 6345 3583
rect 6373 3541 6388 3583
rect 6570 3566 6580 3573
tri 6580 3566 6587 3573 sw
rect 6570 3541 6587 3566
rect 6711 3541 6728 3573
rect 6910 3541 6925 3583
rect 253 3503 285 3517
rect 833 3503 865 3517
rect 1413 3503 1445 3517
rect 1993 3503 2025 3517
rect 2573 3503 2605 3517
rect 3153 3503 3185 3517
rect 3733 3503 3765 3517
rect 4313 3503 4345 3517
rect 4893 3503 4925 3517
rect 5473 3503 5505 3517
rect 6053 3503 6085 3517
rect 6633 3503 6665 3517
rect 67 3417 82 3445
rect 148 3417 163 3445
rect 375 3417 390 3445
rect 457 3417 472 3446
rect 647 3417 662 3445
rect 728 3417 743 3445
rect 955 3417 970 3445
rect 1037 3417 1052 3446
rect 1227 3417 1242 3445
rect 1308 3417 1323 3445
rect 1535 3417 1550 3445
rect 1617 3417 1632 3446
rect 1807 3417 1822 3445
rect 1888 3417 1903 3445
rect 2115 3417 2130 3445
rect 2197 3417 2212 3446
rect 2387 3417 2402 3445
rect 2468 3417 2483 3445
rect 2695 3417 2710 3445
rect 2777 3417 2792 3446
rect 2967 3417 2982 3445
rect 3048 3417 3063 3445
rect 3275 3417 3290 3445
rect 3357 3417 3372 3446
rect 3547 3417 3562 3445
rect 3628 3417 3643 3445
rect 3855 3417 3870 3445
rect 3937 3417 3952 3446
rect 4127 3417 4142 3445
rect 4208 3417 4223 3445
rect 4435 3417 4450 3445
rect 4517 3417 4532 3446
rect 4707 3417 4722 3445
rect 4788 3417 4803 3445
rect 5015 3417 5030 3445
rect 5097 3417 5112 3446
rect 5287 3417 5302 3445
rect 5368 3417 5383 3445
rect 5595 3417 5610 3445
rect 5677 3417 5692 3446
rect 5867 3417 5882 3445
rect 5948 3417 5963 3445
rect 6175 3417 6190 3445
rect 6257 3417 6272 3446
rect 6447 3417 6462 3445
rect 6528 3417 6543 3445
rect 6755 3417 6770 3445
rect 6837 3417 6852 3446
rect -7 3271 8 3313
rect 190 3296 200 3303
tri 200 3296 207 3303 sw
rect 190 3271 207 3296
rect 331 3271 348 3303
rect 530 3271 545 3313
rect 573 3271 588 3313
rect 770 3296 780 3303
tri 780 3296 787 3303 sw
rect 770 3271 787 3296
rect 911 3271 928 3303
rect 1110 3271 1125 3313
rect 1153 3271 1168 3313
rect 1350 3296 1360 3303
tri 1360 3296 1367 3303 sw
rect 1350 3271 1367 3296
rect 1491 3271 1508 3303
rect 1690 3271 1705 3313
rect 1733 3271 1748 3313
rect 1930 3296 1940 3303
tri 1940 3296 1947 3303 sw
rect 1930 3271 1947 3296
rect 2071 3271 2088 3303
rect 2270 3271 2285 3313
rect 2313 3271 2328 3313
rect 2510 3296 2520 3303
tri 2520 3296 2527 3303 sw
rect 2510 3271 2527 3296
rect 2651 3271 2668 3303
rect 2850 3271 2865 3313
rect 2893 3271 2908 3313
rect 3090 3296 3100 3303
tri 3100 3296 3107 3303 sw
rect 3090 3271 3107 3296
rect 3231 3271 3248 3303
rect 3430 3271 3445 3313
rect 3473 3271 3488 3313
rect 3670 3296 3680 3303
tri 3680 3296 3687 3303 sw
rect 3670 3271 3687 3296
rect 3811 3271 3828 3303
rect 4010 3271 4025 3313
rect 4053 3271 4068 3313
rect 4250 3296 4260 3303
tri 4260 3296 4267 3303 sw
rect 4250 3271 4267 3296
rect 4391 3271 4408 3303
rect 4590 3271 4605 3313
rect 4633 3271 4648 3313
rect 4830 3296 4840 3303
tri 4840 3296 4847 3303 sw
rect 4830 3271 4847 3296
rect 4971 3271 4988 3303
rect 5170 3271 5185 3313
rect 5213 3271 5228 3313
rect 5410 3296 5420 3303
tri 5420 3296 5427 3303 sw
rect 5410 3271 5427 3296
rect 5551 3271 5568 3303
rect 5750 3271 5765 3313
rect 5793 3271 5808 3313
rect 5990 3296 6000 3303
tri 6000 3296 6007 3303 sw
rect 5990 3271 6007 3296
rect 6131 3271 6148 3303
rect 6330 3271 6345 3313
rect 6373 3271 6388 3313
rect 6570 3296 6580 3303
tri 6580 3296 6587 3303 sw
rect 6570 3271 6587 3296
rect 6711 3271 6728 3303
rect 6910 3271 6925 3313
rect 253 3233 285 3247
rect 833 3233 865 3247
rect 1413 3233 1445 3247
rect 1993 3233 2025 3247
rect 2573 3233 2605 3247
rect 3153 3233 3185 3247
rect 3733 3233 3765 3247
rect 4313 3233 4345 3247
rect 4893 3233 4925 3247
rect 5473 3233 5505 3247
rect 6053 3233 6085 3247
rect 6633 3233 6665 3247
rect 67 3147 82 3175
rect 148 3147 163 3175
rect 375 3147 390 3175
rect 457 3147 472 3176
rect 647 3147 662 3175
rect 728 3147 743 3175
rect 955 3147 970 3175
rect 1037 3147 1052 3176
rect 1227 3147 1242 3175
rect 1308 3147 1323 3175
rect 1535 3147 1550 3175
rect 1617 3147 1632 3176
rect 1807 3147 1822 3175
rect 1888 3147 1903 3175
rect 2115 3147 2130 3175
rect 2197 3147 2212 3176
rect 2387 3147 2402 3175
rect 2468 3147 2483 3175
rect 2695 3147 2710 3175
rect 2777 3147 2792 3176
rect 2967 3147 2982 3175
rect 3048 3147 3063 3175
rect 3275 3147 3290 3175
rect 3357 3147 3372 3176
rect 3547 3147 3562 3175
rect 3628 3147 3643 3175
rect 3855 3147 3870 3175
rect 3937 3147 3952 3176
rect 4127 3147 4142 3175
rect 4208 3147 4223 3175
rect 4435 3147 4450 3175
rect 4517 3147 4532 3176
rect 4707 3147 4722 3175
rect 4788 3147 4803 3175
rect 5015 3147 5030 3175
rect 5097 3147 5112 3176
rect 5287 3147 5302 3175
rect 5368 3147 5383 3175
rect 5595 3147 5610 3175
rect 5677 3147 5692 3176
rect 5867 3147 5882 3175
rect 5948 3147 5963 3175
rect 6175 3147 6190 3175
rect 6257 3147 6272 3176
rect 6447 3147 6462 3175
rect 6528 3147 6543 3175
rect 6755 3147 6770 3175
rect 6837 3147 6852 3176
rect -7 3001 8 3043
rect 190 3026 200 3033
tri 200 3026 207 3033 sw
rect 190 3001 207 3026
rect 331 3001 348 3033
rect 530 3001 545 3043
rect 573 3001 588 3043
rect 770 3026 780 3033
tri 780 3026 787 3033 sw
rect 770 3001 787 3026
rect 911 3001 928 3033
rect 1110 3001 1125 3043
rect 1153 3001 1168 3043
rect 1350 3026 1360 3033
tri 1360 3026 1367 3033 sw
rect 1350 3001 1367 3026
rect 1491 3001 1508 3033
rect 1690 3001 1705 3043
rect 1733 3001 1748 3043
rect 1930 3026 1940 3033
tri 1940 3026 1947 3033 sw
rect 1930 3001 1947 3026
rect 2071 3001 2088 3033
rect 2270 3001 2285 3043
rect 2313 3001 2328 3043
rect 2510 3026 2520 3033
tri 2520 3026 2527 3033 sw
rect 2510 3001 2527 3026
rect 2651 3001 2668 3033
rect 2850 3001 2865 3043
rect 2893 3001 2908 3043
rect 3090 3026 3100 3033
tri 3100 3026 3107 3033 sw
rect 3090 3001 3107 3026
rect 3231 3001 3248 3033
rect 3430 3001 3445 3043
rect 3473 3001 3488 3043
rect 3670 3026 3680 3033
tri 3680 3026 3687 3033 sw
rect 3670 3001 3687 3026
rect 3811 3001 3828 3033
rect 4010 3001 4025 3043
rect 4053 3001 4068 3043
rect 4250 3026 4260 3033
tri 4260 3026 4267 3033 sw
rect 4250 3001 4267 3026
rect 4391 3001 4408 3033
rect 4590 3001 4605 3043
rect 4633 3001 4648 3043
rect 4830 3026 4840 3033
tri 4840 3026 4847 3033 sw
rect 4830 3001 4847 3026
rect 4971 3001 4988 3033
rect 5170 3001 5185 3043
rect 5213 3001 5228 3043
rect 5410 3026 5420 3033
tri 5420 3026 5427 3033 sw
rect 5410 3001 5427 3026
rect 5551 3001 5568 3033
rect 5750 3001 5765 3043
rect 5793 3001 5808 3043
rect 5990 3026 6000 3033
tri 6000 3026 6007 3033 sw
rect 5990 3001 6007 3026
rect 6131 3001 6148 3033
rect 6330 3001 6345 3043
rect 6373 3001 6388 3043
rect 6570 3026 6580 3033
tri 6580 3026 6587 3033 sw
rect 6570 3001 6587 3026
rect 6711 3001 6728 3033
rect 6910 3001 6925 3043
rect 253 2963 285 2977
rect 833 2963 865 2977
rect 1413 2963 1445 2977
rect 1993 2963 2025 2977
rect 2573 2963 2605 2977
rect 3153 2963 3185 2977
rect 3733 2963 3765 2977
rect 4313 2963 4345 2977
rect 4893 2963 4925 2977
rect 5473 2963 5505 2977
rect 6053 2963 6085 2977
rect 6633 2963 6665 2977
rect 67 2877 82 2905
rect 148 2877 163 2905
rect 375 2877 390 2905
rect 457 2877 472 2906
rect 647 2877 662 2905
rect 728 2877 743 2905
rect 955 2877 970 2905
rect 1037 2877 1052 2906
rect 1227 2877 1242 2905
rect 1308 2877 1323 2905
rect 1535 2877 1550 2905
rect 1617 2877 1632 2906
rect 1807 2877 1822 2905
rect 1888 2877 1903 2905
rect 2115 2877 2130 2905
rect 2197 2877 2212 2906
rect 2387 2877 2402 2905
rect 2468 2877 2483 2905
rect 2695 2877 2710 2905
rect 2777 2877 2792 2906
rect 2967 2877 2982 2905
rect 3048 2877 3063 2905
rect 3275 2877 3290 2905
rect 3357 2877 3372 2906
rect 3547 2877 3562 2905
rect 3628 2877 3643 2905
rect 3855 2877 3870 2905
rect 3937 2877 3952 2906
rect 4127 2877 4142 2905
rect 4208 2877 4223 2905
rect 4435 2877 4450 2905
rect 4517 2877 4532 2906
rect 4707 2877 4722 2905
rect 4788 2877 4803 2905
rect 5015 2877 5030 2905
rect 5097 2877 5112 2906
rect 5287 2877 5302 2905
rect 5368 2877 5383 2905
rect 5595 2877 5610 2905
rect 5677 2877 5692 2906
rect 5867 2877 5882 2905
rect 5948 2877 5963 2905
rect 6175 2877 6190 2905
rect 6257 2877 6272 2906
rect 6447 2877 6462 2905
rect 6528 2877 6543 2905
rect 6755 2877 6770 2905
rect 6837 2877 6852 2906
rect -7 2731 8 2773
rect 190 2756 200 2763
tri 200 2756 207 2763 sw
rect 190 2731 207 2756
rect 331 2731 348 2763
rect 530 2731 545 2773
rect 573 2731 588 2773
rect 770 2756 780 2763
tri 780 2756 787 2763 sw
rect 770 2731 787 2756
rect 911 2731 928 2763
rect 1110 2731 1125 2773
rect 1153 2731 1168 2773
rect 1350 2756 1360 2763
tri 1360 2756 1367 2763 sw
rect 1350 2731 1367 2756
rect 1491 2731 1508 2763
rect 1690 2731 1705 2773
rect 1733 2731 1748 2773
rect 1930 2756 1940 2763
tri 1940 2756 1947 2763 sw
rect 1930 2731 1947 2756
rect 2071 2731 2088 2763
rect 2270 2731 2285 2773
rect 2313 2731 2328 2773
rect 2510 2756 2520 2763
tri 2520 2756 2527 2763 sw
rect 2510 2731 2527 2756
rect 2651 2731 2668 2763
rect 2850 2731 2865 2773
rect 2893 2731 2908 2773
rect 3090 2756 3100 2763
tri 3100 2756 3107 2763 sw
rect 3090 2731 3107 2756
rect 3231 2731 3248 2763
rect 3430 2731 3445 2773
rect 3473 2731 3488 2773
rect 3670 2756 3680 2763
tri 3680 2756 3687 2763 sw
rect 3670 2731 3687 2756
rect 3811 2731 3828 2763
rect 4010 2731 4025 2773
rect 4053 2731 4068 2773
rect 4250 2756 4260 2763
tri 4260 2756 4267 2763 sw
rect 4250 2731 4267 2756
rect 4391 2731 4408 2763
rect 4590 2731 4605 2773
rect 4633 2731 4648 2773
rect 4830 2756 4840 2763
tri 4840 2756 4847 2763 sw
rect 4830 2731 4847 2756
rect 4971 2731 4988 2763
rect 5170 2731 5185 2773
rect 5213 2731 5228 2773
rect 5410 2756 5420 2763
tri 5420 2756 5427 2763 sw
rect 5410 2731 5427 2756
rect 5551 2731 5568 2763
rect 5750 2731 5765 2773
rect 5793 2731 5808 2773
rect 5990 2756 6000 2763
tri 6000 2756 6007 2763 sw
rect 5990 2731 6007 2756
rect 6131 2731 6148 2763
rect 6330 2731 6345 2773
rect 6373 2731 6388 2773
rect 6570 2756 6580 2763
tri 6580 2756 6587 2763 sw
rect 6570 2731 6587 2756
rect 6711 2731 6728 2763
rect 6910 2731 6925 2773
rect 253 2693 285 2707
rect 833 2693 865 2707
rect 1413 2693 1445 2707
rect 1993 2693 2025 2707
rect 2573 2693 2605 2707
rect 3153 2693 3185 2707
rect 3733 2693 3765 2707
rect 4313 2693 4345 2707
rect 4893 2693 4925 2707
rect 5473 2693 5505 2707
rect 6053 2693 6085 2707
rect 6633 2693 6665 2707
rect 67 2607 82 2635
rect 148 2607 163 2635
rect 375 2607 390 2635
rect 457 2607 472 2636
rect 647 2607 662 2635
rect 728 2607 743 2635
rect 955 2607 970 2635
rect 1037 2607 1052 2636
rect 1227 2607 1242 2635
rect 1308 2607 1323 2635
rect 1535 2607 1550 2635
rect 1617 2607 1632 2636
rect 1807 2607 1822 2635
rect 1888 2607 1903 2635
rect 2115 2607 2130 2635
rect 2197 2607 2212 2636
rect 2387 2607 2402 2635
rect 2468 2607 2483 2635
rect 2695 2607 2710 2635
rect 2777 2607 2792 2636
rect 2967 2607 2982 2635
rect 3048 2607 3063 2635
rect 3275 2607 3290 2635
rect 3357 2607 3372 2636
rect 3547 2607 3562 2635
rect 3628 2607 3643 2635
rect 3855 2607 3870 2635
rect 3937 2607 3952 2636
rect 4127 2607 4142 2635
rect 4208 2607 4223 2635
rect 4435 2607 4450 2635
rect 4517 2607 4532 2636
rect 4707 2607 4722 2635
rect 4788 2607 4803 2635
rect 5015 2607 5030 2635
rect 5097 2607 5112 2636
rect 5287 2607 5302 2635
rect 5368 2607 5383 2635
rect 5595 2607 5610 2635
rect 5677 2607 5692 2636
rect 5867 2607 5882 2635
rect 5948 2607 5963 2635
rect 6175 2607 6190 2635
rect 6257 2607 6272 2636
rect 6447 2607 6462 2635
rect 6528 2607 6543 2635
rect 6755 2607 6770 2635
rect 6837 2607 6852 2636
rect -7 2461 8 2503
rect 190 2486 200 2493
tri 200 2486 207 2493 sw
rect 190 2461 207 2486
rect 331 2461 348 2493
rect 530 2461 545 2503
rect 573 2461 588 2503
rect 770 2486 780 2493
tri 780 2486 787 2493 sw
rect 770 2461 787 2486
rect 911 2461 928 2493
rect 1110 2461 1125 2503
rect 1153 2461 1168 2503
rect 1350 2486 1360 2493
tri 1360 2486 1367 2493 sw
rect 1350 2461 1367 2486
rect 1491 2461 1508 2493
rect 1690 2461 1705 2503
rect 1733 2461 1748 2503
rect 1930 2486 1940 2493
tri 1940 2486 1947 2493 sw
rect 1930 2461 1947 2486
rect 2071 2461 2088 2493
rect 2270 2461 2285 2503
rect 2313 2461 2328 2503
rect 2510 2486 2520 2493
tri 2520 2486 2527 2493 sw
rect 2510 2461 2527 2486
rect 2651 2461 2668 2493
rect 2850 2461 2865 2503
rect 2893 2461 2908 2503
rect 3090 2486 3100 2493
tri 3100 2486 3107 2493 sw
rect 3090 2461 3107 2486
rect 3231 2461 3248 2493
rect 3430 2461 3445 2503
rect 3473 2461 3488 2503
rect 3670 2486 3680 2493
tri 3680 2486 3687 2493 sw
rect 3670 2461 3687 2486
rect 3811 2461 3828 2493
rect 4010 2461 4025 2503
rect 4053 2461 4068 2503
rect 4250 2486 4260 2493
tri 4260 2486 4267 2493 sw
rect 4250 2461 4267 2486
rect 4391 2461 4408 2493
rect 4590 2461 4605 2503
rect 4633 2461 4648 2503
rect 4830 2486 4840 2493
tri 4840 2486 4847 2493 sw
rect 4830 2461 4847 2486
rect 4971 2461 4988 2493
rect 5170 2461 5185 2503
rect 5213 2461 5228 2503
rect 5410 2486 5420 2493
tri 5420 2486 5427 2493 sw
rect 5410 2461 5427 2486
rect 5551 2461 5568 2493
rect 5750 2461 5765 2503
rect 5793 2461 5808 2503
rect 5990 2486 6000 2493
tri 6000 2486 6007 2493 sw
rect 5990 2461 6007 2486
rect 6131 2461 6148 2493
rect 6330 2461 6345 2503
rect 6373 2461 6388 2503
rect 6570 2486 6580 2493
tri 6580 2486 6587 2493 sw
rect 6570 2461 6587 2486
rect 6711 2461 6728 2493
rect 6910 2461 6925 2503
rect 253 2423 285 2437
rect 833 2423 865 2437
rect 1413 2423 1445 2437
rect 1993 2423 2025 2437
rect 2573 2423 2605 2437
rect 3153 2423 3185 2437
rect 3733 2423 3765 2437
rect 4313 2423 4345 2437
rect 4893 2423 4925 2437
rect 5473 2423 5505 2437
rect 6053 2423 6085 2437
rect 6633 2423 6665 2437
rect 67 2337 82 2365
rect 148 2337 163 2365
rect 375 2337 390 2365
rect 457 2337 472 2366
rect 647 2337 662 2365
rect 728 2337 743 2365
rect 955 2337 970 2365
rect 1037 2337 1052 2366
rect 1227 2337 1242 2365
rect 1308 2337 1323 2365
rect 1535 2337 1550 2365
rect 1617 2337 1632 2366
rect 1807 2337 1822 2365
rect 1888 2337 1903 2365
rect 2115 2337 2130 2365
rect 2197 2337 2212 2366
rect 2387 2337 2402 2365
rect 2468 2337 2483 2365
rect 2695 2337 2710 2365
rect 2777 2337 2792 2366
rect 2967 2337 2982 2365
rect 3048 2337 3063 2365
rect 3275 2337 3290 2365
rect 3357 2337 3372 2366
rect 3547 2337 3562 2365
rect 3628 2337 3643 2365
rect 3855 2337 3870 2365
rect 3937 2337 3952 2366
rect 4127 2337 4142 2365
rect 4208 2337 4223 2365
rect 4435 2337 4450 2365
rect 4517 2337 4532 2366
rect 4707 2337 4722 2365
rect 4788 2337 4803 2365
rect 5015 2337 5030 2365
rect 5097 2337 5112 2366
rect 5287 2337 5302 2365
rect 5368 2337 5383 2365
rect 5595 2337 5610 2365
rect 5677 2337 5692 2366
rect 5867 2337 5882 2365
rect 5948 2337 5963 2365
rect 6175 2337 6190 2365
rect 6257 2337 6272 2366
rect 6447 2337 6462 2365
rect 6528 2337 6543 2365
rect 6755 2337 6770 2365
rect 6837 2337 6852 2366
rect -7 2191 8 2233
rect 190 2216 200 2223
tri 200 2216 207 2223 sw
rect 190 2191 207 2216
rect 331 2191 348 2223
rect 530 2191 545 2233
rect 573 2191 588 2233
rect 770 2216 780 2223
tri 780 2216 787 2223 sw
rect 770 2191 787 2216
rect 911 2191 928 2223
rect 1110 2191 1125 2233
rect 1153 2191 1168 2233
rect 1350 2216 1360 2223
tri 1360 2216 1367 2223 sw
rect 1350 2191 1367 2216
rect 1491 2191 1508 2223
rect 1690 2191 1705 2233
rect 1733 2191 1748 2233
rect 1930 2216 1940 2223
tri 1940 2216 1947 2223 sw
rect 1930 2191 1947 2216
rect 2071 2191 2088 2223
rect 2270 2191 2285 2233
rect 2313 2191 2328 2233
rect 2510 2216 2520 2223
tri 2520 2216 2527 2223 sw
rect 2510 2191 2527 2216
rect 2651 2191 2668 2223
rect 2850 2191 2865 2233
rect 2893 2191 2908 2233
rect 3090 2216 3100 2223
tri 3100 2216 3107 2223 sw
rect 3090 2191 3107 2216
rect 3231 2191 3248 2223
rect 3430 2191 3445 2233
rect 3473 2191 3488 2233
rect 3670 2216 3680 2223
tri 3680 2216 3687 2223 sw
rect 3670 2191 3687 2216
rect 3811 2191 3828 2223
rect 4010 2191 4025 2233
rect 4053 2191 4068 2233
rect 4250 2216 4260 2223
tri 4260 2216 4267 2223 sw
rect 4250 2191 4267 2216
rect 4391 2191 4408 2223
rect 4590 2191 4605 2233
rect 4633 2191 4648 2233
rect 4830 2216 4840 2223
tri 4840 2216 4847 2223 sw
rect 4830 2191 4847 2216
rect 4971 2191 4988 2223
rect 5170 2191 5185 2233
rect 5213 2191 5228 2233
rect 5410 2216 5420 2223
tri 5420 2216 5427 2223 sw
rect 5410 2191 5427 2216
rect 5551 2191 5568 2223
rect 5750 2191 5765 2233
rect 5793 2191 5808 2233
rect 5990 2216 6000 2223
tri 6000 2216 6007 2223 sw
rect 5990 2191 6007 2216
rect 6131 2191 6148 2223
rect 6330 2191 6345 2233
rect 6373 2191 6388 2233
rect 6570 2216 6580 2223
tri 6580 2216 6587 2223 sw
rect 6570 2191 6587 2216
rect 6711 2191 6728 2223
rect 6910 2191 6925 2233
rect 253 2153 285 2167
rect 833 2153 865 2167
rect 1413 2153 1445 2167
rect 1993 2153 2025 2167
rect 2573 2153 2605 2167
rect 3153 2153 3185 2167
rect 3733 2153 3765 2167
rect 4313 2153 4345 2167
rect 4893 2153 4925 2167
rect 5473 2153 5505 2167
rect 6053 2153 6085 2167
rect 6633 2153 6665 2167
rect 67 2067 82 2095
rect 148 2067 163 2095
rect 375 2067 390 2095
rect 457 2067 472 2096
rect 647 2067 662 2095
rect 728 2067 743 2095
rect 955 2067 970 2095
rect 1037 2067 1052 2096
rect 1227 2067 1242 2095
rect 1308 2067 1323 2095
rect 1535 2067 1550 2095
rect 1617 2067 1632 2096
rect 1807 2067 1822 2095
rect 1888 2067 1903 2095
rect 2115 2067 2130 2095
rect 2197 2067 2212 2096
rect 2387 2067 2402 2095
rect 2468 2067 2483 2095
rect 2695 2067 2710 2095
rect 2777 2067 2792 2096
rect 2967 2067 2982 2095
rect 3048 2067 3063 2095
rect 3275 2067 3290 2095
rect 3357 2067 3372 2096
rect 3547 2067 3562 2095
rect 3628 2067 3643 2095
rect 3855 2067 3870 2095
rect 3937 2067 3952 2096
rect 4127 2067 4142 2095
rect 4208 2067 4223 2095
rect 4435 2067 4450 2095
rect 4517 2067 4532 2096
rect 4707 2067 4722 2095
rect 4788 2067 4803 2095
rect 5015 2067 5030 2095
rect 5097 2067 5112 2096
rect 5287 2067 5302 2095
rect 5368 2067 5383 2095
rect 5595 2067 5610 2095
rect 5677 2067 5692 2096
rect 5867 2067 5882 2095
rect 5948 2067 5963 2095
rect 6175 2067 6190 2095
rect 6257 2067 6272 2096
rect 6447 2067 6462 2095
rect 6528 2067 6543 2095
rect 6755 2067 6770 2095
rect 6837 2067 6852 2096
rect -7 1921 8 1963
rect 190 1946 200 1953
tri 200 1946 207 1953 sw
rect 190 1921 207 1946
rect 331 1921 348 1953
rect 530 1921 545 1963
rect 573 1921 588 1963
rect 770 1946 780 1953
tri 780 1946 787 1953 sw
rect 770 1921 787 1946
rect 911 1921 928 1953
rect 1110 1921 1125 1963
rect 1153 1921 1168 1963
rect 1350 1946 1360 1953
tri 1360 1946 1367 1953 sw
rect 1350 1921 1367 1946
rect 1491 1921 1508 1953
rect 1690 1921 1705 1963
rect 1733 1921 1748 1963
rect 1930 1946 1940 1953
tri 1940 1946 1947 1953 sw
rect 1930 1921 1947 1946
rect 2071 1921 2088 1953
rect 2270 1921 2285 1963
rect 2313 1921 2328 1963
rect 2510 1946 2520 1953
tri 2520 1946 2527 1953 sw
rect 2510 1921 2527 1946
rect 2651 1921 2668 1953
rect 2850 1921 2865 1963
rect 2893 1921 2908 1963
rect 3090 1946 3100 1953
tri 3100 1946 3107 1953 sw
rect 3090 1921 3107 1946
rect 3231 1921 3248 1953
rect 3430 1921 3445 1963
rect 3473 1921 3488 1963
rect 3670 1946 3680 1953
tri 3680 1946 3687 1953 sw
rect 3670 1921 3687 1946
rect 3811 1921 3828 1953
rect 4010 1921 4025 1963
rect 4053 1921 4068 1963
rect 4250 1946 4260 1953
tri 4260 1946 4267 1953 sw
rect 4250 1921 4267 1946
rect 4391 1921 4408 1953
rect 4590 1921 4605 1963
rect 4633 1921 4648 1963
rect 4830 1946 4840 1953
tri 4840 1946 4847 1953 sw
rect 4830 1921 4847 1946
rect 4971 1921 4988 1953
rect 5170 1921 5185 1963
rect 5213 1921 5228 1963
rect 5410 1946 5420 1953
tri 5420 1946 5427 1953 sw
rect 5410 1921 5427 1946
rect 5551 1921 5568 1953
rect 5750 1921 5765 1963
rect 5793 1921 5808 1963
rect 5990 1946 6000 1953
tri 6000 1946 6007 1953 sw
rect 5990 1921 6007 1946
rect 6131 1921 6148 1953
rect 6330 1921 6345 1963
rect 6373 1921 6388 1963
rect 6570 1946 6580 1953
tri 6580 1946 6587 1953 sw
rect 6570 1921 6587 1946
rect 6711 1921 6728 1953
rect 6910 1921 6925 1963
rect 253 1883 285 1897
rect 833 1883 865 1897
rect 1413 1883 1445 1897
rect 1993 1883 2025 1897
rect 2573 1883 2605 1897
rect 3153 1883 3185 1897
rect 3733 1883 3765 1897
rect 4313 1883 4345 1897
rect 4893 1883 4925 1897
rect 5473 1883 5505 1897
rect 6053 1883 6085 1897
rect 6633 1883 6665 1897
rect 67 1797 82 1825
rect 148 1797 163 1825
rect 375 1797 390 1825
rect 457 1797 472 1826
rect 647 1797 662 1825
rect 728 1797 743 1825
rect 955 1797 970 1825
rect 1037 1797 1052 1826
rect 1227 1797 1242 1825
rect 1308 1797 1323 1825
rect 1535 1797 1550 1825
rect 1617 1797 1632 1826
rect 1807 1797 1822 1825
rect 1888 1797 1903 1825
rect 2115 1797 2130 1825
rect 2197 1797 2212 1826
rect 2387 1797 2402 1825
rect 2468 1797 2483 1825
rect 2695 1797 2710 1825
rect 2777 1797 2792 1826
rect 2967 1797 2982 1825
rect 3048 1797 3063 1825
rect 3275 1797 3290 1825
rect 3357 1797 3372 1826
rect 3547 1797 3562 1825
rect 3628 1797 3643 1825
rect 3855 1797 3870 1825
rect 3937 1797 3952 1826
rect 4127 1797 4142 1825
rect 4208 1797 4223 1825
rect 4435 1797 4450 1825
rect 4517 1797 4532 1826
rect 4707 1797 4722 1825
rect 4788 1797 4803 1825
rect 5015 1797 5030 1825
rect 5097 1797 5112 1826
rect 5287 1797 5302 1825
rect 5368 1797 5383 1825
rect 5595 1797 5610 1825
rect 5677 1797 5692 1826
rect 5867 1797 5882 1825
rect 5948 1797 5963 1825
rect 6175 1797 6190 1825
rect 6257 1797 6272 1826
rect 6447 1797 6462 1825
rect 6528 1797 6543 1825
rect 6755 1797 6770 1825
rect 6837 1797 6852 1826
rect -7 1651 8 1693
rect 190 1676 200 1683
tri 200 1676 207 1683 sw
rect 190 1651 207 1676
rect 331 1651 348 1683
rect 530 1651 545 1693
rect 573 1651 588 1693
rect 770 1676 780 1683
tri 780 1676 787 1683 sw
rect 770 1651 787 1676
rect 911 1651 928 1683
rect 1110 1651 1125 1693
rect 1153 1651 1168 1693
rect 1350 1676 1360 1683
tri 1360 1676 1367 1683 sw
rect 1350 1651 1367 1676
rect 1491 1651 1508 1683
rect 1690 1651 1705 1693
rect 1733 1651 1748 1693
rect 1930 1676 1940 1683
tri 1940 1676 1947 1683 sw
rect 1930 1651 1947 1676
rect 2071 1651 2088 1683
rect 2270 1651 2285 1693
rect 2313 1651 2328 1693
rect 2510 1676 2520 1683
tri 2520 1676 2527 1683 sw
rect 2510 1651 2527 1676
rect 2651 1651 2668 1683
rect 2850 1651 2865 1693
rect 2893 1651 2908 1693
rect 3090 1676 3100 1683
tri 3100 1676 3107 1683 sw
rect 3090 1651 3107 1676
rect 3231 1651 3248 1683
rect 3430 1651 3445 1693
rect 3473 1651 3488 1693
rect 3670 1676 3680 1683
tri 3680 1676 3687 1683 sw
rect 3670 1651 3687 1676
rect 3811 1651 3828 1683
rect 4010 1651 4025 1693
rect 4053 1651 4068 1693
rect 4250 1676 4260 1683
tri 4260 1676 4267 1683 sw
rect 4250 1651 4267 1676
rect 4391 1651 4408 1683
rect 4590 1651 4605 1693
rect 4633 1651 4648 1693
rect 4830 1676 4840 1683
tri 4840 1676 4847 1683 sw
rect 4830 1651 4847 1676
rect 4971 1651 4988 1683
rect 5170 1651 5185 1693
rect 5213 1651 5228 1693
rect 5410 1676 5420 1683
tri 5420 1676 5427 1683 sw
rect 5410 1651 5427 1676
rect 5551 1651 5568 1683
rect 5750 1651 5765 1693
rect 5793 1651 5808 1693
rect 5990 1676 6000 1683
tri 6000 1676 6007 1683 sw
rect 5990 1651 6007 1676
rect 6131 1651 6148 1683
rect 6330 1651 6345 1693
rect 6373 1651 6388 1693
rect 6570 1676 6580 1683
tri 6580 1676 6587 1683 sw
rect 6570 1651 6587 1676
rect 6711 1651 6728 1683
rect 6910 1651 6925 1693
rect 253 1613 285 1627
rect 833 1613 865 1627
rect 1413 1613 1445 1627
rect 1993 1613 2025 1627
rect 2573 1613 2605 1627
rect 3153 1613 3185 1627
rect 3733 1613 3765 1627
rect 4313 1613 4345 1627
rect 4893 1613 4925 1627
rect 5473 1613 5505 1627
rect 6053 1613 6085 1627
rect 6633 1613 6665 1627
rect 67 1527 82 1555
rect 148 1527 163 1555
rect 375 1527 390 1555
rect 457 1527 472 1556
rect 647 1527 662 1555
rect 728 1527 743 1555
rect 955 1527 970 1555
rect 1037 1527 1052 1556
rect 1227 1527 1242 1555
rect 1308 1527 1323 1555
rect 1535 1527 1550 1555
rect 1617 1527 1632 1556
rect 1807 1527 1822 1555
rect 1888 1527 1903 1555
rect 2115 1527 2130 1555
rect 2197 1527 2212 1556
rect 2387 1527 2402 1555
rect 2468 1527 2483 1555
rect 2695 1527 2710 1555
rect 2777 1527 2792 1556
rect 2967 1527 2982 1555
rect 3048 1527 3063 1555
rect 3275 1527 3290 1555
rect 3357 1527 3372 1556
rect 3547 1527 3562 1555
rect 3628 1527 3643 1555
rect 3855 1527 3870 1555
rect 3937 1527 3952 1556
rect 4127 1527 4142 1555
rect 4208 1527 4223 1555
rect 4435 1527 4450 1555
rect 4517 1527 4532 1556
rect 4707 1527 4722 1555
rect 4788 1527 4803 1555
rect 5015 1527 5030 1555
rect 5097 1527 5112 1556
rect 5287 1527 5302 1555
rect 5368 1527 5383 1555
rect 5595 1527 5610 1555
rect 5677 1527 5692 1556
rect 5867 1527 5882 1555
rect 5948 1527 5963 1555
rect 6175 1527 6190 1555
rect 6257 1527 6272 1556
rect 6447 1527 6462 1555
rect 6528 1527 6543 1555
rect 6755 1527 6770 1555
rect 6837 1527 6852 1556
rect -7 1381 8 1423
rect 190 1406 200 1413
tri 200 1406 207 1413 sw
rect 190 1381 207 1406
rect 331 1381 348 1413
rect 530 1381 545 1423
rect 573 1381 588 1423
rect 770 1406 780 1413
tri 780 1406 787 1413 sw
rect 770 1381 787 1406
rect 911 1381 928 1413
rect 1110 1381 1125 1423
rect 1153 1381 1168 1423
rect 1350 1406 1360 1413
tri 1360 1406 1367 1413 sw
rect 1350 1381 1367 1406
rect 1491 1381 1508 1413
rect 1690 1381 1705 1423
rect 1733 1381 1748 1423
rect 1930 1406 1940 1413
tri 1940 1406 1947 1413 sw
rect 1930 1381 1947 1406
rect 2071 1381 2088 1413
rect 2270 1381 2285 1423
rect 2313 1381 2328 1423
rect 2510 1406 2520 1413
tri 2520 1406 2527 1413 sw
rect 2510 1381 2527 1406
rect 2651 1381 2668 1413
rect 2850 1381 2865 1423
rect 2893 1381 2908 1423
rect 3090 1406 3100 1413
tri 3100 1406 3107 1413 sw
rect 3090 1381 3107 1406
rect 3231 1381 3248 1413
rect 3430 1381 3445 1423
rect 3473 1381 3488 1423
rect 3670 1406 3680 1413
tri 3680 1406 3687 1413 sw
rect 3670 1381 3687 1406
rect 3811 1381 3828 1413
rect 4010 1381 4025 1423
rect 4053 1381 4068 1423
rect 4250 1406 4260 1413
tri 4260 1406 4267 1413 sw
rect 4250 1381 4267 1406
rect 4391 1381 4408 1413
rect 4590 1381 4605 1423
rect 4633 1381 4648 1423
rect 4830 1406 4840 1413
tri 4840 1406 4847 1413 sw
rect 4830 1381 4847 1406
rect 4971 1381 4988 1413
rect 5170 1381 5185 1423
rect 5213 1381 5228 1423
rect 5410 1406 5420 1413
tri 5420 1406 5427 1413 sw
rect 5410 1381 5427 1406
rect 5551 1381 5568 1413
rect 5750 1381 5765 1423
rect 5793 1381 5808 1423
rect 5990 1406 6000 1413
tri 6000 1406 6007 1413 sw
rect 5990 1381 6007 1406
rect 6131 1381 6148 1413
rect 6330 1381 6345 1423
rect 6373 1381 6388 1423
rect 6570 1406 6580 1413
tri 6580 1406 6587 1413 sw
rect 6570 1381 6587 1406
rect 6711 1381 6728 1413
rect 6910 1381 6925 1423
rect 253 1343 285 1357
rect 833 1343 865 1357
rect 1413 1343 1445 1357
rect 1993 1343 2025 1357
rect 2573 1343 2605 1357
rect 3153 1343 3185 1357
rect 3733 1343 3765 1357
rect 4313 1343 4345 1357
rect 4893 1343 4925 1357
rect 5473 1343 5505 1357
rect 6053 1343 6085 1357
rect 6633 1343 6665 1357
rect 67 1257 82 1285
rect 148 1257 163 1285
rect 375 1257 390 1285
rect 457 1257 472 1286
rect 647 1257 662 1285
rect 728 1257 743 1285
rect 955 1257 970 1285
rect 1037 1257 1052 1286
rect 1227 1257 1242 1285
rect 1308 1257 1323 1285
rect 1535 1257 1550 1285
rect 1617 1257 1632 1286
rect 1807 1257 1822 1285
rect 1888 1257 1903 1285
rect 2115 1257 2130 1285
rect 2197 1257 2212 1286
rect 2387 1257 2402 1285
rect 2468 1257 2483 1285
rect 2695 1257 2710 1285
rect 2777 1257 2792 1286
rect 2967 1257 2982 1285
rect 3048 1257 3063 1285
rect 3275 1257 3290 1285
rect 3357 1257 3372 1286
rect 3547 1257 3562 1285
rect 3628 1257 3643 1285
rect 3855 1257 3870 1285
rect 3937 1257 3952 1286
rect 4127 1257 4142 1285
rect 4208 1257 4223 1285
rect 4435 1257 4450 1285
rect 4517 1257 4532 1286
rect 4707 1257 4722 1285
rect 4788 1257 4803 1285
rect 5015 1257 5030 1285
rect 5097 1257 5112 1286
rect 5287 1257 5302 1285
rect 5368 1257 5383 1285
rect 5595 1257 5610 1285
rect 5677 1257 5692 1286
rect 5867 1257 5882 1285
rect 5948 1257 5963 1285
rect 6175 1257 6190 1285
rect 6257 1257 6272 1286
rect 6447 1257 6462 1285
rect 6528 1257 6543 1285
rect 6755 1257 6770 1285
rect 6837 1257 6852 1286
rect -7 1111 8 1153
rect 190 1136 200 1143
tri 200 1136 207 1143 sw
rect 190 1111 207 1136
rect 331 1111 348 1143
rect 530 1111 545 1153
rect 573 1111 588 1153
rect 770 1136 780 1143
tri 780 1136 787 1143 sw
rect 770 1111 787 1136
rect 911 1111 928 1143
rect 1110 1111 1125 1153
rect 1153 1111 1168 1153
rect 1350 1136 1360 1143
tri 1360 1136 1367 1143 sw
rect 1350 1111 1367 1136
rect 1491 1111 1508 1143
rect 1690 1111 1705 1153
rect 1733 1111 1748 1153
rect 1930 1136 1940 1143
tri 1940 1136 1947 1143 sw
rect 1930 1111 1947 1136
rect 2071 1111 2088 1143
rect 2270 1111 2285 1153
rect 2313 1111 2328 1153
rect 2510 1136 2520 1143
tri 2520 1136 2527 1143 sw
rect 2510 1111 2527 1136
rect 2651 1111 2668 1143
rect 2850 1111 2865 1153
rect 2893 1111 2908 1153
rect 3090 1136 3100 1143
tri 3100 1136 3107 1143 sw
rect 3090 1111 3107 1136
rect 3231 1111 3248 1143
rect 3430 1111 3445 1153
rect 3473 1111 3488 1153
rect 3670 1136 3680 1143
tri 3680 1136 3687 1143 sw
rect 3670 1111 3687 1136
rect 3811 1111 3828 1143
rect 4010 1111 4025 1153
rect 4053 1111 4068 1153
rect 4250 1136 4260 1143
tri 4260 1136 4267 1143 sw
rect 4250 1111 4267 1136
rect 4391 1111 4408 1143
rect 4590 1111 4605 1153
rect 4633 1111 4648 1153
rect 4830 1136 4840 1143
tri 4840 1136 4847 1143 sw
rect 4830 1111 4847 1136
rect 4971 1111 4988 1143
rect 5170 1111 5185 1153
rect 5213 1111 5228 1153
rect 5410 1136 5420 1143
tri 5420 1136 5427 1143 sw
rect 5410 1111 5427 1136
rect 5551 1111 5568 1143
rect 5750 1111 5765 1153
rect 5793 1111 5808 1153
rect 5990 1136 6000 1143
tri 6000 1136 6007 1143 sw
rect 5990 1111 6007 1136
rect 6131 1111 6148 1143
rect 6330 1111 6345 1153
rect 6373 1111 6388 1153
rect 6570 1136 6580 1143
tri 6580 1136 6587 1143 sw
rect 6570 1111 6587 1136
rect 6711 1111 6728 1143
rect 6910 1111 6925 1153
rect 253 1073 285 1087
rect 833 1073 865 1087
rect 1413 1073 1445 1087
rect 1993 1073 2025 1087
rect 2573 1073 2605 1087
rect 3153 1073 3185 1087
rect 3733 1073 3765 1087
rect 4313 1073 4345 1087
rect 4893 1073 4925 1087
rect 5473 1073 5505 1087
rect 6053 1073 6085 1087
rect 6633 1073 6665 1087
rect 67 987 82 1015
rect 148 987 163 1015
rect 375 987 390 1015
rect 457 987 472 1016
rect 647 987 662 1015
rect 728 987 743 1015
rect 955 987 970 1015
rect 1037 987 1052 1016
rect 1227 987 1242 1015
rect 1308 987 1323 1015
rect 1535 987 1550 1015
rect 1617 987 1632 1016
rect 1807 987 1822 1015
rect 1888 987 1903 1015
rect 2115 987 2130 1015
rect 2197 987 2212 1016
rect 2387 987 2402 1015
rect 2468 987 2483 1015
rect 2695 987 2710 1015
rect 2777 987 2792 1016
rect 2967 987 2982 1015
rect 3048 987 3063 1015
rect 3275 987 3290 1015
rect 3357 987 3372 1016
rect 3547 987 3562 1015
rect 3628 987 3643 1015
rect 3855 987 3870 1015
rect 3937 987 3952 1016
rect 4127 987 4142 1015
rect 4208 987 4223 1015
rect 4435 987 4450 1015
rect 4517 987 4532 1016
rect 4707 987 4722 1015
rect 4788 987 4803 1015
rect 5015 987 5030 1015
rect 5097 987 5112 1016
rect 5287 987 5302 1015
rect 5368 987 5383 1015
rect 5595 987 5610 1015
rect 5677 987 5692 1016
rect 5867 987 5882 1015
rect 5948 987 5963 1015
rect 6175 987 6190 1015
rect 6257 987 6272 1016
rect 6447 987 6462 1015
rect 6528 987 6543 1015
rect 6755 987 6770 1015
rect 6837 987 6852 1016
rect -7 841 8 883
rect 190 866 200 873
tri 200 866 207 873 sw
rect 190 841 207 866
rect 331 841 348 873
rect 530 841 545 883
rect 573 841 588 883
rect 770 866 780 873
tri 780 866 787 873 sw
rect 770 841 787 866
rect 911 841 928 873
rect 1110 841 1125 883
rect 1153 841 1168 883
rect 1350 866 1360 873
tri 1360 866 1367 873 sw
rect 1350 841 1367 866
rect 1491 841 1508 873
rect 1690 841 1705 883
rect 1733 841 1748 883
rect 1930 866 1940 873
tri 1940 866 1947 873 sw
rect 1930 841 1947 866
rect 2071 841 2088 873
rect 2270 841 2285 883
rect 2313 841 2328 883
rect 2510 866 2520 873
tri 2520 866 2527 873 sw
rect 2510 841 2527 866
rect 2651 841 2668 873
rect 2850 841 2865 883
rect 2893 841 2908 883
rect 3090 866 3100 873
tri 3100 866 3107 873 sw
rect 3090 841 3107 866
rect 3231 841 3248 873
rect 3430 841 3445 883
rect 3473 841 3488 883
rect 3670 866 3680 873
tri 3680 866 3687 873 sw
rect 3670 841 3687 866
rect 3811 841 3828 873
rect 4010 841 4025 883
rect 4053 841 4068 883
rect 4250 866 4260 873
tri 4260 866 4267 873 sw
rect 4250 841 4267 866
rect 4391 841 4408 873
rect 4590 841 4605 883
rect 4633 841 4648 883
rect 4830 866 4840 873
tri 4840 866 4847 873 sw
rect 4830 841 4847 866
rect 4971 841 4988 873
rect 5170 841 5185 883
rect 5213 841 5228 883
rect 5410 866 5420 873
tri 5420 866 5427 873 sw
rect 5410 841 5427 866
rect 5551 841 5568 873
rect 5750 841 5765 883
rect 5793 841 5808 883
rect 5990 866 6000 873
tri 6000 866 6007 873 sw
rect 5990 841 6007 866
rect 6131 841 6148 873
rect 6330 841 6345 883
rect 6373 841 6388 883
rect 6570 866 6580 873
tri 6580 866 6587 873 sw
rect 6570 841 6587 866
rect 6711 841 6728 873
rect 6910 841 6925 883
rect 253 803 285 817
rect 833 803 865 817
rect 1413 803 1445 817
rect 1993 803 2025 817
rect 2573 803 2605 817
rect 3153 803 3185 817
rect 3733 803 3765 817
rect 4313 803 4345 817
rect 4893 803 4925 817
rect 5473 803 5505 817
rect 6053 803 6085 817
rect 6633 803 6665 817
rect 67 717 82 745
rect 148 717 163 745
rect 375 717 390 745
rect 457 717 472 746
rect 647 717 662 745
rect 728 717 743 745
rect 955 717 970 745
rect 1037 717 1052 746
rect 1227 717 1242 745
rect 1308 717 1323 745
rect 1535 717 1550 745
rect 1617 717 1632 746
rect 1807 717 1822 745
rect 1888 717 1903 745
rect 2115 717 2130 745
rect 2197 717 2212 746
rect 2387 717 2402 745
rect 2468 717 2483 745
rect 2695 717 2710 745
rect 2777 717 2792 746
rect 2967 717 2982 745
rect 3048 717 3063 745
rect 3275 717 3290 745
rect 3357 717 3372 746
rect 3547 717 3562 745
rect 3628 717 3643 745
rect 3855 717 3870 745
rect 3937 717 3952 746
rect 4127 717 4142 745
rect 4208 717 4223 745
rect 4435 717 4450 745
rect 4517 717 4532 746
rect 4707 717 4722 745
rect 4788 717 4803 745
rect 5015 717 5030 745
rect 5097 717 5112 746
rect 5287 717 5302 745
rect 5368 717 5383 745
rect 5595 717 5610 745
rect 5677 717 5692 746
rect 5867 717 5882 745
rect 5948 717 5963 745
rect 6175 717 6190 745
rect 6257 717 6272 746
rect 6447 717 6462 745
rect 6528 717 6543 745
rect 6755 717 6770 745
rect 6837 717 6852 746
rect -7 571 8 613
rect 190 596 200 603
tri 200 596 207 603 sw
rect 190 571 207 596
rect 331 571 348 603
rect 530 571 545 613
rect 573 571 588 613
rect 770 596 780 603
tri 780 596 787 603 sw
rect 770 571 787 596
rect 911 571 928 603
rect 1110 571 1125 613
rect 1153 571 1168 613
rect 1350 596 1360 603
tri 1360 596 1367 603 sw
rect 1350 571 1367 596
rect 1491 571 1508 603
rect 1690 571 1705 613
rect 1733 571 1748 613
rect 1930 596 1940 603
tri 1940 596 1947 603 sw
rect 1930 571 1947 596
rect 2071 571 2088 603
rect 2270 571 2285 613
rect 2313 571 2328 613
rect 2510 596 2520 603
tri 2520 596 2527 603 sw
rect 2510 571 2527 596
rect 2651 571 2668 603
rect 2850 571 2865 613
rect 2893 571 2908 613
rect 3090 596 3100 603
tri 3100 596 3107 603 sw
rect 3090 571 3107 596
rect 3231 571 3248 603
rect 3430 571 3445 613
rect 3473 571 3488 613
rect 3670 596 3680 603
tri 3680 596 3687 603 sw
rect 3670 571 3687 596
rect 3811 571 3828 603
rect 4010 571 4025 613
rect 4053 571 4068 613
rect 4250 596 4260 603
tri 4260 596 4267 603 sw
rect 4250 571 4267 596
rect 4391 571 4408 603
rect 4590 571 4605 613
rect 4633 571 4648 613
rect 4830 596 4840 603
tri 4840 596 4847 603 sw
rect 4830 571 4847 596
rect 4971 571 4988 603
rect 5170 571 5185 613
rect 5213 571 5228 613
rect 5410 596 5420 603
tri 5420 596 5427 603 sw
rect 5410 571 5427 596
rect 5551 571 5568 603
rect 5750 571 5765 613
rect 5793 571 5808 613
rect 5990 596 6000 603
tri 6000 596 6007 603 sw
rect 5990 571 6007 596
rect 6131 571 6148 603
rect 6330 571 6345 613
rect 6373 571 6388 613
rect 6570 596 6580 603
tri 6580 596 6587 603 sw
rect 6570 571 6587 596
rect 6711 571 6728 603
rect 6910 571 6925 613
rect 253 533 285 547
rect 833 533 865 547
rect 1413 533 1445 547
rect 1993 533 2025 547
rect 2573 533 2605 547
rect 3153 533 3185 547
rect 3733 533 3765 547
rect 4313 533 4345 547
rect 4893 533 4925 547
rect 5473 533 5505 547
rect 6053 533 6085 547
rect 6633 533 6665 547
rect 67 447 82 475
rect 148 447 163 475
rect 375 447 390 475
rect 457 447 472 476
rect 647 447 662 475
rect 728 447 743 475
rect 955 447 970 475
rect 1037 447 1052 476
rect 1227 447 1242 475
rect 1308 447 1323 475
rect 1535 447 1550 475
rect 1617 447 1632 476
rect 1807 447 1822 475
rect 1888 447 1903 475
rect 2115 447 2130 475
rect 2197 447 2212 476
rect 2387 447 2402 475
rect 2468 447 2483 475
rect 2695 447 2710 475
rect 2777 447 2792 476
rect 2967 447 2982 475
rect 3048 447 3063 475
rect 3275 447 3290 475
rect 3357 447 3372 476
rect 3547 447 3562 475
rect 3628 447 3643 475
rect 3855 447 3870 475
rect 3937 447 3952 476
rect 4127 447 4142 475
rect 4208 447 4223 475
rect 4435 447 4450 475
rect 4517 447 4532 476
rect 4707 447 4722 475
rect 4788 447 4803 475
rect 5015 447 5030 475
rect 5097 447 5112 476
rect 5287 447 5302 475
rect 5368 447 5383 475
rect 5595 447 5610 475
rect 5677 447 5692 476
rect 5867 447 5882 475
rect 5948 447 5963 475
rect 6175 447 6190 475
rect 6257 447 6272 476
rect 6447 447 6462 475
rect 6528 447 6543 475
rect 6755 447 6770 475
rect 6837 447 6852 476
rect -7 301 8 343
rect 190 326 200 333
tri 200 326 207 333 sw
rect 190 301 207 326
rect 331 301 348 333
rect 530 301 545 343
rect 573 301 588 343
rect 770 326 780 333
tri 780 326 787 333 sw
rect 770 301 787 326
rect 911 301 928 333
rect 1110 301 1125 343
rect 1153 301 1168 343
rect 1350 326 1360 333
tri 1360 326 1367 333 sw
rect 1350 301 1367 326
rect 1491 301 1508 333
rect 1690 301 1705 343
rect 1733 301 1748 343
rect 1930 326 1940 333
tri 1940 326 1947 333 sw
rect 1930 301 1947 326
rect 2071 301 2088 333
rect 2270 301 2285 343
rect 2313 301 2328 343
rect 2510 326 2520 333
tri 2520 326 2527 333 sw
rect 2510 301 2527 326
rect 2651 301 2668 333
rect 2850 301 2865 343
rect 2893 301 2908 343
rect 3090 326 3100 333
tri 3100 326 3107 333 sw
rect 3090 301 3107 326
rect 3231 301 3248 333
rect 3430 301 3445 343
rect 3473 301 3488 343
rect 3670 326 3680 333
tri 3680 326 3687 333 sw
rect 3670 301 3687 326
rect 3811 301 3828 333
rect 4010 301 4025 343
rect 4053 301 4068 343
rect 4250 326 4260 333
tri 4260 326 4267 333 sw
rect 4250 301 4267 326
rect 4391 301 4408 333
rect 4590 301 4605 343
rect 4633 301 4648 343
rect 4830 326 4840 333
tri 4840 326 4847 333 sw
rect 4830 301 4847 326
rect 4971 301 4988 333
rect 5170 301 5185 343
rect 5213 301 5228 343
rect 5410 326 5420 333
tri 5420 326 5427 333 sw
rect 5410 301 5427 326
rect 5551 301 5568 333
rect 5750 301 5765 343
rect 5793 301 5808 343
rect 5990 326 6000 333
tri 6000 326 6007 333 sw
rect 5990 301 6007 326
rect 6131 301 6148 333
rect 6330 301 6345 343
rect 6373 301 6388 343
rect 6570 326 6580 333
tri 6580 326 6587 333 sw
rect 6570 301 6587 326
rect 6711 301 6728 333
rect 6910 301 6925 343
rect 253 263 285 277
rect 833 263 865 277
rect 1413 263 1445 277
rect 1993 263 2025 277
rect 2573 263 2605 277
rect 3153 263 3185 277
rect 3733 263 3765 277
rect 4313 263 4345 277
rect 4893 263 4925 277
rect 5473 263 5505 277
rect 6053 263 6085 277
rect 6633 263 6665 277
rect 67 177 82 205
rect 148 177 163 205
rect 375 177 390 205
rect 457 177 472 206
rect 647 177 662 205
rect 728 177 743 205
rect 955 177 970 205
rect 1037 177 1052 206
rect 1227 177 1242 205
rect 1308 177 1323 205
rect 1535 177 1550 205
rect 1617 177 1632 206
rect 1807 177 1822 205
rect 1888 177 1903 205
rect 2115 177 2130 205
rect 2197 177 2212 206
rect 2387 177 2402 205
rect 2468 177 2483 205
rect 2695 177 2710 205
rect 2777 177 2792 206
rect 2967 177 2982 205
rect 3048 177 3063 205
rect 3275 177 3290 205
rect 3357 177 3372 206
rect 3547 177 3562 205
rect 3628 177 3643 205
rect 3855 177 3870 205
rect 3937 177 3952 206
rect 4127 177 4142 205
rect 4208 177 4223 205
rect 4435 177 4450 205
rect 4517 177 4532 206
rect 4707 177 4722 205
rect 4788 177 4803 205
rect 5015 177 5030 205
rect 5097 177 5112 206
rect 5287 177 5302 205
rect 5368 177 5383 205
rect 5595 177 5610 205
rect 5677 177 5692 206
rect 5867 177 5882 205
rect 5948 177 5963 205
rect 6175 177 6190 205
rect 6257 177 6272 206
rect 6447 177 6462 205
rect 6528 177 6543 205
rect 6755 177 6770 205
rect 6837 177 6852 206
rect -7 31 8 73
rect 190 56 200 63
tri 200 56 207 63 sw
rect 190 31 207 56
rect 331 31 348 63
rect 530 31 545 73
rect 573 31 588 73
rect 770 56 780 63
tri 780 56 787 63 sw
rect 770 31 787 56
rect 911 31 928 63
rect 1110 31 1125 73
rect 1153 31 1168 73
rect 1350 56 1360 63
tri 1360 56 1367 63 sw
rect 1350 31 1367 56
rect 1491 31 1508 63
rect 1690 31 1705 73
rect 1733 31 1748 73
rect 1930 56 1940 63
tri 1940 56 1947 63 sw
rect 1930 31 1947 56
rect 2071 31 2088 63
rect 2270 31 2285 73
rect 2313 31 2328 73
rect 2510 56 2520 63
tri 2520 56 2527 63 sw
rect 2510 31 2527 56
rect 2651 31 2668 63
rect 2850 31 2865 73
rect 2893 31 2908 73
rect 3090 56 3100 63
tri 3100 56 3107 63 sw
rect 3090 31 3107 56
rect 3231 31 3248 63
rect 3430 31 3445 73
rect 3473 31 3488 73
rect 3670 56 3680 63
tri 3680 56 3687 63 sw
rect 3670 31 3687 56
rect 3811 31 3828 63
rect 4010 31 4025 73
rect 4053 31 4068 73
rect 4250 56 4260 63
tri 4260 56 4267 63 sw
rect 4250 31 4267 56
rect 4391 31 4408 63
rect 4590 31 4605 73
rect 4633 31 4648 73
rect 4830 56 4840 63
tri 4840 56 4847 63 sw
rect 4830 31 4847 56
rect 4971 31 4988 63
rect 5170 31 5185 73
rect 5213 31 5228 73
rect 5410 56 5420 63
tri 5420 56 5427 63 sw
rect 5410 31 5427 56
rect 5551 31 5568 63
rect 5750 31 5765 73
rect 5793 31 5808 73
rect 5990 56 6000 63
tri 6000 56 6007 63 sw
rect 5990 31 6007 56
rect 6131 31 6148 63
rect 6330 31 6345 73
rect 6373 31 6388 73
rect 6570 56 6580 63
tri 6580 56 6587 63 sw
rect 6570 31 6587 56
rect 6711 31 6728 63
rect 6910 31 6925 73
rect 253 -7 285 7
rect 833 -7 865 7
rect 1413 -7 1445 7
rect 1993 -7 2025 7
rect 2573 -7 2605 7
rect 3153 -7 3185 7
rect 3733 -7 3765 7
rect 4313 -7 4345 7
rect 4893 -7 4925 7
rect 5473 -7 5505 7
rect 6053 -7 6085 7
rect 6633 -7 6665 7
<< pdiffc >>
rect 253 4269 285 4283
rect 191 4217 206 4245
rect 332 4229 344 4245
tri 332 4217 344 4229 ne
rect 833 4269 865 4283
rect 771 4217 786 4245
rect 912 4229 924 4245
tri 912 4217 924 4229 ne
rect 1413 4269 1445 4283
rect 1351 4217 1366 4245
rect 1492 4229 1504 4245
tri 1492 4217 1504 4229 ne
rect 1993 4269 2025 4283
rect 1931 4217 1946 4245
rect 2072 4229 2084 4245
tri 2072 4217 2084 4229 ne
rect 2573 4269 2605 4283
rect 2511 4217 2526 4245
rect 2652 4229 2664 4245
tri 2652 4217 2664 4229 ne
rect 3153 4269 3185 4283
rect 3091 4217 3106 4245
rect 3232 4229 3244 4245
tri 3232 4217 3244 4229 ne
rect 3733 4269 3765 4283
rect 3671 4217 3686 4245
rect 3812 4229 3824 4245
tri 3812 4217 3824 4229 ne
rect 4313 4269 4345 4283
rect 4251 4217 4266 4245
rect 4392 4229 4404 4245
tri 4392 4217 4404 4229 ne
rect 4893 4269 4925 4283
rect 4831 4217 4846 4245
rect 4972 4229 4984 4245
tri 4972 4217 4984 4229 ne
rect 5473 4269 5505 4283
rect 5411 4217 5426 4245
rect 5552 4229 5564 4245
tri 5552 4217 5564 4229 ne
rect 6053 4269 6085 4283
rect 5991 4217 6006 4245
rect 6132 4229 6144 4245
tri 6132 4217 6144 4229 ne
rect 6633 4269 6665 4283
rect 6571 4217 6586 4245
rect 6712 4229 6724 4245
tri 6712 4217 6724 4229 ne
rect 253 3999 285 4013
rect 191 3947 206 3975
rect 332 3959 344 3975
tri 332 3947 344 3959 ne
rect 833 3999 865 4013
rect 771 3947 786 3975
rect 912 3959 924 3975
tri 912 3947 924 3959 ne
rect 1413 3999 1445 4013
rect 1351 3947 1366 3975
rect 1492 3959 1504 3975
tri 1492 3947 1504 3959 ne
rect 1993 3999 2025 4013
rect 1931 3947 1946 3975
rect 2072 3959 2084 3975
tri 2072 3947 2084 3959 ne
rect 2573 3999 2605 4013
rect 2511 3947 2526 3975
rect 2652 3959 2664 3975
tri 2652 3947 2664 3959 ne
rect 3153 3999 3185 4013
rect 3091 3947 3106 3975
rect 3232 3959 3244 3975
tri 3232 3947 3244 3959 ne
rect 3733 3999 3765 4013
rect 3671 3947 3686 3975
rect 3812 3959 3824 3975
tri 3812 3947 3824 3959 ne
rect 4313 3999 4345 4013
rect 4251 3947 4266 3975
rect 4392 3959 4404 3975
tri 4392 3947 4404 3959 ne
rect 4893 3999 4925 4013
rect 4831 3947 4846 3975
rect 4972 3959 4984 3975
tri 4972 3947 4984 3959 ne
rect 5473 3999 5505 4013
rect 5411 3947 5426 3975
rect 5552 3959 5564 3975
tri 5552 3947 5564 3959 ne
rect 6053 3999 6085 4013
rect 5991 3947 6006 3975
rect 6132 3959 6144 3975
tri 6132 3947 6144 3959 ne
rect 6633 3999 6665 4013
rect 6571 3947 6586 3975
rect 6712 3959 6724 3975
tri 6712 3947 6724 3959 ne
rect 253 3729 285 3743
rect 191 3677 206 3705
rect 332 3689 344 3705
tri 332 3677 344 3689 ne
rect 833 3729 865 3743
rect 771 3677 786 3705
rect 912 3689 924 3705
tri 912 3677 924 3689 ne
rect 1413 3729 1445 3743
rect 1351 3677 1366 3705
rect 1492 3689 1504 3705
tri 1492 3677 1504 3689 ne
rect 1993 3729 2025 3743
rect 1931 3677 1946 3705
rect 2072 3689 2084 3705
tri 2072 3677 2084 3689 ne
rect 2573 3729 2605 3743
rect 2511 3677 2526 3705
rect 2652 3689 2664 3705
tri 2652 3677 2664 3689 ne
rect 3153 3729 3185 3743
rect 3091 3677 3106 3705
rect 3232 3689 3244 3705
tri 3232 3677 3244 3689 ne
rect 3733 3729 3765 3743
rect 3671 3677 3686 3705
rect 3812 3689 3824 3705
tri 3812 3677 3824 3689 ne
rect 4313 3729 4345 3743
rect 4251 3677 4266 3705
rect 4392 3689 4404 3705
tri 4392 3677 4404 3689 ne
rect 4893 3729 4925 3743
rect 4831 3677 4846 3705
rect 4972 3689 4984 3705
tri 4972 3677 4984 3689 ne
rect 5473 3729 5505 3743
rect 5411 3677 5426 3705
rect 5552 3689 5564 3705
tri 5552 3677 5564 3689 ne
rect 6053 3729 6085 3743
rect 5991 3677 6006 3705
rect 6132 3689 6144 3705
tri 6132 3677 6144 3689 ne
rect 6633 3729 6665 3743
rect 6571 3677 6586 3705
rect 6712 3689 6724 3705
tri 6712 3677 6724 3689 ne
rect 253 3459 285 3473
rect 191 3407 206 3435
rect 332 3419 344 3435
tri 332 3407 344 3419 ne
rect 833 3459 865 3473
rect 771 3407 786 3435
rect 912 3419 924 3435
tri 912 3407 924 3419 ne
rect 1413 3459 1445 3473
rect 1351 3407 1366 3435
rect 1492 3419 1504 3435
tri 1492 3407 1504 3419 ne
rect 1993 3459 2025 3473
rect 1931 3407 1946 3435
rect 2072 3419 2084 3435
tri 2072 3407 2084 3419 ne
rect 2573 3459 2605 3473
rect 2511 3407 2526 3435
rect 2652 3419 2664 3435
tri 2652 3407 2664 3419 ne
rect 3153 3459 3185 3473
rect 3091 3407 3106 3435
rect 3232 3419 3244 3435
tri 3232 3407 3244 3419 ne
rect 3733 3459 3765 3473
rect 3671 3407 3686 3435
rect 3812 3419 3824 3435
tri 3812 3407 3824 3419 ne
rect 4313 3459 4345 3473
rect 4251 3407 4266 3435
rect 4392 3419 4404 3435
tri 4392 3407 4404 3419 ne
rect 4893 3459 4925 3473
rect 4831 3407 4846 3435
rect 4972 3419 4984 3435
tri 4972 3407 4984 3419 ne
rect 5473 3459 5505 3473
rect 5411 3407 5426 3435
rect 5552 3419 5564 3435
tri 5552 3407 5564 3419 ne
rect 6053 3459 6085 3473
rect 5991 3407 6006 3435
rect 6132 3419 6144 3435
tri 6132 3407 6144 3419 ne
rect 6633 3459 6665 3473
rect 6571 3407 6586 3435
rect 6712 3419 6724 3435
tri 6712 3407 6724 3419 ne
rect 253 3189 285 3203
rect 191 3137 206 3165
rect 332 3149 344 3165
tri 332 3137 344 3149 ne
rect 833 3189 865 3203
rect 771 3137 786 3165
rect 912 3149 924 3165
tri 912 3137 924 3149 ne
rect 1413 3189 1445 3203
rect 1351 3137 1366 3165
rect 1492 3149 1504 3165
tri 1492 3137 1504 3149 ne
rect 1993 3189 2025 3203
rect 1931 3137 1946 3165
rect 2072 3149 2084 3165
tri 2072 3137 2084 3149 ne
rect 2573 3189 2605 3203
rect 2511 3137 2526 3165
rect 2652 3149 2664 3165
tri 2652 3137 2664 3149 ne
rect 3153 3189 3185 3203
rect 3091 3137 3106 3165
rect 3232 3149 3244 3165
tri 3232 3137 3244 3149 ne
rect 3733 3189 3765 3203
rect 3671 3137 3686 3165
rect 3812 3149 3824 3165
tri 3812 3137 3824 3149 ne
rect 4313 3189 4345 3203
rect 4251 3137 4266 3165
rect 4392 3149 4404 3165
tri 4392 3137 4404 3149 ne
rect 4893 3189 4925 3203
rect 4831 3137 4846 3165
rect 4972 3149 4984 3165
tri 4972 3137 4984 3149 ne
rect 5473 3189 5505 3203
rect 5411 3137 5426 3165
rect 5552 3149 5564 3165
tri 5552 3137 5564 3149 ne
rect 6053 3189 6085 3203
rect 5991 3137 6006 3165
rect 6132 3149 6144 3165
tri 6132 3137 6144 3149 ne
rect 6633 3189 6665 3203
rect 6571 3137 6586 3165
rect 6712 3149 6724 3165
tri 6712 3137 6724 3149 ne
rect 253 2919 285 2933
rect 191 2867 206 2895
rect 332 2879 344 2895
tri 332 2867 344 2879 ne
rect 833 2919 865 2933
rect 771 2867 786 2895
rect 912 2879 924 2895
tri 912 2867 924 2879 ne
rect 1413 2919 1445 2933
rect 1351 2867 1366 2895
rect 1492 2879 1504 2895
tri 1492 2867 1504 2879 ne
rect 1993 2919 2025 2933
rect 1931 2867 1946 2895
rect 2072 2879 2084 2895
tri 2072 2867 2084 2879 ne
rect 2573 2919 2605 2933
rect 2511 2867 2526 2895
rect 2652 2879 2664 2895
tri 2652 2867 2664 2879 ne
rect 3153 2919 3185 2933
rect 3091 2867 3106 2895
rect 3232 2879 3244 2895
tri 3232 2867 3244 2879 ne
rect 3733 2919 3765 2933
rect 3671 2867 3686 2895
rect 3812 2879 3824 2895
tri 3812 2867 3824 2879 ne
rect 4313 2919 4345 2933
rect 4251 2867 4266 2895
rect 4392 2879 4404 2895
tri 4392 2867 4404 2879 ne
rect 4893 2919 4925 2933
rect 4831 2867 4846 2895
rect 4972 2879 4984 2895
tri 4972 2867 4984 2879 ne
rect 5473 2919 5505 2933
rect 5411 2867 5426 2895
rect 5552 2879 5564 2895
tri 5552 2867 5564 2879 ne
rect 6053 2919 6085 2933
rect 5991 2867 6006 2895
rect 6132 2879 6144 2895
tri 6132 2867 6144 2879 ne
rect 6633 2919 6665 2933
rect 6571 2867 6586 2895
rect 6712 2879 6724 2895
tri 6712 2867 6724 2879 ne
rect 253 2649 285 2663
rect 191 2597 206 2625
rect 332 2609 344 2625
tri 332 2597 344 2609 ne
rect 833 2649 865 2663
rect 771 2597 786 2625
rect 912 2609 924 2625
tri 912 2597 924 2609 ne
rect 1413 2649 1445 2663
rect 1351 2597 1366 2625
rect 1492 2609 1504 2625
tri 1492 2597 1504 2609 ne
rect 1993 2649 2025 2663
rect 1931 2597 1946 2625
rect 2072 2609 2084 2625
tri 2072 2597 2084 2609 ne
rect 2573 2649 2605 2663
rect 2511 2597 2526 2625
rect 2652 2609 2664 2625
tri 2652 2597 2664 2609 ne
rect 3153 2649 3185 2663
rect 3091 2597 3106 2625
rect 3232 2609 3244 2625
tri 3232 2597 3244 2609 ne
rect 3733 2649 3765 2663
rect 3671 2597 3686 2625
rect 3812 2609 3824 2625
tri 3812 2597 3824 2609 ne
rect 4313 2649 4345 2663
rect 4251 2597 4266 2625
rect 4392 2609 4404 2625
tri 4392 2597 4404 2609 ne
rect 4893 2649 4925 2663
rect 4831 2597 4846 2625
rect 4972 2609 4984 2625
tri 4972 2597 4984 2609 ne
rect 5473 2649 5505 2663
rect 5411 2597 5426 2625
rect 5552 2609 5564 2625
tri 5552 2597 5564 2609 ne
rect 6053 2649 6085 2663
rect 5991 2597 6006 2625
rect 6132 2609 6144 2625
tri 6132 2597 6144 2609 ne
rect 6633 2649 6665 2663
rect 6571 2597 6586 2625
rect 6712 2609 6724 2625
tri 6712 2597 6724 2609 ne
rect 253 2379 285 2393
rect 191 2327 206 2355
rect 332 2339 344 2355
tri 332 2327 344 2339 ne
rect 833 2379 865 2393
rect 771 2327 786 2355
rect 912 2339 924 2355
tri 912 2327 924 2339 ne
rect 1413 2379 1445 2393
rect 1351 2327 1366 2355
rect 1492 2339 1504 2355
tri 1492 2327 1504 2339 ne
rect 1993 2379 2025 2393
rect 1931 2327 1946 2355
rect 2072 2339 2084 2355
tri 2072 2327 2084 2339 ne
rect 2573 2379 2605 2393
rect 2511 2327 2526 2355
rect 2652 2339 2664 2355
tri 2652 2327 2664 2339 ne
rect 3153 2379 3185 2393
rect 3091 2327 3106 2355
rect 3232 2339 3244 2355
tri 3232 2327 3244 2339 ne
rect 3733 2379 3765 2393
rect 3671 2327 3686 2355
rect 3812 2339 3824 2355
tri 3812 2327 3824 2339 ne
rect 4313 2379 4345 2393
rect 4251 2327 4266 2355
rect 4392 2339 4404 2355
tri 4392 2327 4404 2339 ne
rect 4893 2379 4925 2393
rect 4831 2327 4846 2355
rect 4972 2339 4984 2355
tri 4972 2327 4984 2339 ne
rect 5473 2379 5505 2393
rect 5411 2327 5426 2355
rect 5552 2339 5564 2355
tri 5552 2327 5564 2339 ne
rect 6053 2379 6085 2393
rect 5991 2327 6006 2355
rect 6132 2339 6144 2355
tri 6132 2327 6144 2339 ne
rect 6633 2379 6665 2393
rect 6571 2327 6586 2355
rect 6712 2339 6724 2355
tri 6712 2327 6724 2339 ne
rect 253 2109 285 2123
rect 191 2057 206 2085
rect 332 2069 344 2085
tri 332 2057 344 2069 ne
rect 833 2109 865 2123
rect 771 2057 786 2085
rect 912 2069 924 2085
tri 912 2057 924 2069 ne
rect 1413 2109 1445 2123
rect 1351 2057 1366 2085
rect 1492 2069 1504 2085
tri 1492 2057 1504 2069 ne
rect 1993 2109 2025 2123
rect 1931 2057 1946 2085
rect 2072 2069 2084 2085
tri 2072 2057 2084 2069 ne
rect 2573 2109 2605 2123
rect 2511 2057 2526 2085
rect 2652 2069 2664 2085
tri 2652 2057 2664 2069 ne
rect 3153 2109 3185 2123
rect 3091 2057 3106 2085
rect 3232 2069 3244 2085
tri 3232 2057 3244 2069 ne
rect 3733 2109 3765 2123
rect 3671 2057 3686 2085
rect 3812 2069 3824 2085
tri 3812 2057 3824 2069 ne
rect 4313 2109 4345 2123
rect 4251 2057 4266 2085
rect 4392 2069 4404 2085
tri 4392 2057 4404 2069 ne
rect 4893 2109 4925 2123
rect 4831 2057 4846 2085
rect 4972 2069 4984 2085
tri 4972 2057 4984 2069 ne
rect 5473 2109 5505 2123
rect 5411 2057 5426 2085
rect 5552 2069 5564 2085
tri 5552 2057 5564 2069 ne
rect 6053 2109 6085 2123
rect 5991 2057 6006 2085
rect 6132 2069 6144 2085
tri 6132 2057 6144 2069 ne
rect 6633 2109 6665 2123
rect 6571 2057 6586 2085
rect 6712 2069 6724 2085
tri 6712 2057 6724 2069 ne
rect 253 1839 285 1853
rect 191 1787 206 1815
rect 332 1799 344 1815
tri 332 1787 344 1799 ne
rect 833 1839 865 1853
rect 771 1787 786 1815
rect 912 1799 924 1815
tri 912 1787 924 1799 ne
rect 1413 1839 1445 1853
rect 1351 1787 1366 1815
rect 1492 1799 1504 1815
tri 1492 1787 1504 1799 ne
rect 1993 1839 2025 1853
rect 1931 1787 1946 1815
rect 2072 1799 2084 1815
tri 2072 1787 2084 1799 ne
rect 2573 1839 2605 1853
rect 2511 1787 2526 1815
rect 2652 1799 2664 1815
tri 2652 1787 2664 1799 ne
rect 3153 1839 3185 1853
rect 3091 1787 3106 1815
rect 3232 1799 3244 1815
tri 3232 1787 3244 1799 ne
rect 3733 1839 3765 1853
rect 3671 1787 3686 1815
rect 3812 1799 3824 1815
tri 3812 1787 3824 1799 ne
rect 4313 1839 4345 1853
rect 4251 1787 4266 1815
rect 4392 1799 4404 1815
tri 4392 1787 4404 1799 ne
rect 4893 1839 4925 1853
rect 4831 1787 4846 1815
rect 4972 1799 4984 1815
tri 4972 1787 4984 1799 ne
rect 5473 1839 5505 1853
rect 5411 1787 5426 1815
rect 5552 1799 5564 1815
tri 5552 1787 5564 1799 ne
rect 6053 1839 6085 1853
rect 5991 1787 6006 1815
rect 6132 1799 6144 1815
tri 6132 1787 6144 1799 ne
rect 6633 1839 6665 1853
rect 6571 1787 6586 1815
rect 6712 1799 6724 1815
tri 6712 1787 6724 1799 ne
rect 253 1569 285 1583
rect 191 1517 206 1545
rect 332 1529 344 1545
tri 332 1517 344 1529 ne
rect 833 1569 865 1583
rect 771 1517 786 1545
rect 912 1529 924 1545
tri 912 1517 924 1529 ne
rect 1413 1569 1445 1583
rect 1351 1517 1366 1545
rect 1492 1529 1504 1545
tri 1492 1517 1504 1529 ne
rect 1993 1569 2025 1583
rect 1931 1517 1946 1545
rect 2072 1529 2084 1545
tri 2072 1517 2084 1529 ne
rect 2573 1569 2605 1583
rect 2511 1517 2526 1545
rect 2652 1529 2664 1545
tri 2652 1517 2664 1529 ne
rect 3153 1569 3185 1583
rect 3091 1517 3106 1545
rect 3232 1529 3244 1545
tri 3232 1517 3244 1529 ne
rect 3733 1569 3765 1583
rect 3671 1517 3686 1545
rect 3812 1529 3824 1545
tri 3812 1517 3824 1529 ne
rect 4313 1569 4345 1583
rect 4251 1517 4266 1545
rect 4392 1529 4404 1545
tri 4392 1517 4404 1529 ne
rect 4893 1569 4925 1583
rect 4831 1517 4846 1545
rect 4972 1529 4984 1545
tri 4972 1517 4984 1529 ne
rect 5473 1569 5505 1583
rect 5411 1517 5426 1545
rect 5552 1529 5564 1545
tri 5552 1517 5564 1529 ne
rect 6053 1569 6085 1583
rect 5991 1517 6006 1545
rect 6132 1529 6144 1545
tri 6132 1517 6144 1529 ne
rect 6633 1569 6665 1583
rect 6571 1517 6586 1545
rect 6712 1529 6724 1545
tri 6712 1517 6724 1529 ne
rect 253 1299 285 1313
rect 191 1247 206 1275
rect 332 1259 344 1275
tri 332 1247 344 1259 ne
rect 833 1299 865 1313
rect 771 1247 786 1275
rect 912 1259 924 1275
tri 912 1247 924 1259 ne
rect 1413 1299 1445 1313
rect 1351 1247 1366 1275
rect 1492 1259 1504 1275
tri 1492 1247 1504 1259 ne
rect 1993 1299 2025 1313
rect 1931 1247 1946 1275
rect 2072 1259 2084 1275
tri 2072 1247 2084 1259 ne
rect 2573 1299 2605 1313
rect 2511 1247 2526 1275
rect 2652 1259 2664 1275
tri 2652 1247 2664 1259 ne
rect 3153 1299 3185 1313
rect 3091 1247 3106 1275
rect 3232 1259 3244 1275
tri 3232 1247 3244 1259 ne
rect 3733 1299 3765 1313
rect 3671 1247 3686 1275
rect 3812 1259 3824 1275
tri 3812 1247 3824 1259 ne
rect 4313 1299 4345 1313
rect 4251 1247 4266 1275
rect 4392 1259 4404 1275
tri 4392 1247 4404 1259 ne
rect 4893 1299 4925 1313
rect 4831 1247 4846 1275
rect 4972 1259 4984 1275
tri 4972 1247 4984 1259 ne
rect 5473 1299 5505 1313
rect 5411 1247 5426 1275
rect 5552 1259 5564 1275
tri 5552 1247 5564 1259 ne
rect 6053 1299 6085 1313
rect 5991 1247 6006 1275
rect 6132 1259 6144 1275
tri 6132 1247 6144 1259 ne
rect 6633 1299 6665 1313
rect 6571 1247 6586 1275
rect 6712 1259 6724 1275
tri 6712 1247 6724 1259 ne
rect 253 1029 285 1043
rect 191 977 206 1005
rect 332 989 344 1005
tri 332 977 344 989 ne
rect 833 1029 865 1043
rect 771 977 786 1005
rect 912 989 924 1005
tri 912 977 924 989 ne
rect 1413 1029 1445 1043
rect 1351 977 1366 1005
rect 1492 989 1504 1005
tri 1492 977 1504 989 ne
rect 1993 1029 2025 1043
rect 1931 977 1946 1005
rect 2072 989 2084 1005
tri 2072 977 2084 989 ne
rect 2573 1029 2605 1043
rect 2511 977 2526 1005
rect 2652 989 2664 1005
tri 2652 977 2664 989 ne
rect 3153 1029 3185 1043
rect 3091 977 3106 1005
rect 3232 989 3244 1005
tri 3232 977 3244 989 ne
rect 3733 1029 3765 1043
rect 3671 977 3686 1005
rect 3812 989 3824 1005
tri 3812 977 3824 989 ne
rect 4313 1029 4345 1043
rect 4251 977 4266 1005
rect 4392 989 4404 1005
tri 4392 977 4404 989 ne
rect 4893 1029 4925 1043
rect 4831 977 4846 1005
rect 4972 989 4984 1005
tri 4972 977 4984 989 ne
rect 5473 1029 5505 1043
rect 5411 977 5426 1005
rect 5552 989 5564 1005
tri 5552 977 5564 989 ne
rect 6053 1029 6085 1043
rect 5991 977 6006 1005
rect 6132 989 6144 1005
tri 6132 977 6144 989 ne
rect 6633 1029 6665 1043
rect 6571 977 6586 1005
rect 6712 989 6724 1005
tri 6712 977 6724 989 ne
rect 253 759 285 773
rect 191 707 206 735
rect 332 719 344 735
tri 332 707 344 719 ne
rect 833 759 865 773
rect 771 707 786 735
rect 912 719 924 735
tri 912 707 924 719 ne
rect 1413 759 1445 773
rect 1351 707 1366 735
rect 1492 719 1504 735
tri 1492 707 1504 719 ne
rect 1993 759 2025 773
rect 1931 707 1946 735
rect 2072 719 2084 735
tri 2072 707 2084 719 ne
rect 2573 759 2605 773
rect 2511 707 2526 735
rect 2652 719 2664 735
tri 2652 707 2664 719 ne
rect 3153 759 3185 773
rect 3091 707 3106 735
rect 3232 719 3244 735
tri 3232 707 3244 719 ne
rect 3733 759 3765 773
rect 3671 707 3686 735
rect 3812 719 3824 735
tri 3812 707 3824 719 ne
rect 4313 759 4345 773
rect 4251 707 4266 735
rect 4392 719 4404 735
tri 4392 707 4404 719 ne
rect 4893 759 4925 773
rect 4831 707 4846 735
rect 4972 719 4984 735
tri 4972 707 4984 719 ne
rect 5473 759 5505 773
rect 5411 707 5426 735
rect 5552 719 5564 735
tri 5552 707 5564 719 ne
rect 6053 759 6085 773
rect 5991 707 6006 735
rect 6132 719 6144 735
tri 6132 707 6144 719 ne
rect 6633 759 6665 773
rect 6571 707 6586 735
rect 6712 719 6724 735
tri 6712 707 6724 719 ne
rect 253 489 285 503
rect 191 437 206 465
rect 332 449 344 465
tri 332 437 344 449 ne
rect 833 489 865 503
rect 771 437 786 465
rect 912 449 924 465
tri 912 437 924 449 ne
rect 1413 489 1445 503
rect 1351 437 1366 465
rect 1492 449 1504 465
tri 1492 437 1504 449 ne
rect 1993 489 2025 503
rect 1931 437 1946 465
rect 2072 449 2084 465
tri 2072 437 2084 449 ne
rect 2573 489 2605 503
rect 2511 437 2526 465
rect 2652 449 2664 465
tri 2652 437 2664 449 ne
rect 3153 489 3185 503
rect 3091 437 3106 465
rect 3232 449 3244 465
tri 3232 437 3244 449 ne
rect 3733 489 3765 503
rect 3671 437 3686 465
rect 3812 449 3824 465
tri 3812 437 3824 449 ne
rect 4313 489 4345 503
rect 4251 437 4266 465
rect 4392 449 4404 465
tri 4392 437 4404 449 ne
rect 4893 489 4925 503
rect 4831 437 4846 465
rect 4972 449 4984 465
tri 4972 437 4984 449 ne
rect 5473 489 5505 503
rect 5411 437 5426 465
rect 5552 449 5564 465
tri 5552 437 5564 449 ne
rect 6053 489 6085 503
rect 5991 437 6006 465
rect 6132 449 6144 465
tri 6132 437 6144 449 ne
rect 6633 489 6665 503
rect 6571 437 6586 465
rect 6712 449 6724 465
tri 6712 437 6724 449 ne
rect 253 219 285 233
rect 191 167 206 195
rect 332 179 344 195
tri 332 167 344 179 ne
rect 833 219 865 233
rect 771 167 786 195
rect 912 179 924 195
tri 912 167 924 179 ne
rect 1413 219 1445 233
rect 1351 167 1366 195
rect 1492 179 1504 195
tri 1492 167 1504 179 ne
rect 1993 219 2025 233
rect 1931 167 1946 195
rect 2072 179 2084 195
tri 2072 167 2084 179 ne
rect 2573 219 2605 233
rect 2511 167 2526 195
rect 2652 179 2664 195
tri 2652 167 2664 179 ne
rect 3153 219 3185 233
rect 3091 167 3106 195
rect 3232 179 3244 195
tri 3232 167 3244 179 ne
rect 3733 219 3765 233
rect 3671 167 3686 195
rect 3812 179 3824 195
tri 3812 167 3824 179 ne
rect 4313 219 4345 233
rect 4251 167 4266 195
rect 4392 179 4404 195
tri 4392 167 4404 179 ne
rect 4893 219 4925 233
rect 4831 167 4846 195
rect 4972 179 4984 195
tri 4972 167 4984 179 ne
rect 5473 219 5505 233
rect 5411 167 5426 195
rect 5552 179 5564 195
tri 5552 167 5564 179 ne
rect 6053 219 6085 233
rect 5991 167 6006 195
rect 6132 179 6144 195
tri 6132 167 6144 179 ne
rect 6633 219 6665 233
rect 6571 167 6586 195
rect 6712 179 6724 195
tri 6712 167 6724 179 ne
<< psubdiffcont >>
rect 255 4057 283 4059
rect 835 4057 863 4059
rect 1415 4057 1443 4059
rect 1995 4057 2023 4059
rect 2575 4057 2603 4059
rect 3155 4057 3183 4059
rect 3735 4057 3763 4059
rect 4315 4057 4343 4059
rect 4895 4057 4923 4059
rect 5475 4057 5503 4059
rect 6055 4057 6083 4059
rect 6635 4057 6663 4059
rect 255 3787 283 3789
rect 835 3787 863 3789
rect 1415 3787 1443 3789
rect 1995 3787 2023 3789
rect 2575 3787 2603 3789
rect 3155 3787 3183 3789
rect 3735 3787 3763 3789
rect 4315 3787 4343 3789
rect 4895 3787 4923 3789
rect 5475 3787 5503 3789
rect 6055 3787 6083 3789
rect 6635 3787 6663 3789
rect 255 3517 283 3519
rect 835 3517 863 3519
rect 1415 3517 1443 3519
rect 1995 3517 2023 3519
rect 2575 3517 2603 3519
rect 3155 3517 3183 3519
rect 3735 3517 3763 3519
rect 4315 3517 4343 3519
rect 4895 3517 4923 3519
rect 5475 3517 5503 3519
rect 6055 3517 6083 3519
rect 6635 3517 6663 3519
rect 255 3247 283 3249
rect 835 3247 863 3249
rect 1415 3247 1443 3249
rect 1995 3247 2023 3249
rect 2575 3247 2603 3249
rect 3155 3247 3183 3249
rect 3735 3247 3763 3249
rect 4315 3247 4343 3249
rect 4895 3247 4923 3249
rect 5475 3247 5503 3249
rect 6055 3247 6083 3249
rect 6635 3247 6663 3249
rect 255 2977 283 2979
rect 835 2977 863 2979
rect 1415 2977 1443 2979
rect 1995 2977 2023 2979
rect 2575 2977 2603 2979
rect 3155 2977 3183 2979
rect 3735 2977 3763 2979
rect 4315 2977 4343 2979
rect 4895 2977 4923 2979
rect 5475 2977 5503 2979
rect 6055 2977 6083 2979
rect 6635 2977 6663 2979
rect 255 2707 283 2709
rect 835 2707 863 2709
rect 1415 2707 1443 2709
rect 1995 2707 2023 2709
rect 2575 2707 2603 2709
rect 3155 2707 3183 2709
rect 3735 2707 3763 2709
rect 4315 2707 4343 2709
rect 4895 2707 4923 2709
rect 5475 2707 5503 2709
rect 6055 2707 6083 2709
rect 6635 2707 6663 2709
rect 255 2437 283 2439
rect 835 2437 863 2439
rect 1415 2437 1443 2439
rect 1995 2437 2023 2439
rect 2575 2437 2603 2439
rect 3155 2437 3183 2439
rect 3735 2437 3763 2439
rect 4315 2437 4343 2439
rect 4895 2437 4923 2439
rect 5475 2437 5503 2439
rect 6055 2437 6083 2439
rect 6635 2437 6663 2439
rect 255 2167 283 2169
rect 835 2167 863 2169
rect 1415 2167 1443 2169
rect 1995 2167 2023 2169
rect 2575 2167 2603 2169
rect 3155 2167 3183 2169
rect 3735 2167 3763 2169
rect 4315 2167 4343 2169
rect 4895 2167 4923 2169
rect 5475 2167 5503 2169
rect 6055 2167 6083 2169
rect 6635 2167 6663 2169
rect 255 1897 283 1899
rect 835 1897 863 1899
rect 1415 1897 1443 1899
rect 1995 1897 2023 1899
rect 2575 1897 2603 1899
rect 3155 1897 3183 1899
rect 3735 1897 3763 1899
rect 4315 1897 4343 1899
rect 4895 1897 4923 1899
rect 5475 1897 5503 1899
rect 6055 1897 6083 1899
rect 6635 1897 6663 1899
rect 255 1627 283 1629
rect 835 1627 863 1629
rect 1415 1627 1443 1629
rect 1995 1627 2023 1629
rect 2575 1627 2603 1629
rect 3155 1627 3183 1629
rect 3735 1627 3763 1629
rect 4315 1627 4343 1629
rect 4895 1627 4923 1629
rect 5475 1627 5503 1629
rect 6055 1627 6083 1629
rect 6635 1627 6663 1629
rect 255 1357 283 1359
rect 835 1357 863 1359
rect 1415 1357 1443 1359
rect 1995 1357 2023 1359
rect 2575 1357 2603 1359
rect 3155 1357 3183 1359
rect 3735 1357 3763 1359
rect 4315 1357 4343 1359
rect 4895 1357 4923 1359
rect 5475 1357 5503 1359
rect 6055 1357 6083 1359
rect 6635 1357 6663 1359
rect 255 1087 283 1089
rect 835 1087 863 1089
rect 1415 1087 1443 1089
rect 1995 1087 2023 1089
rect 2575 1087 2603 1089
rect 3155 1087 3183 1089
rect 3735 1087 3763 1089
rect 4315 1087 4343 1089
rect 4895 1087 4923 1089
rect 5475 1087 5503 1089
rect 6055 1087 6083 1089
rect 6635 1087 6663 1089
rect 255 817 283 819
rect 835 817 863 819
rect 1415 817 1443 819
rect 1995 817 2023 819
rect 2575 817 2603 819
rect 3155 817 3183 819
rect 3735 817 3763 819
rect 4315 817 4343 819
rect 4895 817 4923 819
rect 5475 817 5503 819
rect 6055 817 6083 819
rect 6635 817 6663 819
rect 255 547 283 549
rect 835 547 863 549
rect 1415 547 1443 549
rect 1995 547 2023 549
rect 2575 547 2603 549
rect 3155 547 3183 549
rect 3735 547 3763 549
rect 4315 547 4343 549
rect 4895 547 4923 549
rect 5475 547 5503 549
rect 6055 547 6083 549
rect 6635 547 6663 549
rect 255 277 283 279
rect 835 277 863 279
rect 1415 277 1443 279
rect 1995 277 2023 279
rect 2575 277 2603 279
rect 3155 277 3183 279
rect 3735 277 3763 279
rect 4315 277 4343 279
rect 4895 277 4923 279
rect 5475 277 5503 279
rect 6055 277 6083 279
rect 6635 277 6663 279
rect 255 7 283 9
rect 835 7 863 9
rect 1415 7 1443 9
rect 1995 7 2023 9
rect 2575 7 2603 9
rect 3155 7 3183 9
rect 3735 7 3763 9
rect 4315 7 4343 9
rect 4895 7 4923 9
rect 5475 7 5503 9
rect 6055 7 6083 9
rect 6635 7 6663 9
<< nsubdiffcont >>
rect 255 4267 283 4269
rect 835 4267 863 4269
rect 1415 4267 1443 4269
rect 1995 4267 2023 4269
rect 2575 4267 2603 4269
rect 3155 4267 3183 4269
rect 3735 4267 3763 4269
rect 4315 4267 4343 4269
rect 4895 4267 4923 4269
rect 5475 4267 5503 4269
rect 6055 4267 6083 4269
rect 6635 4267 6663 4269
rect 255 3997 283 3999
rect 835 3997 863 3999
rect 1415 3997 1443 3999
rect 1995 3997 2023 3999
rect 2575 3997 2603 3999
rect 3155 3997 3183 3999
rect 3735 3997 3763 3999
rect 4315 3997 4343 3999
rect 4895 3997 4923 3999
rect 5475 3997 5503 3999
rect 6055 3997 6083 3999
rect 6635 3997 6663 3999
rect 255 3727 283 3729
rect 835 3727 863 3729
rect 1415 3727 1443 3729
rect 1995 3727 2023 3729
rect 2575 3727 2603 3729
rect 3155 3727 3183 3729
rect 3735 3727 3763 3729
rect 4315 3727 4343 3729
rect 4895 3727 4923 3729
rect 5475 3727 5503 3729
rect 6055 3727 6083 3729
rect 6635 3727 6663 3729
rect 255 3457 283 3459
rect 835 3457 863 3459
rect 1415 3457 1443 3459
rect 1995 3457 2023 3459
rect 2575 3457 2603 3459
rect 3155 3457 3183 3459
rect 3735 3457 3763 3459
rect 4315 3457 4343 3459
rect 4895 3457 4923 3459
rect 5475 3457 5503 3459
rect 6055 3457 6083 3459
rect 6635 3457 6663 3459
rect 255 3187 283 3189
rect 835 3187 863 3189
rect 1415 3187 1443 3189
rect 1995 3187 2023 3189
rect 2575 3187 2603 3189
rect 3155 3187 3183 3189
rect 3735 3187 3763 3189
rect 4315 3187 4343 3189
rect 4895 3187 4923 3189
rect 5475 3187 5503 3189
rect 6055 3187 6083 3189
rect 6635 3187 6663 3189
rect 255 2917 283 2919
rect 835 2917 863 2919
rect 1415 2917 1443 2919
rect 1995 2917 2023 2919
rect 2575 2917 2603 2919
rect 3155 2917 3183 2919
rect 3735 2917 3763 2919
rect 4315 2917 4343 2919
rect 4895 2917 4923 2919
rect 5475 2917 5503 2919
rect 6055 2917 6083 2919
rect 6635 2917 6663 2919
rect 255 2647 283 2649
rect 835 2647 863 2649
rect 1415 2647 1443 2649
rect 1995 2647 2023 2649
rect 2575 2647 2603 2649
rect 3155 2647 3183 2649
rect 3735 2647 3763 2649
rect 4315 2647 4343 2649
rect 4895 2647 4923 2649
rect 5475 2647 5503 2649
rect 6055 2647 6083 2649
rect 6635 2647 6663 2649
rect 255 2377 283 2379
rect 835 2377 863 2379
rect 1415 2377 1443 2379
rect 1995 2377 2023 2379
rect 2575 2377 2603 2379
rect 3155 2377 3183 2379
rect 3735 2377 3763 2379
rect 4315 2377 4343 2379
rect 4895 2377 4923 2379
rect 5475 2377 5503 2379
rect 6055 2377 6083 2379
rect 6635 2377 6663 2379
rect 255 2107 283 2109
rect 835 2107 863 2109
rect 1415 2107 1443 2109
rect 1995 2107 2023 2109
rect 2575 2107 2603 2109
rect 3155 2107 3183 2109
rect 3735 2107 3763 2109
rect 4315 2107 4343 2109
rect 4895 2107 4923 2109
rect 5475 2107 5503 2109
rect 6055 2107 6083 2109
rect 6635 2107 6663 2109
rect 255 1837 283 1839
rect 835 1837 863 1839
rect 1415 1837 1443 1839
rect 1995 1837 2023 1839
rect 2575 1837 2603 1839
rect 3155 1837 3183 1839
rect 3735 1837 3763 1839
rect 4315 1837 4343 1839
rect 4895 1837 4923 1839
rect 5475 1837 5503 1839
rect 6055 1837 6083 1839
rect 6635 1837 6663 1839
rect 255 1567 283 1569
rect 835 1567 863 1569
rect 1415 1567 1443 1569
rect 1995 1567 2023 1569
rect 2575 1567 2603 1569
rect 3155 1567 3183 1569
rect 3735 1567 3763 1569
rect 4315 1567 4343 1569
rect 4895 1567 4923 1569
rect 5475 1567 5503 1569
rect 6055 1567 6083 1569
rect 6635 1567 6663 1569
rect 255 1297 283 1299
rect 835 1297 863 1299
rect 1415 1297 1443 1299
rect 1995 1297 2023 1299
rect 2575 1297 2603 1299
rect 3155 1297 3183 1299
rect 3735 1297 3763 1299
rect 4315 1297 4343 1299
rect 4895 1297 4923 1299
rect 5475 1297 5503 1299
rect 6055 1297 6083 1299
rect 6635 1297 6663 1299
rect 255 1027 283 1029
rect 835 1027 863 1029
rect 1415 1027 1443 1029
rect 1995 1027 2023 1029
rect 2575 1027 2603 1029
rect 3155 1027 3183 1029
rect 3735 1027 3763 1029
rect 4315 1027 4343 1029
rect 4895 1027 4923 1029
rect 5475 1027 5503 1029
rect 6055 1027 6083 1029
rect 6635 1027 6663 1029
rect 255 757 283 759
rect 835 757 863 759
rect 1415 757 1443 759
rect 1995 757 2023 759
rect 2575 757 2603 759
rect 3155 757 3183 759
rect 3735 757 3763 759
rect 4315 757 4343 759
rect 4895 757 4923 759
rect 5475 757 5503 759
rect 6055 757 6083 759
rect 6635 757 6663 759
rect 255 487 283 489
rect 835 487 863 489
rect 1415 487 1443 489
rect 1995 487 2023 489
rect 2575 487 2603 489
rect 3155 487 3183 489
rect 3735 487 3763 489
rect 4315 487 4343 489
rect 4895 487 4923 489
rect 5475 487 5503 489
rect 6055 487 6083 489
rect 6635 487 6663 489
rect 255 217 283 219
rect 835 217 863 219
rect 1415 217 1443 219
rect 1995 217 2023 219
rect 2575 217 2603 219
rect 3155 217 3183 219
rect 3735 217 3763 219
rect 4315 217 4343 219
rect 4895 217 4923 219
rect 5475 217 5503 219
rect 6055 217 6083 219
rect 6635 217 6663 219
<< poly >>
rect -43 4283 6925 4313
rect 100 4255 130 4283
rect 215 4245 245 4267
rect 293 4245 323 4267
rect 408 4255 438 4283
rect 100 4205 130 4227
rect 680 4255 710 4283
rect 795 4245 825 4267
rect 873 4245 903 4267
rect 988 4255 1018 4283
rect 215 4184 245 4217
rect 36 4123 66 4145
rect 122 4123 137 4157
rect 215 4123 245 4150
rect 293 4184 323 4217
rect 408 4205 438 4227
rect 680 4205 710 4227
rect 1260 4255 1290 4283
rect 1375 4245 1405 4267
rect 1453 4245 1483 4267
rect 1568 4255 1598 4283
rect 795 4184 825 4217
rect 293 4123 323 4150
rect 401 4123 416 4157
rect 472 4123 502 4145
rect 616 4123 646 4145
rect 702 4123 717 4157
rect 795 4123 825 4150
rect 873 4184 903 4217
rect 988 4205 1018 4227
rect 1260 4205 1290 4227
rect 1840 4255 1870 4283
rect 1955 4245 1985 4267
rect 2033 4245 2063 4267
rect 2148 4255 2178 4283
rect 1375 4184 1405 4217
rect 873 4123 903 4150
rect 981 4123 996 4157
rect 1052 4123 1082 4145
rect 1196 4123 1226 4145
rect 1282 4123 1297 4157
rect 1375 4123 1405 4150
rect 1453 4184 1483 4217
rect 1568 4205 1598 4227
rect 1840 4205 1870 4227
rect 2420 4255 2450 4283
rect 2535 4245 2565 4267
rect 2613 4245 2643 4267
rect 2728 4255 2758 4283
rect 1955 4184 1985 4217
rect 1453 4123 1483 4150
rect 1561 4123 1576 4157
rect 1632 4123 1662 4145
rect 1776 4123 1806 4145
rect 1862 4123 1877 4157
rect 1955 4123 1985 4150
rect 2033 4184 2063 4217
rect 2148 4205 2178 4227
rect 2420 4205 2450 4227
rect 3000 4255 3030 4283
rect 3115 4245 3145 4267
rect 3193 4245 3223 4267
rect 3308 4255 3338 4283
rect 2535 4184 2565 4217
rect 2033 4123 2063 4150
rect 2141 4123 2156 4157
rect 2212 4123 2242 4145
rect 2356 4123 2386 4145
rect 2442 4123 2457 4157
rect 2535 4123 2565 4150
rect 2613 4184 2643 4217
rect 2728 4205 2758 4227
rect 3000 4205 3030 4227
rect 3580 4255 3610 4283
rect 3695 4245 3725 4267
rect 3773 4245 3803 4267
rect 3888 4255 3918 4283
rect 3115 4184 3145 4217
rect 2613 4123 2643 4150
rect 2721 4123 2736 4157
rect 2792 4123 2822 4145
rect 2936 4123 2966 4145
rect 3022 4123 3037 4157
rect 3115 4123 3145 4150
rect 3193 4184 3223 4217
rect 3308 4205 3338 4227
rect 3580 4205 3610 4227
rect 4160 4255 4190 4283
rect 4275 4245 4305 4267
rect 4353 4245 4383 4267
rect 4468 4255 4498 4283
rect 3695 4184 3725 4217
rect 3193 4123 3223 4150
rect 3301 4123 3316 4157
rect 3372 4123 3402 4145
rect 3516 4123 3546 4145
rect 3602 4123 3617 4157
rect 3695 4123 3725 4150
rect 3773 4184 3803 4217
rect 3888 4205 3918 4227
rect 4160 4205 4190 4227
rect 4740 4255 4770 4283
rect 4855 4245 4885 4267
rect 4933 4245 4963 4267
rect 5048 4255 5078 4283
rect 4275 4184 4305 4217
rect 3773 4123 3803 4150
rect 3881 4123 3896 4157
rect 3952 4123 3982 4145
rect 4096 4123 4126 4145
rect 4182 4123 4197 4157
rect 4275 4123 4305 4150
rect 4353 4184 4383 4217
rect 4468 4205 4498 4227
rect 4740 4205 4770 4227
rect 5320 4255 5350 4283
rect 5435 4245 5465 4267
rect 5513 4245 5543 4267
rect 5628 4255 5658 4283
rect 4855 4184 4885 4217
rect 4353 4123 4383 4150
rect 4461 4123 4476 4157
rect 4532 4123 4562 4145
rect 4676 4123 4706 4145
rect 4762 4123 4777 4157
rect 4855 4123 4885 4150
rect 4933 4184 4963 4217
rect 5048 4205 5078 4227
rect 5320 4205 5350 4227
rect 5900 4255 5930 4283
rect 6015 4245 6045 4267
rect 6093 4245 6123 4267
rect 6208 4255 6238 4283
rect 5435 4184 5465 4217
rect 4933 4123 4963 4150
rect 5041 4123 5056 4157
rect 5112 4123 5142 4145
rect 5256 4123 5286 4145
rect 5342 4123 5357 4157
rect 5435 4123 5465 4150
rect 5513 4184 5543 4217
rect 5628 4205 5658 4227
rect 5900 4205 5930 4227
rect 6480 4255 6510 4283
rect 6595 4245 6625 4267
rect 6673 4245 6703 4267
rect 6788 4255 6818 4283
rect 6015 4184 6045 4217
rect 5513 4123 5543 4150
rect 5621 4123 5636 4157
rect 5692 4123 5722 4145
rect 5836 4123 5866 4145
rect 5922 4123 5937 4157
rect 6015 4123 6045 4150
rect 6093 4184 6123 4217
rect 6208 4205 6238 4227
rect 6480 4205 6510 4227
rect 6595 4184 6625 4217
rect 6093 4123 6123 4150
rect 6201 4123 6216 4157
rect 6272 4123 6302 4145
rect 6416 4123 6446 4145
rect 6502 4123 6517 4157
rect 6595 4123 6625 4150
rect 6673 4184 6703 4217
rect 6788 4205 6818 4227
rect 6673 4123 6703 4150
rect 6781 4123 6796 4157
rect 6852 4123 6882 4145
rect 122 4109 152 4123
rect 386 4109 416 4123
rect 702 4109 732 4123
rect 966 4109 996 4123
rect 1282 4109 1312 4123
rect 1546 4109 1576 4123
rect 1862 4109 1892 4123
rect 2126 4109 2156 4123
rect 2442 4109 2472 4123
rect 2706 4109 2736 4123
rect 3022 4109 3052 4123
rect 3286 4109 3316 4123
rect 3602 4109 3632 4123
rect 3866 4109 3896 4123
rect 4182 4109 4212 4123
rect 4446 4109 4476 4123
rect 4762 4109 4792 4123
rect 5026 4109 5056 4123
rect 5342 4109 5372 4123
rect 5606 4109 5636 4123
rect 5922 4109 5952 4123
rect 6186 4109 6216 4123
rect 6502 4109 6532 4123
rect 6766 4109 6796 4123
rect 36 4059 66 4081
rect 122 4059 152 4081
rect 215 4059 245 4081
rect 293 4059 323 4081
rect 386 4059 416 4081
rect 472 4059 502 4081
rect 616 4059 646 4081
rect 702 4059 732 4081
rect 795 4059 825 4081
rect 873 4059 903 4081
rect 966 4059 996 4081
rect 1052 4059 1082 4081
rect 1196 4059 1226 4081
rect 1282 4059 1312 4081
rect 1375 4059 1405 4081
rect 1453 4059 1483 4081
rect 1546 4059 1576 4081
rect 1632 4059 1662 4081
rect 1776 4059 1806 4081
rect 1862 4059 1892 4081
rect 1955 4059 1985 4081
rect 2033 4059 2063 4081
rect 2126 4059 2156 4081
rect 2212 4059 2242 4081
rect 2356 4059 2386 4081
rect 2442 4059 2472 4081
rect 2535 4059 2565 4081
rect 2613 4059 2643 4081
rect 2706 4059 2736 4081
rect 2792 4059 2822 4081
rect 2936 4059 2966 4081
rect 3022 4059 3052 4081
rect 3115 4059 3145 4081
rect 3193 4059 3223 4081
rect 3286 4059 3316 4081
rect 3372 4059 3402 4081
rect 3516 4059 3546 4081
rect 3602 4059 3632 4081
rect 3695 4059 3725 4081
rect 3773 4059 3803 4081
rect 3866 4059 3896 4081
rect 3952 4059 3982 4081
rect 4096 4059 4126 4081
rect 4182 4059 4212 4081
rect 4275 4059 4305 4081
rect 4353 4059 4383 4081
rect 4446 4059 4476 4081
rect 4532 4059 4562 4081
rect 4676 4059 4706 4081
rect 4762 4059 4792 4081
rect 4855 4059 4885 4081
rect 4933 4059 4963 4081
rect 5026 4059 5056 4081
rect 5112 4059 5142 4081
rect 5256 4059 5286 4081
rect 5342 4059 5372 4081
rect 5435 4059 5465 4081
rect 5513 4059 5543 4081
rect 5606 4059 5636 4081
rect 5692 4059 5722 4081
rect 5836 4059 5866 4081
rect 5922 4059 5952 4081
rect 6015 4059 6045 4081
rect 6093 4059 6123 4081
rect 6186 4059 6216 4081
rect 6272 4059 6302 4081
rect 6416 4059 6446 4081
rect 6502 4059 6532 4081
rect 6595 4059 6625 4081
rect 6673 4059 6703 4081
rect 6766 4059 6796 4081
rect 6852 4059 6882 4081
rect -43 4013 6925 4043
rect 100 3985 130 4013
rect 215 3975 245 3997
rect 293 3975 323 3997
rect 408 3985 438 4013
rect 100 3935 130 3957
rect 680 3985 710 4013
rect 795 3975 825 3997
rect 873 3975 903 3997
rect 988 3985 1018 4013
rect 215 3914 245 3947
rect 36 3853 66 3875
rect 122 3853 137 3887
rect 215 3853 245 3880
rect 293 3914 323 3947
rect 408 3935 438 3957
rect 680 3935 710 3957
rect 1260 3985 1290 4013
rect 1375 3975 1405 3997
rect 1453 3975 1483 3997
rect 1568 3985 1598 4013
rect 795 3914 825 3947
rect 293 3853 323 3880
rect 401 3853 416 3887
rect 472 3853 502 3875
rect 616 3853 646 3875
rect 702 3853 717 3887
rect 795 3853 825 3880
rect 873 3914 903 3947
rect 988 3935 1018 3957
rect 1260 3935 1290 3957
rect 1840 3985 1870 4013
rect 1955 3975 1985 3997
rect 2033 3975 2063 3997
rect 2148 3985 2178 4013
rect 1375 3914 1405 3947
rect 873 3853 903 3880
rect 981 3853 996 3887
rect 1052 3853 1082 3875
rect 1196 3853 1226 3875
rect 1282 3853 1297 3887
rect 1375 3853 1405 3880
rect 1453 3914 1483 3947
rect 1568 3935 1598 3957
rect 1840 3935 1870 3957
rect 2420 3985 2450 4013
rect 2535 3975 2565 3997
rect 2613 3975 2643 3997
rect 2728 3985 2758 4013
rect 1955 3914 1985 3947
rect 1453 3853 1483 3880
rect 1561 3853 1576 3887
rect 1632 3853 1662 3875
rect 1776 3853 1806 3875
rect 1862 3853 1877 3887
rect 1955 3853 1985 3880
rect 2033 3914 2063 3947
rect 2148 3935 2178 3957
rect 2420 3935 2450 3957
rect 3000 3985 3030 4013
rect 3115 3975 3145 3997
rect 3193 3975 3223 3997
rect 3308 3985 3338 4013
rect 2535 3914 2565 3947
rect 2033 3853 2063 3880
rect 2141 3853 2156 3887
rect 2212 3853 2242 3875
rect 2356 3853 2386 3875
rect 2442 3853 2457 3887
rect 2535 3853 2565 3880
rect 2613 3914 2643 3947
rect 2728 3935 2758 3957
rect 3000 3935 3030 3957
rect 3580 3985 3610 4013
rect 3695 3975 3725 3997
rect 3773 3975 3803 3997
rect 3888 3985 3918 4013
rect 3115 3914 3145 3947
rect 2613 3853 2643 3880
rect 2721 3853 2736 3887
rect 2792 3853 2822 3875
rect 2936 3853 2966 3875
rect 3022 3853 3037 3887
rect 3115 3853 3145 3880
rect 3193 3914 3223 3947
rect 3308 3935 3338 3957
rect 3580 3935 3610 3957
rect 4160 3985 4190 4013
rect 4275 3975 4305 3997
rect 4353 3975 4383 3997
rect 4468 3985 4498 4013
rect 3695 3914 3725 3947
rect 3193 3853 3223 3880
rect 3301 3853 3316 3887
rect 3372 3853 3402 3875
rect 3516 3853 3546 3875
rect 3602 3853 3617 3887
rect 3695 3853 3725 3880
rect 3773 3914 3803 3947
rect 3888 3935 3918 3957
rect 4160 3935 4190 3957
rect 4740 3985 4770 4013
rect 4855 3975 4885 3997
rect 4933 3975 4963 3997
rect 5048 3985 5078 4013
rect 4275 3914 4305 3947
rect 3773 3853 3803 3880
rect 3881 3853 3896 3887
rect 3952 3853 3982 3875
rect 4096 3853 4126 3875
rect 4182 3853 4197 3887
rect 4275 3853 4305 3880
rect 4353 3914 4383 3947
rect 4468 3935 4498 3957
rect 4740 3935 4770 3957
rect 5320 3985 5350 4013
rect 5435 3975 5465 3997
rect 5513 3975 5543 3997
rect 5628 3985 5658 4013
rect 4855 3914 4885 3947
rect 4353 3853 4383 3880
rect 4461 3853 4476 3887
rect 4532 3853 4562 3875
rect 4676 3853 4706 3875
rect 4762 3853 4777 3887
rect 4855 3853 4885 3880
rect 4933 3914 4963 3947
rect 5048 3935 5078 3957
rect 5320 3935 5350 3957
rect 5900 3985 5930 4013
rect 6015 3975 6045 3997
rect 6093 3975 6123 3997
rect 6208 3985 6238 4013
rect 5435 3914 5465 3947
rect 4933 3853 4963 3880
rect 5041 3853 5056 3887
rect 5112 3853 5142 3875
rect 5256 3853 5286 3875
rect 5342 3853 5357 3887
rect 5435 3853 5465 3880
rect 5513 3914 5543 3947
rect 5628 3935 5658 3957
rect 5900 3935 5930 3957
rect 6480 3985 6510 4013
rect 6595 3975 6625 3997
rect 6673 3975 6703 3997
rect 6788 3985 6818 4013
rect 6015 3914 6045 3947
rect 5513 3853 5543 3880
rect 5621 3853 5636 3887
rect 5692 3853 5722 3875
rect 5836 3853 5866 3875
rect 5922 3853 5937 3887
rect 6015 3853 6045 3880
rect 6093 3914 6123 3947
rect 6208 3935 6238 3957
rect 6480 3935 6510 3957
rect 6595 3914 6625 3947
rect 6093 3853 6123 3880
rect 6201 3853 6216 3887
rect 6272 3853 6302 3875
rect 6416 3853 6446 3875
rect 6502 3853 6517 3887
rect 6595 3853 6625 3880
rect 6673 3914 6703 3947
rect 6788 3935 6818 3957
rect 6673 3853 6703 3880
rect 6781 3853 6796 3887
rect 6852 3853 6882 3875
rect 122 3839 152 3853
rect 386 3839 416 3853
rect 702 3839 732 3853
rect 966 3839 996 3853
rect 1282 3839 1312 3853
rect 1546 3839 1576 3853
rect 1862 3839 1892 3853
rect 2126 3839 2156 3853
rect 2442 3839 2472 3853
rect 2706 3839 2736 3853
rect 3022 3839 3052 3853
rect 3286 3839 3316 3853
rect 3602 3839 3632 3853
rect 3866 3839 3896 3853
rect 4182 3839 4212 3853
rect 4446 3839 4476 3853
rect 4762 3839 4792 3853
rect 5026 3839 5056 3853
rect 5342 3839 5372 3853
rect 5606 3839 5636 3853
rect 5922 3839 5952 3853
rect 6186 3839 6216 3853
rect 6502 3839 6532 3853
rect 6766 3839 6796 3853
rect 36 3789 66 3811
rect 122 3789 152 3811
rect 215 3789 245 3811
rect 293 3789 323 3811
rect 386 3789 416 3811
rect 472 3789 502 3811
rect 616 3789 646 3811
rect 702 3789 732 3811
rect 795 3789 825 3811
rect 873 3789 903 3811
rect 966 3789 996 3811
rect 1052 3789 1082 3811
rect 1196 3789 1226 3811
rect 1282 3789 1312 3811
rect 1375 3789 1405 3811
rect 1453 3789 1483 3811
rect 1546 3789 1576 3811
rect 1632 3789 1662 3811
rect 1776 3789 1806 3811
rect 1862 3789 1892 3811
rect 1955 3789 1985 3811
rect 2033 3789 2063 3811
rect 2126 3789 2156 3811
rect 2212 3789 2242 3811
rect 2356 3789 2386 3811
rect 2442 3789 2472 3811
rect 2535 3789 2565 3811
rect 2613 3789 2643 3811
rect 2706 3789 2736 3811
rect 2792 3789 2822 3811
rect 2936 3789 2966 3811
rect 3022 3789 3052 3811
rect 3115 3789 3145 3811
rect 3193 3789 3223 3811
rect 3286 3789 3316 3811
rect 3372 3789 3402 3811
rect 3516 3789 3546 3811
rect 3602 3789 3632 3811
rect 3695 3789 3725 3811
rect 3773 3789 3803 3811
rect 3866 3789 3896 3811
rect 3952 3789 3982 3811
rect 4096 3789 4126 3811
rect 4182 3789 4212 3811
rect 4275 3789 4305 3811
rect 4353 3789 4383 3811
rect 4446 3789 4476 3811
rect 4532 3789 4562 3811
rect 4676 3789 4706 3811
rect 4762 3789 4792 3811
rect 4855 3789 4885 3811
rect 4933 3789 4963 3811
rect 5026 3789 5056 3811
rect 5112 3789 5142 3811
rect 5256 3789 5286 3811
rect 5342 3789 5372 3811
rect 5435 3789 5465 3811
rect 5513 3789 5543 3811
rect 5606 3789 5636 3811
rect 5692 3789 5722 3811
rect 5836 3789 5866 3811
rect 5922 3789 5952 3811
rect 6015 3789 6045 3811
rect 6093 3789 6123 3811
rect 6186 3789 6216 3811
rect 6272 3789 6302 3811
rect 6416 3789 6446 3811
rect 6502 3789 6532 3811
rect 6595 3789 6625 3811
rect 6673 3789 6703 3811
rect 6766 3789 6796 3811
rect 6852 3789 6882 3811
rect -43 3743 6925 3773
rect 100 3715 130 3743
rect 215 3705 245 3727
rect 293 3705 323 3727
rect 408 3715 438 3743
rect 100 3665 130 3687
rect 680 3715 710 3743
rect 795 3705 825 3727
rect 873 3705 903 3727
rect 988 3715 1018 3743
rect 215 3644 245 3677
rect 36 3583 66 3605
rect 122 3583 137 3617
rect 215 3583 245 3610
rect 293 3644 323 3677
rect 408 3665 438 3687
rect 680 3665 710 3687
rect 1260 3715 1290 3743
rect 1375 3705 1405 3727
rect 1453 3705 1483 3727
rect 1568 3715 1598 3743
rect 795 3644 825 3677
rect 293 3583 323 3610
rect 401 3583 416 3617
rect 472 3583 502 3605
rect 616 3583 646 3605
rect 702 3583 717 3617
rect 795 3583 825 3610
rect 873 3644 903 3677
rect 988 3665 1018 3687
rect 1260 3665 1290 3687
rect 1840 3715 1870 3743
rect 1955 3705 1985 3727
rect 2033 3705 2063 3727
rect 2148 3715 2178 3743
rect 1375 3644 1405 3677
rect 873 3583 903 3610
rect 981 3583 996 3617
rect 1052 3583 1082 3605
rect 1196 3583 1226 3605
rect 1282 3583 1297 3617
rect 1375 3583 1405 3610
rect 1453 3644 1483 3677
rect 1568 3665 1598 3687
rect 1840 3665 1870 3687
rect 2420 3715 2450 3743
rect 2535 3705 2565 3727
rect 2613 3705 2643 3727
rect 2728 3715 2758 3743
rect 1955 3644 1985 3677
rect 1453 3583 1483 3610
rect 1561 3583 1576 3617
rect 1632 3583 1662 3605
rect 1776 3583 1806 3605
rect 1862 3583 1877 3617
rect 1955 3583 1985 3610
rect 2033 3644 2063 3677
rect 2148 3665 2178 3687
rect 2420 3665 2450 3687
rect 3000 3715 3030 3743
rect 3115 3705 3145 3727
rect 3193 3705 3223 3727
rect 3308 3715 3338 3743
rect 2535 3644 2565 3677
rect 2033 3583 2063 3610
rect 2141 3583 2156 3617
rect 2212 3583 2242 3605
rect 2356 3583 2386 3605
rect 2442 3583 2457 3617
rect 2535 3583 2565 3610
rect 2613 3644 2643 3677
rect 2728 3665 2758 3687
rect 3000 3665 3030 3687
rect 3580 3715 3610 3743
rect 3695 3705 3725 3727
rect 3773 3705 3803 3727
rect 3888 3715 3918 3743
rect 3115 3644 3145 3677
rect 2613 3583 2643 3610
rect 2721 3583 2736 3617
rect 2792 3583 2822 3605
rect 2936 3583 2966 3605
rect 3022 3583 3037 3617
rect 3115 3583 3145 3610
rect 3193 3644 3223 3677
rect 3308 3665 3338 3687
rect 3580 3665 3610 3687
rect 4160 3715 4190 3743
rect 4275 3705 4305 3727
rect 4353 3705 4383 3727
rect 4468 3715 4498 3743
rect 3695 3644 3725 3677
rect 3193 3583 3223 3610
rect 3301 3583 3316 3617
rect 3372 3583 3402 3605
rect 3516 3583 3546 3605
rect 3602 3583 3617 3617
rect 3695 3583 3725 3610
rect 3773 3644 3803 3677
rect 3888 3665 3918 3687
rect 4160 3665 4190 3687
rect 4740 3715 4770 3743
rect 4855 3705 4885 3727
rect 4933 3705 4963 3727
rect 5048 3715 5078 3743
rect 4275 3644 4305 3677
rect 3773 3583 3803 3610
rect 3881 3583 3896 3617
rect 3952 3583 3982 3605
rect 4096 3583 4126 3605
rect 4182 3583 4197 3617
rect 4275 3583 4305 3610
rect 4353 3644 4383 3677
rect 4468 3665 4498 3687
rect 4740 3665 4770 3687
rect 5320 3715 5350 3743
rect 5435 3705 5465 3727
rect 5513 3705 5543 3727
rect 5628 3715 5658 3743
rect 4855 3644 4885 3677
rect 4353 3583 4383 3610
rect 4461 3583 4476 3617
rect 4532 3583 4562 3605
rect 4676 3583 4706 3605
rect 4762 3583 4777 3617
rect 4855 3583 4885 3610
rect 4933 3644 4963 3677
rect 5048 3665 5078 3687
rect 5320 3665 5350 3687
rect 5900 3715 5930 3743
rect 6015 3705 6045 3727
rect 6093 3705 6123 3727
rect 6208 3715 6238 3743
rect 5435 3644 5465 3677
rect 4933 3583 4963 3610
rect 5041 3583 5056 3617
rect 5112 3583 5142 3605
rect 5256 3583 5286 3605
rect 5342 3583 5357 3617
rect 5435 3583 5465 3610
rect 5513 3644 5543 3677
rect 5628 3665 5658 3687
rect 5900 3665 5930 3687
rect 6480 3715 6510 3743
rect 6595 3705 6625 3727
rect 6673 3705 6703 3727
rect 6788 3715 6818 3743
rect 6015 3644 6045 3677
rect 5513 3583 5543 3610
rect 5621 3583 5636 3617
rect 5692 3583 5722 3605
rect 5836 3583 5866 3605
rect 5922 3583 5937 3617
rect 6015 3583 6045 3610
rect 6093 3644 6123 3677
rect 6208 3665 6238 3687
rect 6480 3665 6510 3687
rect 6595 3644 6625 3677
rect 6093 3583 6123 3610
rect 6201 3583 6216 3617
rect 6272 3583 6302 3605
rect 6416 3583 6446 3605
rect 6502 3583 6517 3617
rect 6595 3583 6625 3610
rect 6673 3644 6703 3677
rect 6788 3665 6818 3687
rect 6673 3583 6703 3610
rect 6781 3583 6796 3617
rect 6852 3583 6882 3605
rect 122 3569 152 3583
rect 386 3569 416 3583
rect 702 3569 732 3583
rect 966 3569 996 3583
rect 1282 3569 1312 3583
rect 1546 3569 1576 3583
rect 1862 3569 1892 3583
rect 2126 3569 2156 3583
rect 2442 3569 2472 3583
rect 2706 3569 2736 3583
rect 3022 3569 3052 3583
rect 3286 3569 3316 3583
rect 3602 3569 3632 3583
rect 3866 3569 3896 3583
rect 4182 3569 4212 3583
rect 4446 3569 4476 3583
rect 4762 3569 4792 3583
rect 5026 3569 5056 3583
rect 5342 3569 5372 3583
rect 5606 3569 5636 3583
rect 5922 3569 5952 3583
rect 6186 3569 6216 3583
rect 6502 3569 6532 3583
rect 6766 3569 6796 3583
rect 36 3519 66 3541
rect 122 3519 152 3541
rect 215 3519 245 3541
rect 293 3519 323 3541
rect 386 3519 416 3541
rect 472 3519 502 3541
rect 616 3519 646 3541
rect 702 3519 732 3541
rect 795 3519 825 3541
rect 873 3519 903 3541
rect 966 3519 996 3541
rect 1052 3519 1082 3541
rect 1196 3519 1226 3541
rect 1282 3519 1312 3541
rect 1375 3519 1405 3541
rect 1453 3519 1483 3541
rect 1546 3519 1576 3541
rect 1632 3519 1662 3541
rect 1776 3519 1806 3541
rect 1862 3519 1892 3541
rect 1955 3519 1985 3541
rect 2033 3519 2063 3541
rect 2126 3519 2156 3541
rect 2212 3519 2242 3541
rect 2356 3519 2386 3541
rect 2442 3519 2472 3541
rect 2535 3519 2565 3541
rect 2613 3519 2643 3541
rect 2706 3519 2736 3541
rect 2792 3519 2822 3541
rect 2936 3519 2966 3541
rect 3022 3519 3052 3541
rect 3115 3519 3145 3541
rect 3193 3519 3223 3541
rect 3286 3519 3316 3541
rect 3372 3519 3402 3541
rect 3516 3519 3546 3541
rect 3602 3519 3632 3541
rect 3695 3519 3725 3541
rect 3773 3519 3803 3541
rect 3866 3519 3896 3541
rect 3952 3519 3982 3541
rect 4096 3519 4126 3541
rect 4182 3519 4212 3541
rect 4275 3519 4305 3541
rect 4353 3519 4383 3541
rect 4446 3519 4476 3541
rect 4532 3519 4562 3541
rect 4676 3519 4706 3541
rect 4762 3519 4792 3541
rect 4855 3519 4885 3541
rect 4933 3519 4963 3541
rect 5026 3519 5056 3541
rect 5112 3519 5142 3541
rect 5256 3519 5286 3541
rect 5342 3519 5372 3541
rect 5435 3519 5465 3541
rect 5513 3519 5543 3541
rect 5606 3519 5636 3541
rect 5692 3519 5722 3541
rect 5836 3519 5866 3541
rect 5922 3519 5952 3541
rect 6015 3519 6045 3541
rect 6093 3519 6123 3541
rect 6186 3519 6216 3541
rect 6272 3519 6302 3541
rect 6416 3519 6446 3541
rect 6502 3519 6532 3541
rect 6595 3519 6625 3541
rect 6673 3519 6703 3541
rect 6766 3519 6796 3541
rect 6852 3519 6882 3541
rect -43 3473 6925 3503
rect 100 3445 130 3473
rect 215 3435 245 3457
rect 293 3435 323 3457
rect 408 3445 438 3473
rect 100 3395 130 3417
rect 680 3445 710 3473
rect 795 3435 825 3457
rect 873 3435 903 3457
rect 988 3445 1018 3473
rect 215 3374 245 3407
rect 36 3313 66 3335
rect 122 3313 137 3347
rect 215 3313 245 3340
rect 293 3374 323 3407
rect 408 3395 438 3417
rect 680 3395 710 3417
rect 1260 3445 1290 3473
rect 1375 3435 1405 3457
rect 1453 3435 1483 3457
rect 1568 3445 1598 3473
rect 795 3374 825 3407
rect 293 3313 323 3340
rect 401 3313 416 3347
rect 472 3313 502 3335
rect 616 3313 646 3335
rect 702 3313 717 3347
rect 795 3313 825 3340
rect 873 3374 903 3407
rect 988 3395 1018 3417
rect 1260 3395 1290 3417
rect 1840 3445 1870 3473
rect 1955 3435 1985 3457
rect 2033 3435 2063 3457
rect 2148 3445 2178 3473
rect 1375 3374 1405 3407
rect 873 3313 903 3340
rect 981 3313 996 3347
rect 1052 3313 1082 3335
rect 1196 3313 1226 3335
rect 1282 3313 1297 3347
rect 1375 3313 1405 3340
rect 1453 3374 1483 3407
rect 1568 3395 1598 3417
rect 1840 3395 1870 3417
rect 2420 3445 2450 3473
rect 2535 3435 2565 3457
rect 2613 3435 2643 3457
rect 2728 3445 2758 3473
rect 1955 3374 1985 3407
rect 1453 3313 1483 3340
rect 1561 3313 1576 3347
rect 1632 3313 1662 3335
rect 1776 3313 1806 3335
rect 1862 3313 1877 3347
rect 1955 3313 1985 3340
rect 2033 3374 2063 3407
rect 2148 3395 2178 3417
rect 2420 3395 2450 3417
rect 3000 3445 3030 3473
rect 3115 3435 3145 3457
rect 3193 3435 3223 3457
rect 3308 3445 3338 3473
rect 2535 3374 2565 3407
rect 2033 3313 2063 3340
rect 2141 3313 2156 3347
rect 2212 3313 2242 3335
rect 2356 3313 2386 3335
rect 2442 3313 2457 3347
rect 2535 3313 2565 3340
rect 2613 3374 2643 3407
rect 2728 3395 2758 3417
rect 3000 3395 3030 3417
rect 3580 3445 3610 3473
rect 3695 3435 3725 3457
rect 3773 3435 3803 3457
rect 3888 3445 3918 3473
rect 3115 3374 3145 3407
rect 2613 3313 2643 3340
rect 2721 3313 2736 3347
rect 2792 3313 2822 3335
rect 2936 3313 2966 3335
rect 3022 3313 3037 3347
rect 3115 3313 3145 3340
rect 3193 3374 3223 3407
rect 3308 3395 3338 3417
rect 3580 3395 3610 3417
rect 4160 3445 4190 3473
rect 4275 3435 4305 3457
rect 4353 3435 4383 3457
rect 4468 3445 4498 3473
rect 3695 3374 3725 3407
rect 3193 3313 3223 3340
rect 3301 3313 3316 3347
rect 3372 3313 3402 3335
rect 3516 3313 3546 3335
rect 3602 3313 3617 3347
rect 3695 3313 3725 3340
rect 3773 3374 3803 3407
rect 3888 3395 3918 3417
rect 4160 3395 4190 3417
rect 4740 3445 4770 3473
rect 4855 3435 4885 3457
rect 4933 3435 4963 3457
rect 5048 3445 5078 3473
rect 4275 3374 4305 3407
rect 3773 3313 3803 3340
rect 3881 3313 3896 3347
rect 3952 3313 3982 3335
rect 4096 3313 4126 3335
rect 4182 3313 4197 3347
rect 4275 3313 4305 3340
rect 4353 3374 4383 3407
rect 4468 3395 4498 3417
rect 4740 3395 4770 3417
rect 5320 3445 5350 3473
rect 5435 3435 5465 3457
rect 5513 3435 5543 3457
rect 5628 3445 5658 3473
rect 4855 3374 4885 3407
rect 4353 3313 4383 3340
rect 4461 3313 4476 3347
rect 4532 3313 4562 3335
rect 4676 3313 4706 3335
rect 4762 3313 4777 3347
rect 4855 3313 4885 3340
rect 4933 3374 4963 3407
rect 5048 3395 5078 3417
rect 5320 3395 5350 3417
rect 5900 3445 5930 3473
rect 6015 3435 6045 3457
rect 6093 3435 6123 3457
rect 6208 3445 6238 3473
rect 5435 3374 5465 3407
rect 4933 3313 4963 3340
rect 5041 3313 5056 3347
rect 5112 3313 5142 3335
rect 5256 3313 5286 3335
rect 5342 3313 5357 3347
rect 5435 3313 5465 3340
rect 5513 3374 5543 3407
rect 5628 3395 5658 3417
rect 5900 3395 5930 3417
rect 6480 3445 6510 3473
rect 6595 3435 6625 3457
rect 6673 3435 6703 3457
rect 6788 3445 6818 3473
rect 6015 3374 6045 3407
rect 5513 3313 5543 3340
rect 5621 3313 5636 3347
rect 5692 3313 5722 3335
rect 5836 3313 5866 3335
rect 5922 3313 5937 3347
rect 6015 3313 6045 3340
rect 6093 3374 6123 3407
rect 6208 3395 6238 3417
rect 6480 3395 6510 3417
rect 6595 3374 6625 3407
rect 6093 3313 6123 3340
rect 6201 3313 6216 3347
rect 6272 3313 6302 3335
rect 6416 3313 6446 3335
rect 6502 3313 6517 3347
rect 6595 3313 6625 3340
rect 6673 3374 6703 3407
rect 6788 3395 6818 3417
rect 6673 3313 6703 3340
rect 6781 3313 6796 3347
rect 6852 3313 6882 3335
rect 122 3299 152 3313
rect 386 3299 416 3313
rect 702 3299 732 3313
rect 966 3299 996 3313
rect 1282 3299 1312 3313
rect 1546 3299 1576 3313
rect 1862 3299 1892 3313
rect 2126 3299 2156 3313
rect 2442 3299 2472 3313
rect 2706 3299 2736 3313
rect 3022 3299 3052 3313
rect 3286 3299 3316 3313
rect 3602 3299 3632 3313
rect 3866 3299 3896 3313
rect 4182 3299 4212 3313
rect 4446 3299 4476 3313
rect 4762 3299 4792 3313
rect 5026 3299 5056 3313
rect 5342 3299 5372 3313
rect 5606 3299 5636 3313
rect 5922 3299 5952 3313
rect 6186 3299 6216 3313
rect 6502 3299 6532 3313
rect 6766 3299 6796 3313
rect 36 3249 66 3271
rect 122 3249 152 3271
rect 215 3249 245 3271
rect 293 3249 323 3271
rect 386 3249 416 3271
rect 472 3249 502 3271
rect 616 3249 646 3271
rect 702 3249 732 3271
rect 795 3249 825 3271
rect 873 3249 903 3271
rect 966 3249 996 3271
rect 1052 3249 1082 3271
rect 1196 3249 1226 3271
rect 1282 3249 1312 3271
rect 1375 3249 1405 3271
rect 1453 3249 1483 3271
rect 1546 3249 1576 3271
rect 1632 3249 1662 3271
rect 1776 3249 1806 3271
rect 1862 3249 1892 3271
rect 1955 3249 1985 3271
rect 2033 3249 2063 3271
rect 2126 3249 2156 3271
rect 2212 3249 2242 3271
rect 2356 3249 2386 3271
rect 2442 3249 2472 3271
rect 2535 3249 2565 3271
rect 2613 3249 2643 3271
rect 2706 3249 2736 3271
rect 2792 3249 2822 3271
rect 2936 3249 2966 3271
rect 3022 3249 3052 3271
rect 3115 3249 3145 3271
rect 3193 3249 3223 3271
rect 3286 3249 3316 3271
rect 3372 3249 3402 3271
rect 3516 3249 3546 3271
rect 3602 3249 3632 3271
rect 3695 3249 3725 3271
rect 3773 3249 3803 3271
rect 3866 3249 3896 3271
rect 3952 3249 3982 3271
rect 4096 3249 4126 3271
rect 4182 3249 4212 3271
rect 4275 3249 4305 3271
rect 4353 3249 4383 3271
rect 4446 3249 4476 3271
rect 4532 3249 4562 3271
rect 4676 3249 4706 3271
rect 4762 3249 4792 3271
rect 4855 3249 4885 3271
rect 4933 3249 4963 3271
rect 5026 3249 5056 3271
rect 5112 3249 5142 3271
rect 5256 3249 5286 3271
rect 5342 3249 5372 3271
rect 5435 3249 5465 3271
rect 5513 3249 5543 3271
rect 5606 3249 5636 3271
rect 5692 3249 5722 3271
rect 5836 3249 5866 3271
rect 5922 3249 5952 3271
rect 6015 3249 6045 3271
rect 6093 3249 6123 3271
rect 6186 3249 6216 3271
rect 6272 3249 6302 3271
rect 6416 3249 6446 3271
rect 6502 3249 6532 3271
rect 6595 3249 6625 3271
rect 6673 3249 6703 3271
rect 6766 3249 6796 3271
rect 6852 3249 6882 3271
rect -43 3203 6925 3233
rect 100 3175 130 3203
rect 215 3165 245 3187
rect 293 3165 323 3187
rect 408 3175 438 3203
rect 100 3125 130 3147
rect 680 3175 710 3203
rect 795 3165 825 3187
rect 873 3165 903 3187
rect 988 3175 1018 3203
rect 215 3104 245 3137
rect 36 3043 66 3065
rect 122 3043 137 3077
rect 215 3043 245 3070
rect 293 3104 323 3137
rect 408 3125 438 3147
rect 680 3125 710 3147
rect 1260 3175 1290 3203
rect 1375 3165 1405 3187
rect 1453 3165 1483 3187
rect 1568 3175 1598 3203
rect 795 3104 825 3137
rect 293 3043 323 3070
rect 401 3043 416 3077
rect 472 3043 502 3065
rect 616 3043 646 3065
rect 702 3043 717 3077
rect 795 3043 825 3070
rect 873 3104 903 3137
rect 988 3125 1018 3147
rect 1260 3125 1290 3147
rect 1840 3175 1870 3203
rect 1955 3165 1985 3187
rect 2033 3165 2063 3187
rect 2148 3175 2178 3203
rect 1375 3104 1405 3137
rect 873 3043 903 3070
rect 981 3043 996 3077
rect 1052 3043 1082 3065
rect 1196 3043 1226 3065
rect 1282 3043 1297 3077
rect 1375 3043 1405 3070
rect 1453 3104 1483 3137
rect 1568 3125 1598 3147
rect 1840 3125 1870 3147
rect 2420 3175 2450 3203
rect 2535 3165 2565 3187
rect 2613 3165 2643 3187
rect 2728 3175 2758 3203
rect 1955 3104 1985 3137
rect 1453 3043 1483 3070
rect 1561 3043 1576 3077
rect 1632 3043 1662 3065
rect 1776 3043 1806 3065
rect 1862 3043 1877 3077
rect 1955 3043 1985 3070
rect 2033 3104 2063 3137
rect 2148 3125 2178 3147
rect 2420 3125 2450 3147
rect 3000 3175 3030 3203
rect 3115 3165 3145 3187
rect 3193 3165 3223 3187
rect 3308 3175 3338 3203
rect 2535 3104 2565 3137
rect 2033 3043 2063 3070
rect 2141 3043 2156 3077
rect 2212 3043 2242 3065
rect 2356 3043 2386 3065
rect 2442 3043 2457 3077
rect 2535 3043 2565 3070
rect 2613 3104 2643 3137
rect 2728 3125 2758 3147
rect 3000 3125 3030 3147
rect 3580 3175 3610 3203
rect 3695 3165 3725 3187
rect 3773 3165 3803 3187
rect 3888 3175 3918 3203
rect 3115 3104 3145 3137
rect 2613 3043 2643 3070
rect 2721 3043 2736 3077
rect 2792 3043 2822 3065
rect 2936 3043 2966 3065
rect 3022 3043 3037 3077
rect 3115 3043 3145 3070
rect 3193 3104 3223 3137
rect 3308 3125 3338 3147
rect 3580 3125 3610 3147
rect 4160 3175 4190 3203
rect 4275 3165 4305 3187
rect 4353 3165 4383 3187
rect 4468 3175 4498 3203
rect 3695 3104 3725 3137
rect 3193 3043 3223 3070
rect 3301 3043 3316 3077
rect 3372 3043 3402 3065
rect 3516 3043 3546 3065
rect 3602 3043 3617 3077
rect 3695 3043 3725 3070
rect 3773 3104 3803 3137
rect 3888 3125 3918 3147
rect 4160 3125 4190 3147
rect 4740 3175 4770 3203
rect 4855 3165 4885 3187
rect 4933 3165 4963 3187
rect 5048 3175 5078 3203
rect 4275 3104 4305 3137
rect 3773 3043 3803 3070
rect 3881 3043 3896 3077
rect 3952 3043 3982 3065
rect 4096 3043 4126 3065
rect 4182 3043 4197 3077
rect 4275 3043 4305 3070
rect 4353 3104 4383 3137
rect 4468 3125 4498 3147
rect 4740 3125 4770 3147
rect 5320 3175 5350 3203
rect 5435 3165 5465 3187
rect 5513 3165 5543 3187
rect 5628 3175 5658 3203
rect 4855 3104 4885 3137
rect 4353 3043 4383 3070
rect 4461 3043 4476 3077
rect 4532 3043 4562 3065
rect 4676 3043 4706 3065
rect 4762 3043 4777 3077
rect 4855 3043 4885 3070
rect 4933 3104 4963 3137
rect 5048 3125 5078 3147
rect 5320 3125 5350 3147
rect 5900 3175 5930 3203
rect 6015 3165 6045 3187
rect 6093 3165 6123 3187
rect 6208 3175 6238 3203
rect 5435 3104 5465 3137
rect 4933 3043 4963 3070
rect 5041 3043 5056 3077
rect 5112 3043 5142 3065
rect 5256 3043 5286 3065
rect 5342 3043 5357 3077
rect 5435 3043 5465 3070
rect 5513 3104 5543 3137
rect 5628 3125 5658 3147
rect 5900 3125 5930 3147
rect 6480 3175 6510 3203
rect 6595 3165 6625 3187
rect 6673 3165 6703 3187
rect 6788 3175 6818 3203
rect 6015 3104 6045 3137
rect 5513 3043 5543 3070
rect 5621 3043 5636 3077
rect 5692 3043 5722 3065
rect 5836 3043 5866 3065
rect 5922 3043 5937 3077
rect 6015 3043 6045 3070
rect 6093 3104 6123 3137
rect 6208 3125 6238 3147
rect 6480 3125 6510 3147
rect 6595 3104 6625 3137
rect 6093 3043 6123 3070
rect 6201 3043 6216 3077
rect 6272 3043 6302 3065
rect 6416 3043 6446 3065
rect 6502 3043 6517 3077
rect 6595 3043 6625 3070
rect 6673 3104 6703 3137
rect 6788 3125 6818 3147
rect 6673 3043 6703 3070
rect 6781 3043 6796 3077
rect 6852 3043 6882 3065
rect 122 3029 152 3043
rect 386 3029 416 3043
rect 702 3029 732 3043
rect 966 3029 996 3043
rect 1282 3029 1312 3043
rect 1546 3029 1576 3043
rect 1862 3029 1892 3043
rect 2126 3029 2156 3043
rect 2442 3029 2472 3043
rect 2706 3029 2736 3043
rect 3022 3029 3052 3043
rect 3286 3029 3316 3043
rect 3602 3029 3632 3043
rect 3866 3029 3896 3043
rect 4182 3029 4212 3043
rect 4446 3029 4476 3043
rect 4762 3029 4792 3043
rect 5026 3029 5056 3043
rect 5342 3029 5372 3043
rect 5606 3029 5636 3043
rect 5922 3029 5952 3043
rect 6186 3029 6216 3043
rect 6502 3029 6532 3043
rect 6766 3029 6796 3043
rect 36 2979 66 3001
rect 122 2979 152 3001
rect 215 2979 245 3001
rect 293 2979 323 3001
rect 386 2979 416 3001
rect 472 2979 502 3001
rect 616 2979 646 3001
rect 702 2979 732 3001
rect 795 2979 825 3001
rect 873 2979 903 3001
rect 966 2979 996 3001
rect 1052 2979 1082 3001
rect 1196 2979 1226 3001
rect 1282 2979 1312 3001
rect 1375 2979 1405 3001
rect 1453 2979 1483 3001
rect 1546 2979 1576 3001
rect 1632 2979 1662 3001
rect 1776 2979 1806 3001
rect 1862 2979 1892 3001
rect 1955 2979 1985 3001
rect 2033 2979 2063 3001
rect 2126 2979 2156 3001
rect 2212 2979 2242 3001
rect 2356 2979 2386 3001
rect 2442 2979 2472 3001
rect 2535 2979 2565 3001
rect 2613 2979 2643 3001
rect 2706 2979 2736 3001
rect 2792 2979 2822 3001
rect 2936 2979 2966 3001
rect 3022 2979 3052 3001
rect 3115 2979 3145 3001
rect 3193 2979 3223 3001
rect 3286 2979 3316 3001
rect 3372 2979 3402 3001
rect 3516 2979 3546 3001
rect 3602 2979 3632 3001
rect 3695 2979 3725 3001
rect 3773 2979 3803 3001
rect 3866 2979 3896 3001
rect 3952 2979 3982 3001
rect 4096 2979 4126 3001
rect 4182 2979 4212 3001
rect 4275 2979 4305 3001
rect 4353 2979 4383 3001
rect 4446 2979 4476 3001
rect 4532 2979 4562 3001
rect 4676 2979 4706 3001
rect 4762 2979 4792 3001
rect 4855 2979 4885 3001
rect 4933 2979 4963 3001
rect 5026 2979 5056 3001
rect 5112 2979 5142 3001
rect 5256 2979 5286 3001
rect 5342 2979 5372 3001
rect 5435 2979 5465 3001
rect 5513 2979 5543 3001
rect 5606 2979 5636 3001
rect 5692 2979 5722 3001
rect 5836 2979 5866 3001
rect 5922 2979 5952 3001
rect 6015 2979 6045 3001
rect 6093 2979 6123 3001
rect 6186 2979 6216 3001
rect 6272 2979 6302 3001
rect 6416 2979 6446 3001
rect 6502 2979 6532 3001
rect 6595 2979 6625 3001
rect 6673 2979 6703 3001
rect 6766 2979 6796 3001
rect 6852 2979 6882 3001
rect -43 2933 6925 2963
rect 100 2905 130 2933
rect 215 2895 245 2917
rect 293 2895 323 2917
rect 408 2905 438 2933
rect 100 2855 130 2877
rect 680 2905 710 2933
rect 795 2895 825 2917
rect 873 2895 903 2917
rect 988 2905 1018 2933
rect 215 2834 245 2867
rect 36 2773 66 2795
rect 122 2773 137 2807
rect 215 2773 245 2800
rect 293 2834 323 2867
rect 408 2855 438 2877
rect 680 2855 710 2877
rect 1260 2905 1290 2933
rect 1375 2895 1405 2917
rect 1453 2895 1483 2917
rect 1568 2905 1598 2933
rect 795 2834 825 2867
rect 293 2773 323 2800
rect 401 2773 416 2807
rect 472 2773 502 2795
rect 616 2773 646 2795
rect 702 2773 717 2807
rect 795 2773 825 2800
rect 873 2834 903 2867
rect 988 2855 1018 2877
rect 1260 2855 1290 2877
rect 1840 2905 1870 2933
rect 1955 2895 1985 2917
rect 2033 2895 2063 2917
rect 2148 2905 2178 2933
rect 1375 2834 1405 2867
rect 873 2773 903 2800
rect 981 2773 996 2807
rect 1052 2773 1082 2795
rect 1196 2773 1226 2795
rect 1282 2773 1297 2807
rect 1375 2773 1405 2800
rect 1453 2834 1483 2867
rect 1568 2855 1598 2877
rect 1840 2855 1870 2877
rect 2420 2905 2450 2933
rect 2535 2895 2565 2917
rect 2613 2895 2643 2917
rect 2728 2905 2758 2933
rect 1955 2834 1985 2867
rect 1453 2773 1483 2800
rect 1561 2773 1576 2807
rect 1632 2773 1662 2795
rect 1776 2773 1806 2795
rect 1862 2773 1877 2807
rect 1955 2773 1985 2800
rect 2033 2834 2063 2867
rect 2148 2855 2178 2877
rect 2420 2855 2450 2877
rect 3000 2905 3030 2933
rect 3115 2895 3145 2917
rect 3193 2895 3223 2917
rect 3308 2905 3338 2933
rect 2535 2834 2565 2867
rect 2033 2773 2063 2800
rect 2141 2773 2156 2807
rect 2212 2773 2242 2795
rect 2356 2773 2386 2795
rect 2442 2773 2457 2807
rect 2535 2773 2565 2800
rect 2613 2834 2643 2867
rect 2728 2855 2758 2877
rect 3000 2855 3030 2877
rect 3580 2905 3610 2933
rect 3695 2895 3725 2917
rect 3773 2895 3803 2917
rect 3888 2905 3918 2933
rect 3115 2834 3145 2867
rect 2613 2773 2643 2800
rect 2721 2773 2736 2807
rect 2792 2773 2822 2795
rect 2936 2773 2966 2795
rect 3022 2773 3037 2807
rect 3115 2773 3145 2800
rect 3193 2834 3223 2867
rect 3308 2855 3338 2877
rect 3580 2855 3610 2877
rect 4160 2905 4190 2933
rect 4275 2895 4305 2917
rect 4353 2895 4383 2917
rect 4468 2905 4498 2933
rect 3695 2834 3725 2867
rect 3193 2773 3223 2800
rect 3301 2773 3316 2807
rect 3372 2773 3402 2795
rect 3516 2773 3546 2795
rect 3602 2773 3617 2807
rect 3695 2773 3725 2800
rect 3773 2834 3803 2867
rect 3888 2855 3918 2877
rect 4160 2855 4190 2877
rect 4740 2905 4770 2933
rect 4855 2895 4885 2917
rect 4933 2895 4963 2917
rect 5048 2905 5078 2933
rect 4275 2834 4305 2867
rect 3773 2773 3803 2800
rect 3881 2773 3896 2807
rect 3952 2773 3982 2795
rect 4096 2773 4126 2795
rect 4182 2773 4197 2807
rect 4275 2773 4305 2800
rect 4353 2834 4383 2867
rect 4468 2855 4498 2877
rect 4740 2855 4770 2877
rect 5320 2905 5350 2933
rect 5435 2895 5465 2917
rect 5513 2895 5543 2917
rect 5628 2905 5658 2933
rect 4855 2834 4885 2867
rect 4353 2773 4383 2800
rect 4461 2773 4476 2807
rect 4532 2773 4562 2795
rect 4676 2773 4706 2795
rect 4762 2773 4777 2807
rect 4855 2773 4885 2800
rect 4933 2834 4963 2867
rect 5048 2855 5078 2877
rect 5320 2855 5350 2877
rect 5900 2905 5930 2933
rect 6015 2895 6045 2917
rect 6093 2895 6123 2917
rect 6208 2905 6238 2933
rect 5435 2834 5465 2867
rect 4933 2773 4963 2800
rect 5041 2773 5056 2807
rect 5112 2773 5142 2795
rect 5256 2773 5286 2795
rect 5342 2773 5357 2807
rect 5435 2773 5465 2800
rect 5513 2834 5543 2867
rect 5628 2855 5658 2877
rect 5900 2855 5930 2877
rect 6480 2905 6510 2933
rect 6595 2895 6625 2917
rect 6673 2895 6703 2917
rect 6788 2905 6818 2933
rect 6015 2834 6045 2867
rect 5513 2773 5543 2800
rect 5621 2773 5636 2807
rect 5692 2773 5722 2795
rect 5836 2773 5866 2795
rect 5922 2773 5937 2807
rect 6015 2773 6045 2800
rect 6093 2834 6123 2867
rect 6208 2855 6238 2877
rect 6480 2855 6510 2877
rect 6595 2834 6625 2867
rect 6093 2773 6123 2800
rect 6201 2773 6216 2807
rect 6272 2773 6302 2795
rect 6416 2773 6446 2795
rect 6502 2773 6517 2807
rect 6595 2773 6625 2800
rect 6673 2834 6703 2867
rect 6788 2855 6818 2877
rect 6673 2773 6703 2800
rect 6781 2773 6796 2807
rect 6852 2773 6882 2795
rect 122 2759 152 2773
rect 386 2759 416 2773
rect 702 2759 732 2773
rect 966 2759 996 2773
rect 1282 2759 1312 2773
rect 1546 2759 1576 2773
rect 1862 2759 1892 2773
rect 2126 2759 2156 2773
rect 2442 2759 2472 2773
rect 2706 2759 2736 2773
rect 3022 2759 3052 2773
rect 3286 2759 3316 2773
rect 3602 2759 3632 2773
rect 3866 2759 3896 2773
rect 4182 2759 4212 2773
rect 4446 2759 4476 2773
rect 4762 2759 4792 2773
rect 5026 2759 5056 2773
rect 5342 2759 5372 2773
rect 5606 2759 5636 2773
rect 5922 2759 5952 2773
rect 6186 2759 6216 2773
rect 6502 2759 6532 2773
rect 6766 2759 6796 2773
rect 36 2709 66 2731
rect 122 2709 152 2731
rect 215 2709 245 2731
rect 293 2709 323 2731
rect 386 2709 416 2731
rect 472 2709 502 2731
rect 616 2709 646 2731
rect 702 2709 732 2731
rect 795 2709 825 2731
rect 873 2709 903 2731
rect 966 2709 996 2731
rect 1052 2709 1082 2731
rect 1196 2709 1226 2731
rect 1282 2709 1312 2731
rect 1375 2709 1405 2731
rect 1453 2709 1483 2731
rect 1546 2709 1576 2731
rect 1632 2709 1662 2731
rect 1776 2709 1806 2731
rect 1862 2709 1892 2731
rect 1955 2709 1985 2731
rect 2033 2709 2063 2731
rect 2126 2709 2156 2731
rect 2212 2709 2242 2731
rect 2356 2709 2386 2731
rect 2442 2709 2472 2731
rect 2535 2709 2565 2731
rect 2613 2709 2643 2731
rect 2706 2709 2736 2731
rect 2792 2709 2822 2731
rect 2936 2709 2966 2731
rect 3022 2709 3052 2731
rect 3115 2709 3145 2731
rect 3193 2709 3223 2731
rect 3286 2709 3316 2731
rect 3372 2709 3402 2731
rect 3516 2709 3546 2731
rect 3602 2709 3632 2731
rect 3695 2709 3725 2731
rect 3773 2709 3803 2731
rect 3866 2709 3896 2731
rect 3952 2709 3982 2731
rect 4096 2709 4126 2731
rect 4182 2709 4212 2731
rect 4275 2709 4305 2731
rect 4353 2709 4383 2731
rect 4446 2709 4476 2731
rect 4532 2709 4562 2731
rect 4676 2709 4706 2731
rect 4762 2709 4792 2731
rect 4855 2709 4885 2731
rect 4933 2709 4963 2731
rect 5026 2709 5056 2731
rect 5112 2709 5142 2731
rect 5256 2709 5286 2731
rect 5342 2709 5372 2731
rect 5435 2709 5465 2731
rect 5513 2709 5543 2731
rect 5606 2709 5636 2731
rect 5692 2709 5722 2731
rect 5836 2709 5866 2731
rect 5922 2709 5952 2731
rect 6015 2709 6045 2731
rect 6093 2709 6123 2731
rect 6186 2709 6216 2731
rect 6272 2709 6302 2731
rect 6416 2709 6446 2731
rect 6502 2709 6532 2731
rect 6595 2709 6625 2731
rect 6673 2709 6703 2731
rect 6766 2709 6796 2731
rect 6852 2709 6882 2731
rect -43 2663 6925 2693
rect 100 2635 130 2663
rect 215 2625 245 2647
rect 293 2625 323 2647
rect 408 2635 438 2663
rect 100 2585 130 2607
rect 680 2635 710 2663
rect 795 2625 825 2647
rect 873 2625 903 2647
rect 988 2635 1018 2663
rect 215 2564 245 2597
rect 36 2503 66 2525
rect 122 2503 137 2537
rect 215 2503 245 2530
rect 293 2564 323 2597
rect 408 2585 438 2607
rect 680 2585 710 2607
rect 1260 2635 1290 2663
rect 1375 2625 1405 2647
rect 1453 2625 1483 2647
rect 1568 2635 1598 2663
rect 795 2564 825 2597
rect 293 2503 323 2530
rect 401 2503 416 2537
rect 472 2503 502 2525
rect 616 2503 646 2525
rect 702 2503 717 2537
rect 795 2503 825 2530
rect 873 2564 903 2597
rect 988 2585 1018 2607
rect 1260 2585 1290 2607
rect 1840 2635 1870 2663
rect 1955 2625 1985 2647
rect 2033 2625 2063 2647
rect 2148 2635 2178 2663
rect 1375 2564 1405 2597
rect 873 2503 903 2530
rect 981 2503 996 2537
rect 1052 2503 1082 2525
rect 1196 2503 1226 2525
rect 1282 2503 1297 2537
rect 1375 2503 1405 2530
rect 1453 2564 1483 2597
rect 1568 2585 1598 2607
rect 1840 2585 1870 2607
rect 2420 2635 2450 2663
rect 2535 2625 2565 2647
rect 2613 2625 2643 2647
rect 2728 2635 2758 2663
rect 1955 2564 1985 2597
rect 1453 2503 1483 2530
rect 1561 2503 1576 2537
rect 1632 2503 1662 2525
rect 1776 2503 1806 2525
rect 1862 2503 1877 2537
rect 1955 2503 1985 2530
rect 2033 2564 2063 2597
rect 2148 2585 2178 2607
rect 2420 2585 2450 2607
rect 3000 2635 3030 2663
rect 3115 2625 3145 2647
rect 3193 2625 3223 2647
rect 3308 2635 3338 2663
rect 2535 2564 2565 2597
rect 2033 2503 2063 2530
rect 2141 2503 2156 2537
rect 2212 2503 2242 2525
rect 2356 2503 2386 2525
rect 2442 2503 2457 2537
rect 2535 2503 2565 2530
rect 2613 2564 2643 2597
rect 2728 2585 2758 2607
rect 3000 2585 3030 2607
rect 3580 2635 3610 2663
rect 3695 2625 3725 2647
rect 3773 2625 3803 2647
rect 3888 2635 3918 2663
rect 3115 2564 3145 2597
rect 2613 2503 2643 2530
rect 2721 2503 2736 2537
rect 2792 2503 2822 2525
rect 2936 2503 2966 2525
rect 3022 2503 3037 2537
rect 3115 2503 3145 2530
rect 3193 2564 3223 2597
rect 3308 2585 3338 2607
rect 3580 2585 3610 2607
rect 4160 2635 4190 2663
rect 4275 2625 4305 2647
rect 4353 2625 4383 2647
rect 4468 2635 4498 2663
rect 3695 2564 3725 2597
rect 3193 2503 3223 2530
rect 3301 2503 3316 2537
rect 3372 2503 3402 2525
rect 3516 2503 3546 2525
rect 3602 2503 3617 2537
rect 3695 2503 3725 2530
rect 3773 2564 3803 2597
rect 3888 2585 3918 2607
rect 4160 2585 4190 2607
rect 4740 2635 4770 2663
rect 4855 2625 4885 2647
rect 4933 2625 4963 2647
rect 5048 2635 5078 2663
rect 4275 2564 4305 2597
rect 3773 2503 3803 2530
rect 3881 2503 3896 2537
rect 3952 2503 3982 2525
rect 4096 2503 4126 2525
rect 4182 2503 4197 2537
rect 4275 2503 4305 2530
rect 4353 2564 4383 2597
rect 4468 2585 4498 2607
rect 4740 2585 4770 2607
rect 5320 2635 5350 2663
rect 5435 2625 5465 2647
rect 5513 2625 5543 2647
rect 5628 2635 5658 2663
rect 4855 2564 4885 2597
rect 4353 2503 4383 2530
rect 4461 2503 4476 2537
rect 4532 2503 4562 2525
rect 4676 2503 4706 2525
rect 4762 2503 4777 2537
rect 4855 2503 4885 2530
rect 4933 2564 4963 2597
rect 5048 2585 5078 2607
rect 5320 2585 5350 2607
rect 5900 2635 5930 2663
rect 6015 2625 6045 2647
rect 6093 2625 6123 2647
rect 6208 2635 6238 2663
rect 5435 2564 5465 2597
rect 4933 2503 4963 2530
rect 5041 2503 5056 2537
rect 5112 2503 5142 2525
rect 5256 2503 5286 2525
rect 5342 2503 5357 2537
rect 5435 2503 5465 2530
rect 5513 2564 5543 2597
rect 5628 2585 5658 2607
rect 5900 2585 5930 2607
rect 6480 2635 6510 2663
rect 6595 2625 6625 2647
rect 6673 2625 6703 2647
rect 6788 2635 6818 2663
rect 6015 2564 6045 2597
rect 5513 2503 5543 2530
rect 5621 2503 5636 2537
rect 5692 2503 5722 2525
rect 5836 2503 5866 2525
rect 5922 2503 5937 2537
rect 6015 2503 6045 2530
rect 6093 2564 6123 2597
rect 6208 2585 6238 2607
rect 6480 2585 6510 2607
rect 6595 2564 6625 2597
rect 6093 2503 6123 2530
rect 6201 2503 6216 2537
rect 6272 2503 6302 2525
rect 6416 2503 6446 2525
rect 6502 2503 6517 2537
rect 6595 2503 6625 2530
rect 6673 2564 6703 2597
rect 6788 2585 6818 2607
rect 6673 2503 6703 2530
rect 6781 2503 6796 2537
rect 6852 2503 6882 2525
rect 122 2489 152 2503
rect 386 2489 416 2503
rect 702 2489 732 2503
rect 966 2489 996 2503
rect 1282 2489 1312 2503
rect 1546 2489 1576 2503
rect 1862 2489 1892 2503
rect 2126 2489 2156 2503
rect 2442 2489 2472 2503
rect 2706 2489 2736 2503
rect 3022 2489 3052 2503
rect 3286 2489 3316 2503
rect 3602 2489 3632 2503
rect 3866 2489 3896 2503
rect 4182 2489 4212 2503
rect 4446 2489 4476 2503
rect 4762 2489 4792 2503
rect 5026 2489 5056 2503
rect 5342 2489 5372 2503
rect 5606 2489 5636 2503
rect 5922 2489 5952 2503
rect 6186 2489 6216 2503
rect 6502 2489 6532 2503
rect 6766 2489 6796 2503
rect 36 2439 66 2461
rect 122 2439 152 2461
rect 215 2439 245 2461
rect 293 2439 323 2461
rect 386 2439 416 2461
rect 472 2439 502 2461
rect 616 2439 646 2461
rect 702 2439 732 2461
rect 795 2439 825 2461
rect 873 2439 903 2461
rect 966 2439 996 2461
rect 1052 2439 1082 2461
rect 1196 2439 1226 2461
rect 1282 2439 1312 2461
rect 1375 2439 1405 2461
rect 1453 2439 1483 2461
rect 1546 2439 1576 2461
rect 1632 2439 1662 2461
rect 1776 2439 1806 2461
rect 1862 2439 1892 2461
rect 1955 2439 1985 2461
rect 2033 2439 2063 2461
rect 2126 2439 2156 2461
rect 2212 2439 2242 2461
rect 2356 2439 2386 2461
rect 2442 2439 2472 2461
rect 2535 2439 2565 2461
rect 2613 2439 2643 2461
rect 2706 2439 2736 2461
rect 2792 2439 2822 2461
rect 2936 2439 2966 2461
rect 3022 2439 3052 2461
rect 3115 2439 3145 2461
rect 3193 2439 3223 2461
rect 3286 2439 3316 2461
rect 3372 2439 3402 2461
rect 3516 2439 3546 2461
rect 3602 2439 3632 2461
rect 3695 2439 3725 2461
rect 3773 2439 3803 2461
rect 3866 2439 3896 2461
rect 3952 2439 3982 2461
rect 4096 2439 4126 2461
rect 4182 2439 4212 2461
rect 4275 2439 4305 2461
rect 4353 2439 4383 2461
rect 4446 2439 4476 2461
rect 4532 2439 4562 2461
rect 4676 2439 4706 2461
rect 4762 2439 4792 2461
rect 4855 2439 4885 2461
rect 4933 2439 4963 2461
rect 5026 2439 5056 2461
rect 5112 2439 5142 2461
rect 5256 2439 5286 2461
rect 5342 2439 5372 2461
rect 5435 2439 5465 2461
rect 5513 2439 5543 2461
rect 5606 2439 5636 2461
rect 5692 2439 5722 2461
rect 5836 2439 5866 2461
rect 5922 2439 5952 2461
rect 6015 2439 6045 2461
rect 6093 2439 6123 2461
rect 6186 2439 6216 2461
rect 6272 2439 6302 2461
rect 6416 2439 6446 2461
rect 6502 2439 6532 2461
rect 6595 2439 6625 2461
rect 6673 2439 6703 2461
rect 6766 2439 6796 2461
rect 6852 2439 6882 2461
rect -43 2393 6925 2423
rect 100 2365 130 2393
rect 215 2355 245 2377
rect 293 2355 323 2377
rect 408 2365 438 2393
rect 100 2315 130 2337
rect 680 2365 710 2393
rect 795 2355 825 2377
rect 873 2355 903 2377
rect 988 2365 1018 2393
rect 215 2294 245 2327
rect 36 2233 66 2255
rect 122 2233 137 2267
rect 215 2233 245 2260
rect 293 2294 323 2327
rect 408 2315 438 2337
rect 680 2315 710 2337
rect 1260 2365 1290 2393
rect 1375 2355 1405 2377
rect 1453 2355 1483 2377
rect 1568 2365 1598 2393
rect 795 2294 825 2327
rect 293 2233 323 2260
rect 401 2233 416 2267
rect 472 2233 502 2255
rect 616 2233 646 2255
rect 702 2233 717 2267
rect 795 2233 825 2260
rect 873 2294 903 2327
rect 988 2315 1018 2337
rect 1260 2315 1290 2337
rect 1840 2365 1870 2393
rect 1955 2355 1985 2377
rect 2033 2355 2063 2377
rect 2148 2365 2178 2393
rect 1375 2294 1405 2327
rect 873 2233 903 2260
rect 981 2233 996 2267
rect 1052 2233 1082 2255
rect 1196 2233 1226 2255
rect 1282 2233 1297 2267
rect 1375 2233 1405 2260
rect 1453 2294 1483 2327
rect 1568 2315 1598 2337
rect 1840 2315 1870 2337
rect 2420 2365 2450 2393
rect 2535 2355 2565 2377
rect 2613 2355 2643 2377
rect 2728 2365 2758 2393
rect 1955 2294 1985 2327
rect 1453 2233 1483 2260
rect 1561 2233 1576 2267
rect 1632 2233 1662 2255
rect 1776 2233 1806 2255
rect 1862 2233 1877 2267
rect 1955 2233 1985 2260
rect 2033 2294 2063 2327
rect 2148 2315 2178 2337
rect 2420 2315 2450 2337
rect 3000 2365 3030 2393
rect 3115 2355 3145 2377
rect 3193 2355 3223 2377
rect 3308 2365 3338 2393
rect 2535 2294 2565 2327
rect 2033 2233 2063 2260
rect 2141 2233 2156 2267
rect 2212 2233 2242 2255
rect 2356 2233 2386 2255
rect 2442 2233 2457 2267
rect 2535 2233 2565 2260
rect 2613 2294 2643 2327
rect 2728 2315 2758 2337
rect 3000 2315 3030 2337
rect 3580 2365 3610 2393
rect 3695 2355 3725 2377
rect 3773 2355 3803 2377
rect 3888 2365 3918 2393
rect 3115 2294 3145 2327
rect 2613 2233 2643 2260
rect 2721 2233 2736 2267
rect 2792 2233 2822 2255
rect 2936 2233 2966 2255
rect 3022 2233 3037 2267
rect 3115 2233 3145 2260
rect 3193 2294 3223 2327
rect 3308 2315 3338 2337
rect 3580 2315 3610 2337
rect 4160 2365 4190 2393
rect 4275 2355 4305 2377
rect 4353 2355 4383 2377
rect 4468 2365 4498 2393
rect 3695 2294 3725 2327
rect 3193 2233 3223 2260
rect 3301 2233 3316 2267
rect 3372 2233 3402 2255
rect 3516 2233 3546 2255
rect 3602 2233 3617 2267
rect 3695 2233 3725 2260
rect 3773 2294 3803 2327
rect 3888 2315 3918 2337
rect 4160 2315 4190 2337
rect 4740 2365 4770 2393
rect 4855 2355 4885 2377
rect 4933 2355 4963 2377
rect 5048 2365 5078 2393
rect 4275 2294 4305 2327
rect 3773 2233 3803 2260
rect 3881 2233 3896 2267
rect 3952 2233 3982 2255
rect 4096 2233 4126 2255
rect 4182 2233 4197 2267
rect 4275 2233 4305 2260
rect 4353 2294 4383 2327
rect 4468 2315 4498 2337
rect 4740 2315 4770 2337
rect 5320 2365 5350 2393
rect 5435 2355 5465 2377
rect 5513 2355 5543 2377
rect 5628 2365 5658 2393
rect 4855 2294 4885 2327
rect 4353 2233 4383 2260
rect 4461 2233 4476 2267
rect 4532 2233 4562 2255
rect 4676 2233 4706 2255
rect 4762 2233 4777 2267
rect 4855 2233 4885 2260
rect 4933 2294 4963 2327
rect 5048 2315 5078 2337
rect 5320 2315 5350 2337
rect 5900 2365 5930 2393
rect 6015 2355 6045 2377
rect 6093 2355 6123 2377
rect 6208 2365 6238 2393
rect 5435 2294 5465 2327
rect 4933 2233 4963 2260
rect 5041 2233 5056 2267
rect 5112 2233 5142 2255
rect 5256 2233 5286 2255
rect 5342 2233 5357 2267
rect 5435 2233 5465 2260
rect 5513 2294 5543 2327
rect 5628 2315 5658 2337
rect 5900 2315 5930 2337
rect 6480 2365 6510 2393
rect 6595 2355 6625 2377
rect 6673 2355 6703 2377
rect 6788 2365 6818 2393
rect 6015 2294 6045 2327
rect 5513 2233 5543 2260
rect 5621 2233 5636 2267
rect 5692 2233 5722 2255
rect 5836 2233 5866 2255
rect 5922 2233 5937 2267
rect 6015 2233 6045 2260
rect 6093 2294 6123 2327
rect 6208 2315 6238 2337
rect 6480 2315 6510 2337
rect 6595 2294 6625 2327
rect 6093 2233 6123 2260
rect 6201 2233 6216 2267
rect 6272 2233 6302 2255
rect 6416 2233 6446 2255
rect 6502 2233 6517 2267
rect 6595 2233 6625 2260
rect 6673 2294 6703 2327
rect 6788 2315 6818 2337
rect 6673 2233 6703 2260
rect 6781 2233 6796 2267
rect 6852 2233 6882 2255
rect 122 2219 152 2233
rect 386 2219 416 2233
rect 702 2219 732 2233
rect 966 2219 996 2233
rect 1282 2219 1312 2233
rect 1546 2219 1576 2233
rect 1862 2219 1892 2233
rect 2126 2219 2156 2233
rect 2442 2219 2472 2233
rect 2706 2219 2736 2233
rect 3022 2219 3052 2233
rect 3286 2219 3316 2233
rect 3602 2219 3632 2233
rect 3866 2219 3896 2233
rect 4182 2219 4212 2233
rect 4446 2219 4476 2233
rect 4762 2219 4792 2233
rect 5026 2219 5056 2233
rect 5342 2219 5372 2233
rect 5606 2219 5636 2233
rect 5922 2219 5952 2233
rect 6186 2219 6216 2233
rect 6502 2219 6532 2233
rect 6766 2219 6796 2233
rect 36 2169 66 2191
rect 122 2169 152 2191
rect 215 2169 245 2191
rect 293 2169 323 2191
rect 386 2169 416 2191
rect 472 2169 502 2191
rect 616 2169 646 2191
rect 702 2169 732 2191
rect 795 2169 825 2191
rect 873 2169 903 2191
rect 966 2169 996 2191
rect 1052 2169 1082 2191
rect 1196 2169 1226 2191
rect 1282 2169 1312 2191
rect 1375 2169 1405 2191
rect 1453 2169 1483 2191
rect 1546 2169 1576 2191
rect 1632 2169 1662 2191
rect 1776 2169 1806 2191
rect 1862 2169 1892 2191
rect 1955 2169 1985 2191
rect 2033 2169 2063 2191
rect 2126 2169 2156 2191
rect 2212 2169 2242 2191
rect 2356 2169 2386 2191
rect 2442 2169 2472 2191
rect 2535 2169 2565 2191
rect 2613 2169 2643 2191
rect 2706 2169 2736 2191
rect 2792 2169 2822 2191
rect 2936 2169 2966 2191
rect 3022 2169 3052 2191
rect 3115 2169 3145 2191
rect 3193 2169 3223 2191
rect 3286 2169 3316 2191
rect 3372 2169 3402 2191
rect 3516 2169 3546 2191
rect 3602 2169 3632 2191
rect 3695 2169 3725 2191
rect 3773 2169 3803 2191
rect 3866 2169 3896 2191
rect 3952 2169 3982 2191
rect 4096 2169 4126 2191
rect 4182 2169 4212 2191
rect 4275 2169 4305 2191
rect 4353 2169 4383 2191
rect 4446 2169 4476 2191
rect 4532 2169 4562 2191
rect 4676 2169 4706 2191
rect 4762 2169 4792 2191
rect 4855 2169 4885 2191
rect 4933 2169 4963 2191
rect 5026 2169 5056 2191
rect 5112 2169 5142 2191
rect 5256 2169 5286 2191
rect 5342 2169 5372 2191
rect 5435 2169 5465 2191
rect 5513 2169 5543 2191
rect 5606 2169 5636 2191
rect 5692 2169 5722 2191
rect 5836 2169 5866 2191
rect 5922 2169 5952 2191
rect 6015 2169 6045 2191
rect 6093 2169 6123 2191
rect 6186 2169 6216 2191
rect 6272 2169 6302 2191
rect 6416 2169 6446 2191
rect 6502 2169 6532 2191
rect 6595 2169 6625 2191
rect 6673 2169 6703 2191
rect 6766 2169 6796 2191
rect 6852 2169 6882 2191
rect -43 2123 6925 2153
rect 100 2095 130 2123
rect 215 2085 245 2107
rect 293 2085 323 2107
rect 408 2095 438 2123
rect 100 2045 130 2067
rect 680 2095 710 2123
rect 795 2085 825 2107
rect 873 2085 903 2107
rect 988 2095 1018 2123
rect 215 2024 245 2057
rect 36 1963 66 1985
rect 122 1963 137 1997
rect 215 1963 245 1990
rect 293 2024 323 2057
rect 408 2045 438 2067
rect 680 2045 710 2067
rect 1260 2095 1290 2123
rect 1375 2085 1405 2107
rect 1453 2085 1483 2107
rect 1568 2095 1598 2123
rect 795 2024 825 2057
rect 293 1963 323 1990
rect 401 1963 416 1997
rect 472 1963 502 1985
rect 616 1963 646 1985
rect 702 1963 717 1997
rect 795 1963 825 1990
rect 873 2024 903 2057
rect 988 2045 1018 2067
rect 1260 2045 1290 2067
rect 1840 2095 1870 2123
rect 1955 2085 1985 2107
rect 2033 2085 2063 2107
rect 2148 2095 2178 2123
rect 1375 2024 1405 2057
rect 873 1963 903 1990
rect 981 1963 996 1997
rect 1052 1963 1082 1985
rect 1196 1963 1226 1985
rect 1282 1963 1297 1997
rect 1375 1963 1405 1990
rect 1453 2024 1483 2057
rect 1568 2045 1598 2067
rect 1840 2045 1870 2067
rect 2420 2095 2450 2123
rect 2535 2085 2565 2107
rect 2613 2085 2643 2107
rect 2728 2095 2758 2123
rect 1955 2024 1985 2057
rect 1453 1963 1483 1990
rect 1561 1963 1576 1997
rect 1632 1963 1662 1985
rect 1776 1963 1806 1985
rect 1862 1963 1877 1997
rect 1955 1963 1985 1990
rect 2033 2024 2063 2057
rect 2148 2045 2178 2067
rect 2420 2045 2450 2067
rect 3000 2095 3030 2123
rect 3115 2085 3145 2107
rect 3193 2085 3223 2107
rect 3308 2095 3338 2123
rect 2535 2024 2565 2057
rect 2033 1963 2063 1990
rect 2141 1963 2156 1997
rect 2212 1963 2242 1985
rect 2356 1963 2386 1985
rect 2442 1963 2457 1997
rect 2535 1963 2565 1990
rect 2613 2024 2643 2057
rect 2728 2045 2758 2067
rect 3000 2045 3030 2067
rect 3580 2095 3610 2123
rect 3695 2085 3725 2107
rect 3773 2085 3803 2107
rect 3888 2095 3918 2123
rect 3115 2024 3145 2057
rect 2613 1963 2643 1990
rect 2721 1963 2736 1997
rect 2792 1963 2822 1985
rect 2936 1963 2966 1985
rect 3022 1963 3037 1997
rect 3115 1963 3145 1990
rect 3193 2024 3223 2057
rect 3308 2045 3338 2067
rect 3580 2045 3610 2067
rect 4160 2095 4190 2123
rect 4275 2085 4305 2107
rect 4353 2085 4383 2107
rect 4468 2095 4498 2123
rect 3695 2024 3725 2057
rect 3193 1963 3223 1990
rect 3301 1963 3316 1997
rect 3372 1963 3402 1985
rect 3516 1963 3546 1985
rect 3602 1963 3617 1997
rect 3695 1963 3725 1990
rect 3773 2024 3803 2057
rect 3888 2045 3918 2067
rect 4160 2045 4190 2067
rect 4740 2095 4770 2123
rect 4855 2085 4885 2107
rect 4933 2085 4963 2107
rect 5048 2095 5078 2123
rect 4275 2024 4305 2057
rect 3773 1963 3803 1990
rect 3881 1963 3896 1997
rect 3952 1963 3982 1985
rect 4096 1963 4126 1985
rect 4182 1963 4197 1997
rect 4275 1963 4305 1990
rect 4353 2024 4383 2057
rect 4468 2045 4498 2067
rect 4740 2045 4770 2067
rect 5320 2095 5350 2123
rect 5435 2085 5465 2107
rect 5513 2085 5543 2107
rect 5628 2095 5658 2123
rect 4855 2024 4885 2057
rect 4353 1963 4383 1990
rect 4461 1963 4476 1997
rect 4532 1963 4562 1985
rect 4676 1963 4706 1985
rect 4762 1963 4777 1997
rect 4855 1963 4885 1990
rect 4933 2024 4963 2057
rect 5048 2045 5078 2067
rect 5320 2045 5350 2067
rect 5900 2095 5930 2123
rect 6015 2085 6045 2107
rect 6093 2085 6123 2107
rect 6208 2095 6238 2123
rect 5435 2024 5465 2057
rect 4933 1963 4963 1990
rect 5041 1963 5056 1997
rect 5112 1963 5142 1985
rect 5256 1963 5286 1985
rect 5342 1963 5357 1997
rect 5435 1963 5465 1990
rect 5513 2024 5543 2057
rect 5628 2045 5658 2067
rect 5900 2045 5930 2067
rect 6480 2095 6510 2123
rect 6595 2085 6625 2107
rect 6673 2085 6703 2107
rect 6788 2095 6818 2123
rect 6015 2024 6045 2057
rect 5513 1963 5543 1990
rect 5621 1963 5636 1997
rect 5692 1963 5722 1985
rect 5836 1963 5866 1985
rect 5922 1963 5937 1997
rect 6015 1963 6045 1990
rect 6093 2024 6123 2057
rect 6208 2045 6238 2067
rect 6480 2045 6510 2067
rect 6595 2024 6625 2057
rect 6093 1963 6123 1990
rect 6201 1963 6216 1997
rect 6272 1963 6302 1985
rect 6416 1963 6446 1985
rect 6502 1963 6517 1997
rect 6595 1963 6625 1990
rect 6673 2024 6703 2057
rect 6788 2045 6818 2067
rect 6673 1963 6703 1990
rect 6781 1963 6796 1997
rect 6852 1963 6882 1985
rect 122 1949 152 1963
rect 386 1949 416 1963
rect 702 1949 732 1963
rect 966 1949 996 1963
rect 1282 1949 1312 1963
rect 1546 1949 1576 1963
rect 1862 1949 1892 1963
rect 2126 1949 2156 1963
rect 2442 1949 2472 1963
rect 2706 1949 2736 1963
rect 3022 1949 3052 1963
rect 3286 1949 3316 1963
rect 3602 1949 3632 1963
rect 3866 1949 3896 1963
rect 4182 1949 4212 1963
rect 4446 1949 4476 1963
rect 4762 1949 4792 1963
rect 5026 1949 5056 1963
rect 5342 1949 5372 1963
rect 5606 1949 5636 1963
rect 5922 1949 5952 1963
rect 6186 1949 6216 1963
rect 6502 1949 6532 1963
rect 6766 1949 6796 1963
rect 36 1899 66 1921
rect 122 1899 152 1921
rect 215 1899 245 1921
rect 293 1899 323 1921
rect 386 1899 416 1921
rect 472 1899 502 1921
rect 616 1899 646 1921
rect 702 1899 732 1921
rect 795 1899 825 1921
rect 873 1899 903 1921
rect 966 1899 996 1921
rect 1052 1899 1082 1921
rect 1196 1899 1226 1921
rect 1282 1899 1312 1921
rect 1375 1899 1405 1921
rect 1453 1899 1483 1921
rect 1546 1899 1576 1921
rect 1632 1899 1662 1921
rect 1776 1899 1806 1921
rect 1862 1899 1892 1921
rect 1955 1899 1985 1921
rect 2033 1899 2063 1921
rect 2126 1899 2156 1921
rect 2212 1899 2242 1921
rect 2356 1899 2386 1921
rect 2442 1899 2472 1921
rect 2535 1899 2565 1921
rect 2613 1899 2643 1921
rect 2706 1899 2736 1921
rect 2792 1899 2822 1921
rect 2936 1899 2966 1921
rect 3022 1899 3052 1921
rect 3115 1899 3145 1921
rect 3193 1899 3223 1921
rect 3286 1899 3316 1921
rect 3372 1899 3402 1921
rect 3516 1899 3546 1921
rect 3602 1899 3632 1921
rect 3695 1899 3725 1921
rect 3773 1899 3803 1921
rect 3866 1899 3896 1921
rect 3952 1899 3982 1921
rect 4096 1899 4126 1921
rect 4182 1899 4212 1921
rect 4275 1899 4305 1921
rect 4353 1899 4383 1921
rect 4446 1899 4476 1921
rect 4532 1899 4562 1921
rect 4676 1899 4706 1921
rect 4762 1899 4792 1921
rect 4855 1899 4885 1921
rect 4933 1899 4963 1921
rect 5026 1899 5056 1921
rect 5112 1899 5142 1921
rect 5256 1899 5286 1921
rect 5342 1899 5372 1921
rect 5435 1899 5465 1921
rect 5513 1899 5543 1921
rect 5606 1899 5636 1921
rect 5692 1899 5722 1921
rect 5836 1899 5866 1921
rect 5922 1899 5952 1921
rect 6015 1899 6045 1921
rect 6093 1899 6123 1921
rect 6186 1899 6216 1921
rect 6272 1899 6302 1921
rect 6416 1899 6446 1921
rect 6502 1899 6532 1921
rect 6595 1899 6625 1921
rect 6673 1899 6703 1921
rect 6766 1899 6796 1921
rect 6852 1899 6882 1921
rect -43 1853 6925 1883
rect 100 1825 130 1853
rect 215 1815 245 1837
rect 293 1815 323 1837
rect 408 1825 438 1853
rect 100 1775 130 1797
rect 680 1825 710 1853
rect 795 1815 825 1837
rect 873 1815 903 1837
rect 988 1825 1018 1853
rect 215 1754 245 1787
rect 36 1693 66 1715
rect 122 1693 137 1727
rect 215 1693 245 1720
rect 293 1754 323 1787
rect 408 1775 438 1797
rect 680 1775 710 1797
rect 1260 1825 1290 1853
rect 1375 1815 1405 1837
rect 1453 1815 1483 1837
rect 1568 1825 1598 1853
rect 795 1754 825 1787
rect 293 1693 323 1720
rect 401 1693 416 1727
rect 472 1693 502 1715
rect 616 1693 646 1715
rect 702 1693 717 1727
rect 795 1693 825 1720
rect 873 1754 903 1787
rect 988 1775 1018 1797
rect 1260 1775 1290 1797
rect 1840 1825 1870 1853
rect 1955 1815 1985 1837
rect 2033 1815 2063 1837
rect 2148 1825 2178 1853
rect 1375 1754 1405 1787
rect 873 1693 903 1720
rect 981 1693 996 1727
rect 1052 1693 1082 1715
rect 1196 1693 1226 1715
rect 1282 1693 1297 1727
rect 1375 1693 1405 1720
rect 1453 1754 1483 1787
rect 1568 1775 1598 1797
rect 1840 1775 1870 1797
rect 2420 1825 2450 1853
rect 2535 1815 2565 1837
rect 2613 1815 2643 1837
rect 2728 1825 2758 1853
rect 1955 1754 1985 1787
rect 1453 1693 1483 1720
rect 1561 1693 1576 1727
rect 1632 1693 1662 1715
rect 1776 1693 1806 1715
rect 1862 1693 1877 1727
rect 1955 1693 1985 1720
rect 2033 1754 2063 1787
rect 2148 1775 2178 1797
rect 2420 1775 2450 1797
rect 3000 1825 3030 1853
rect 3115 1815 3145 1837
rect 3193 1815 3223 1837
rect 3308 1825 3338 1853
rect 2535 1754 2565 1787
rect 2033 1693 2063 1720
rect 2141 1693 2156 1727
rect 2212 1693 2242 1715
rect 2356 1693 2386 1715
rect 2442 1693 2457 1727
rect 2535 1693 2565 1720
rect 2613 1754 2643 1787
rect 2728 1775 2758 1797
rect 3000 1775 3030 1797
rect 3580 1825 3610 1853
rect 3695 1815 3725 1837
rect 3773 1815 3803 1837
rect 3888 1825 3918 1853
rect 3115 1754 3145 1787
rect 2613 1693 2643 1720
rect 2721 1693 2736 1727
rect 2792 1693 2822 1715
rect 2936 1693 2966 1715
rect 3022 1693 3037 1727
rect 3115 1693 3145 1720
rect 3193 1754 3223 1787
rect 3308 1775 3338 1797
rect 3580 1775 3610 1797
rect 4160 1825 4190 1853
rect 4275 1815 4305 1837
rect 4353 1815 4383 1837
rect 4468 1825 4498 1853
rect 3695 1754 3725 1787
rect 3193 1693 3223 1720
rect 3301 1693 3316 1727
rect 3372 1693 3402 1715
rect 3516 1693 3546 1715
rect 3602 1693 3617 1727
rect 3695 1693 3725 1720
rect 3773 1754 3803 1787
rect 3888 1775 3918 1797
rect 4160 1775 4190 1797
rect 4740 1825 4770 1853
rect 4855 1815 4885 1837
rect 4933 1815 4963 1837
rect 5048 1825 5078 1853
rect 4275 1754 4305 1787
rect 3773 1693 3803 1720
rect 3881 1693 3896 1727
rect 3952 1693 3982 1715
rect 4096 1693 4126 1715
rect 4182 1693 4197 1727
rect 4275 1693 4305 1720
rect 4353 1754 4383 1787
rect 4468 1775 4498 1797
rect 4740 1775 4770 1797
rect 5320 1825 5350 1853
rect 5435 1815 5465 1837
rect 5513 1815 5543 1837
rect 5628 1825 5658 1853
rect 4855 1754 4885 1787
rect 4353 1693 4383 1720
rect 4461 1693 4476 1727
rect 4532 1693 4562 1715
rect 4676 1693 4706 1715
rect 4762 1693 4777 1727
rect 4855 1693 4885 1720
rect 4933 1754 4963 1787
rect 5048 1775 5078 1797
rect 5320 1775 5350 1797
rect 5900 1825 5930 1853
rect 6015 1815 6045 1837
rect 6093 1815 6123 1837
rect 6208 1825 6238 1853
rect 5435 1754 5465 1787
rect 4933 1693 4963 1720
rect 5041 1693 5056 1727
rect 5112 1693 5142 1715
rect 5256 1693 5286 1715
rect 5342 1693 5357 1727
rect 5435 1693 5465 1720
rect 5513 1754 5543 1787
rect 5628 1775 5658 1797
rect 5900 1775 5930 1797
rect 6480 1825 6510 1853
rect 6595 1815 6625 1837
rect 6673 1815 6703 1837
rect 6788 1825 6818 1853
rect 6015 1754 6045 1787
rect 5513 1693 5543 1720
rect 5621 1693 5636 1727
rect 5692 1693 5722 1715
rect 5836 1693 5866 1715
rect 5922 1693 5937 1727
rect 6015 1693 6045 1720
rect 6093 1754 6123 1787
rect 6208 1775 6238 1797
rect 6480 1775 6510 1797
rect 6595 1754 6625 1787
rect 6093 1693 6123 1720
rect 6201 1693 6216 1727
rect 6272 1693 6302 1715
rect 6416 1693 6446 1715
rect 6502 1693 6517 1727
rect 6595 1693 6625 1720
rect 6673 1754 6703 1787
rect 6788 1775 6818 1797
rect 6673 1693 6703 1720
rect 6781 1693 6796 1727
rect 6852 1693 6882 1715
rect 122 1679 152 1693
rect 386 1679 416 1693
rect 702 1679 732 1693
rect 966 1679 996 1693
rect 1282 1679 1312 1693
rect 1546 1679 1576 1693
rect 1862 1679 1892 1693
rect 2126 1679 2156 1693
rect 2442 1679 2472 1693
rect 2706 1679 2736 1693
rect 3022 1679 3052 1693
rect 3286 1679 3316 1693
rect 3602 1679 3632 1693
rect 3866 1679 3896 1693
rect 4182 1679 4212 1693
rect 4446 1679 4476 1693
rect 4762 1679 4792 1693
rect 5026 1679 5056 1693
rect 5342 1679 5372 1693
rect 5606 1679 5636 1693
rect 5922 1679 5952 1693
rect 6186 1679 6216 1693
rect 6502 1679 6532 1693
rect 6766 1679 6796 1693
rect 36 1629 66 1651
rect 122 1629 152 1651
rect 215 1629 245 1651
rect 293 1629 323 1651
rect 386 1629 416 1651
rect 472 1629 502 1651
rect 616 1629 646 1651
rect 702 1629 732 1651
rect 795 1629 825 1651
rect 873 1629 903 1651
rect 966 1629 996 1651
rect 1052 1629 1082 1651
rect 1196 1629 1226 1651
rect 1282 1629 1312 1651
rect 1375 1629 1405 1651
rect 1453 1629 1483 1651
rect 1546 1629 1576 1651
rect 1632 1629 1662 1651
rect 1776 1629 1806 1651
rect 1862 1629 1892 1651
rect 1955 1629 1985 1651
rect 2033 1629 2063 1651
rect 2126 1629 2156 1651
rect 2212 1629 2242 1651
rect 2356 1629 2386 1651
rect 2442 1629 2472 1651
rect 2535 1629 2565 1651
rect 2613 1629 2643 1651
rect 2706 1629 2736 1651
rect 2792 1629 2822 1651
rect 2936 1629 2966 1651
rect 3022 1629 3052 1651
rect 3115 1629 3145 1651
rect 3193 1629 3223 1651
rect 3286 1629 3316 1651
rect 3372 1629 3402 1651
rect 3516 1629 3546 1651
rect 3602 1629 3632 1651
rect 3695 1629 3725 1651
rect 3773 1629 3803 1651
rect 3866 1629 3896 1651
rect 3952 1629 3982 1651
rect 4096 1629 4126 1651
rect 4182 1629 4212 1651
rect 4275 1629 4305 1651
rect 4353 1629 4383 1651
rect 4446 1629 4476 1651
rect 4532 1629 4562 1651
rect 4676 1629 4706 1651
rect 4762 1629 4792 1651
rect 4855 1629 4885 1651
rect 4933 1629 4963 1651
rect 5026 1629 5056 1651
rect 5112 1629 5142 1651
rect 5256 1629 5286 1651
rect 5342 1629 5372 1651
rect 5435 1629 5465 1651
rect 5513 1629 5543 1651
rect 5606 1629 5636 1651
rect 5692 1629 5722 1651
rect 5836 1629 5866 1651
rect 5922 1629 5952 1651
rect 6015 1629 6045 1651
rect 6093 1629 6123 1651
rect 6186 1629 6216 1651
rect 6272 1629 6302 1651
rect 6416 1629 6446 1651
rect 6502 1629 6532 1651
rect 6595 1629 6625 1651
rect 6673 1629 6703 1651
rect 6766 1629 6796 1651
rect 6852 1629 6882 1651
rect -43 1583 6925 1613
rect 100 1555 130 1583
rect 215 1545 245 1567
rect 293 1545 323 1567
rect 408 1555 438 1583
rect 100 1505 130 1527
rect 680 1555 710 1583
rect 795 1545 825 1567
rect 873 1545 903 1567
rect 988 1555 1018 1583
rect 215 1484 245 1517
rect 36 1423 66 1445
rect 122 1423 137 1457
rect 215 1423 245 1450
rect 293 1484 323 1517
rect 408 1505 438 1527
rect 680 1505 710 1527
rect 1260 1555 1290 1583
rect 1375 1545 1405 1567
rect 1453 1545 1483 1567
rect 1568 1555 1598 1583
rect 795 1484 825 1517
rect 293 1423 323 1450
rect 401 1423 416 1457
rect 472 1423 502 1445
rect 616 1423 646 1445
rect 702 1423 717 1457
rect 795 1423 825 1450
rect 873 1484 903 1517
rect 988 1505 1018 1527
rect 1260 1505 1290 1527
rect 1840 1555 1870 1583
rect 1955 1545 1985 1567
rect 2033 1545 2063 1567
rect 2148 1555 2178 1583
rect 1375 1484 1405 1517
rect 873 1423 903 1450
rect 981 1423 996 1457
rect 1052 1423 1082 1445
rect 1196 1423 1226 1445
rect 1282 1423 1297 1457
rect 1375 1423 1405 1450
rect 1453 1484 1483 1517
rect 1568 1505 1598 1527
rect 1840 1505 1870 1527
rect 2420 1555 2450 1583
rect 2535 1545 2565 1567
rect 2613 1545 2643 1567
rect 2728 1555 2758 1583
rect 1955 1484 1985 1517
rect 1453 1423 1483 1450
rect 1561 1423 1576 1457
rect 1632 1423 1662 1445
rect 1776 1423 1806 1445
rect 1862 1423 1877 1457
rect 1955 1423 1985 1450
rect 2033 1484 2063 1517
rect 2148 1505 2178 1527
rect 2420 1505 2450 1527
rect 3000 1555 3030 1583
rect 3115 1545 3145 1567
rect 3193 1545 3223 1567
rect 3308 1555 3338 1583
rect 2535 1484 2565 1517
rect 2033 1423 2063 1450
rect 2141 1423 2156 1457
rect 2212 1423 2242 1445
rect 2356 1423 2386 1445
rect 2442 1423 2457 1457
rect 2535 1423 2565 1450
rect 2613 1484 2643 1517
rect 2728 1505 2758 1527
rect 3000 1505 3030 1527
rect 3580 1555 3610 1583
rect 3695 1545 3725 1567
rect 3773 1545 3803 1567
rect 3888 1555 3918 1583
rect 3115 1484 3145 1517
rect 2613 1423 2643 1450
rect 2721 1423 2736 1457
rect 2792 1423 2822 1445
rect 2936 1423 2966 1445
rect 3022 1423 3037 1457
rect 3115 1423 3145 1450
rect 3193 1484 3223 1517
rect 3308 1505 3338 1527
rect 3580 1505 3610 1527
rect 4160 1555 4190 1583
rect 4275 1545 4305 1567
rect 4353 1545 4383 1567
rect 4468 1555 4498 1583
rect 3695 1484 3725 1517
rect 3193 1423 3223 1450
rect 3301 1423 3316 1457
rect 3372 1423 3402 1445
rect 3516 1423 3546 1445
rect 3602 1423 3617 1457
rect 3695 1423 3725 1450
rect 3773 1484 3803 1517
rect 3888 1505 3918 1527
rect 4160 1505 4190 1527
rect 4740 1555 4770 1583
rect 4855 1545 4885 1567
rect 4933 1545 4963 1567
rect 5048 1555 5078 1583
rect 4275 1484 4305 1517
rect 3773 1423 3803 1450
rect 3881 1423 3896 1457
rect 3952 1423 3982 1445
rect 4096 1423 4126 1445
rect 4182 1423 4197 1457
rect 4275 1423 4305 1450
rect 4353 1484 4383 1517
rect 4468 1505 4498 1527
rect 4740 1505 4770 1527
rect 5320 1555 5350 1583
rect 5435 1545 5465 1567
rect 5513 1545 5543 1567
rect 5628 1555 5658 1583
rect 4855 1484 4885 1517
rect 4353 1423 4383 1450
rect 4461 1423 4476 1457
rect 4532 1423 4562 1445
rect 4676 1423 4706 1445
rect 4762 1423 4777 1457
rect 4855 1423 4885 1450
rect 4933 1484 4963 1517
rect 5048 1505 5078 1527
rect 5320 1505 5350 1527
rect 5900 1555 5930 1583
rect 6015 1545 6045 1567
rect 6093 1545 6123 1567
rect 6208 1555 6238 1583
rect 5435 1484 5465 1517
rect 4933 1423 4963 1450
rect 5041 1423 5056 1457
rect 5112 1423 5142 1445
rect 5256 1423 5286 1445
rect 5342 1423 5357 1457
rect 5435 1423 5465 1450
rect 5513 1484 5543 1517
rect 5628 1505 5658 1527
rect 5900 1505 5930 1527
rect 6480 1555 6510 1583
rect 6595 1545 6625 1567
rect 6673 1545 6703 1567
rect 6788 1555 6818 1583
rect 6015 1484 6045 1517
rect 5513 1423 5543 1450
rect 5621 1423 5636 1457
rect 5692 1423 5722 1445
rect 5836 1423 5866 1445
rect 5922 1423 5937 1457
rect 6015 1423 6045 1450
rect 6093 1484 6123 1517
rect 6208 1505 6238 1527
rect 6480 1505 6510 1527
rect 6595 1484 6625 1517
rect 6093 1423 6123 1450
rect 6201 1423 6216 1457
rect 6272 1423 6302 1445
rect 6416 1423 6446 1445
rect 6502 1423 6517 1457
rect 6595 1423 6625 1450
rect 6673 1484 6703 1517
rect 6788 1505 6818 1527
rect 6673 1423 6703 1450
rect 6781 1423 6796 1457
rect 6852 1423 6882 1445
rect 122 1409 152 1423
rect 386 1409 416 1423
rect 702 1409 732 1423
rect 966 1409 996 1423
rect 1282 1409 1312 1423
rect 1546 1409 1576 1423
rect 1862 1409 1892 1423
rect 2126 1409 2156 1423
rect 2442 1409 2472 1423
rect 2706 1409 2736 1423
rect 3022 1409 3052 1423
rect 3286 1409 3316 1423
rect 3602 1409 3632 1423
rect 3866 1409 3896 1423
rect 4182 1409 4212 1423
rect 4446 1409 4476 1423
rect 4762 1409 4792 1423
rect 5026 1409 5056 1423
rect 5342 1409 5372 1423
rect 5606 1409 5636 1423
rect 5922 1409 5952 1423
rect 6186 1409 6216 1423
rect 6502 1409 6532 1423
rect 6766 1409 6796 1423
rect 36 1359 66 1381
rect 122 1359 152 1381
rect 215 1359 245 1381
rect 293 1359 323 1381
rect 386 1359 416 1381
rect 472 1359 502 1381
rect 616 1359 646 1381
rect 702 1359 732 1381
rect 795 1359 825 1381
rect 873 1359 903 1381
rect 966 1359 996 1381
rect 1052 1359 1082 1381
rect 1196 1359 1226 1381
rect 1282 1359 1312 1381
rect 1375 1359 1405 1381
rect 1453 1359 1483 1381
rect 1546 1359 1576 1381
rect 1632 1359 1662 1381
rect 1776 1359 1806 1381
rect 1862 1359 1892 1381
rect 1955 1359 1985 1381
rect 2033 1359 2063 1381
rect 2126 1359 2156 1381
rect 2212 1359 2242 1381
rect 2356 1359 2386 1381
rect 2442 1359 2472 1381
rect 2535 1359 2565 1381
rect 2613 1359 2643 1381
rect 2706 1359 2736 1381
rect 2792 1359 2822 1381
rect 2936 1359 2966 1381
rect 3022 1359 3052 1381
rect 3115 1359 3145 1381
rect 3193 1359 3223 1381
rect 3286 1359 3316 1381
rect 3372 1359 3402 1381
rect 3516 1359 3546 1381
rect 3602 1359 3632 1381
rect 3695 1359 3725 1381
rect 3773 1359 3803 1381
rect 3866 1359 3896 1381
rect 3952 1359 3982 1381
rect 4096 1359 4126 1381
rect 4182 1359 4212 1381
rect 4275 1359 4305 1381
rect 4353 1359 4383 1381
rect 4446 1359 4476 1381
rect 4532 1359 4562 1381
rect 4676 1359 4706 1381
rect 4762 1359 4792 1381
rect 4855 1359 4885 1381
rect 4933 1359 4963 1381
rect 5026 1359 5056 1381
rect 5112 1359 5142 1381
rect 5256 1359 5286 1381
rect 5342 1359 5372 1381
rect 5435 1359 5465 1381
rect 5513 1359 5543 1381
rect 5606 1359 5636 1381
rect 5692 1359 5722 1381
rect 5836 1359 5866 1381
rect 5922 1359 5952 1381
rect 6015 1359 6045 1381
rect 6093 1359 6123 1381
rect 6186 1359 6216 1381
rect 6272 1359 6302 1381
rect 6416 1359 6446 1381
rect 6502 1359 6532 1381
rect 6595 1359 6625 1381
rect 6673 1359 6703 1381
rect 6766 1359 6796 1381
rect 6852 1359 6882 1381
rect -43 1313 6925 1343
rect 100 1285 130 1313
rect 215 1275 245 1297
rect 293 1275 323 1297
rect 408 1285 438 1313
rect 100 1235 130 1257
rect 680 1285 710 1313
rect 795 1275 825 1297
rect 873 1275 903 1297
rect 988 1285 1018 1313
rect 215 1214 245 1247
rect 36 1153 66 1175
rect 122 1153 137 1187
rect 215 1153 245 1180
rect 293 1214 323 1247
rect 408 1235 438 1257
rect 680 1235 710 1257
rect 1260 1285 1290 1313
rect 1375 1275 1405 1297
rect 1453 1275 1483 1297
rect 1568 1285 1598 1313
rect 795 1214 825 1247
rect 293 1153 323 1180
rect 401 1153 416 1187
rect 472 1153 502 1175
rect 616 1153 646 1175
rect 702 1153 717 1187
rect 795 1153 825 1180
rect 873 1214 903 1247
rect 988 1235 1018 1257
rect 1260 1235 1290 1257
rect 1840 1285 1870 1313
rect 1955 1275 1985 1297
rect 2033 1275 2063 1297
rect 2148 1285 2178 1313
rect 1375 1214 1405 1247
rect 873 1153 903 1180
rect 981 1153 996 1187
rect 1052 1153 1082 1175
rect 1196 1153 1226 1175
rect 1282 1153 1297 1187
rect 1375 1153 1405 1180
rect 1453 1214 1483 1247
rect 1568 1235 1598 1257
rect 1840 1235 1870 1257
rect 2420 1285 2450 1313
rect 2535 1275 2565 1297
rect 2613 1275 2643 1297
rect 2728 1285 2758 1313
rect 1955 1214 1985 1247
rect 1453 1153 1483 1180
rect 1561 1153 1576 1187
rect 1632 1153 1662 1175
rect 1776 1153 1806 1175
rect 1862 1153 1877 1187
rect 1955 1153 1985 1180
rect 2033 1214 2063 1247
rect 2148 1235 2178 1257
rect 2420 1235 2450 1257
rect 3000 1285 3030 1313
rect 3115 1275 3145 1297
rect 3193 1275 3223 1297
rect 3308 1285 3338 1313
rect 2535 1214 2565 1247
rect 2033 1153 2063 1180
rect 2141 1153 2156 1187
rect 2212 1153 2242 1175
rect 2356 1153 2386 1175
rect 2442 1153 2457 1187
rect 2535 1153 2565 1180
rect 2613 1214 2643 1247
rect 2728 1235 2758 1257
rect 3000 1235 3030 1257
rect 3580 1285 3610 1313
rect 3695 1275 3725 1297
rect 3773 1275 3803 1297
rect 3888 1285 3918 1313
rect 3115 1214 3145 1247
rect 2613 1153 2643 1180
rect 2721 1153 2736 1187
rect 2792 1153 2822 1175
rect 2936 1153 2966 1175
rect 3022 1153 3037 1187
rect 3115 1153 3145 1180
rect 3193 1214 3223 1247
rect 3308 1235 3338 1257
rect 3580 1235 3610 1257
rect 4160 1285 4190 1313
rect 4275 1275 4305 1297
rect 4353 1275 4383 1297
rect 4468 1285 4498 1313
rect 3695 1214 3725 1247
rect 3193 1153 3223 1180
rect 3301 1153 3316 1187
rect 3372 1153 3402 1175
rect 3516 1153 3546 1175
rect 3602 1153 3617 1187
rect 3695 1153 3725 1180
rect 3773 1214 3803 1247
rect 3888 1235 3918 1257
rect 4160 1235 4190 1257
rect 4740 1285 4770 1313
rect 4855 1275 4885 1297
rect 4933 1275 4963 1297
rect 5048 1285 5078 1313
rect 4275 1214 4305 1247
rect 3773 1153 3803 1180
rect 3881 1153 3896 1187
rect 3952 1153 3982 1175
rect 4096 1153 4126 1175
rect 4182 1153 4197 1187
rect 4275 1153 4305 1180
rect 4353 1214 4383 1247
rect 4468 1235 4498 1257
rect 4740 1235 4770 1257
rect 5320 1285 5350 1313
rect 5435 1275 5465 1297
rect 5513 1275 5543 1297
rect 5628 1285 5658 1313
rect 4855 1214 4885 1247
rect 4353 1153 4383 1180
rect 4461 1153 4476 1187
rect 4532 1153 4562 1175
rect 4676 1153 4706 1175
rect 4762 1153 4777 1187
rect 4855 1153 4885 1180
rect 4933 1214 4963 1247
rect 5048 1235 5078 1257
rect 5320 1235 5350 1257
rect 5900 1285 5930 1313
rect 6015 1275 6045 1297
rect 6093 1275 6123 1297
rect 6208 1285 6238 1313
rect 5435 1214 5465 1247
rect 4933 1153 4963 1180
rect 5041 1153 5056 1187
rect 5112 1153 5142 1175
rect 5256 1153 5286 1175
rect 5342 1153 5357 1187
rect 5435 1153 5465 1180
rect 5513 1214 5543 1247
rect 5628 1235 5658 1257
rect 5900 1235 5930 1257
rect 6480 1285 6510 1313
rect 6595 1275 6625 1297
rect 6673 1275 6703 1297
rect 6788 1285 6818 1313
rect 6015 1214 6045 1247
rect 5513 1153 5543 1180
rect 5621 1153 5636 1187
rect 5692 1153 5722 1175
rect 5836 1153 5866 1175
rect 5922 1153 5937 1187
rect 6015 1153 6045 1180
rect 6093 1214 6123 1247
rect 6208 1235 6238 1257
rect 6480 1235 6510 1257
rect 6595 1214 6625 1247
rect 6093 1153 6123 1180
rect 6201 1153 6216 1187
rect 6272 1153 6302 1175
rect 6416 1153 6446 1175
rect 6502 1153 6517 1187
rect 6595 1153 6625 1180
rect 6673 1214 6703 1247
rect 6788 1235 6818 1257
rect 6673 1153 6703 1180
rect 6781 1153 6796 1187
rect 6852 1153 6882 1175
rect 122 1139 152 1153
rect 386 1139 416 1153
rect 702 1139 732 1153
rect 966 1139 996 1153
rect 1282 1139 1312 1153
rect 1546 1139 1576 1153
rect 1862 1139 1892 1153
rect 2126 1139 2156 1153
rect 2442 1139 2472 1153
rect 2706 1139 2736 1153
rect 3022 1139 3052 1153
rect 3286 1139 3316 1153
rect 3602 1139 3632 1153
rect 3866 1139 3896 1153
rect 4182 1139 4212 1153
rect 4446 1139 4476 1153
rect 4762 1139 4792 1153
rect 5026 1139 5056 1153
rect 5342 1139 5372 1153
rect 5606 1139 5636 1153
rect 5922 1139 5952 1153
rect 6186 1139 6216 1153
rect 6502 1139 6532 1153
rect 6766 1139 6796 1153
rect 36 1089 66 1111
rect 122 1089 152 1111
rect 215 1089 245 1111
rect 293 1089 323 1111
rect 386 1089 416 1111
rect 472 1089 502 1111
rect 616 1089 646 1111
rect 702 1089 732 1111
rect 795 1089 825 1111
rect 873 1089 903 1111
rect 966 1089 996 1111
rect 1052 1089 1082 1111
rect 1196 1089 1226 1111
rect 1282 1089 1312 1111
rect 1375 1089 1405 1111
rect 1453 1089 1483 1111
rect 1546 1089 1576 1111
rect 1632 1089 1662 1111
rect 1776 1089 1806 1111
rect 1862 1089 1892 1111
rect 1955 1089 1985 1111
rect 2033 1089 2063 1111
rect 2126 1089 2156 1111
rect 2212 1089 2242 1111
rect 2356 1089 2386 1111
rect 2442 1089 2472 1111
rect 2535 1089 2565 1111
rect 2613 1089 2643 1111
rect 2706 1089 2736 1111
rect 2792 1089 2822 1111
rect 2936 1089 2966 1111
rect 3022 1089 3052 1111
rect 3115 1089 3145 1111
rect 3193 1089 3223 1111
rect 3286 1089 3316 1111
rect 3372 1089 3402 1111
rect 3516 1089 3546 1111
rect 3602 1089 3632 1111
rect 3695 1089 3725 1111
rect 3773 1089 3803 1111
rect 3866 1089 3896 1111
rect 3952 1089 3982 1111
rect 4096 1089 4126 1111
rect 4182 1089 4212 1111
rect 4275 1089 4305 1111
rect 4353 1089 4383 1111
rect 4446 1089 4476 1111
rect 4532 1089 4562 1111
rect 4676 1089 4706 1111
rect 4762 1089 4792 1111
rect 4855 1089 4885 1111
rect 4933 1089 4963 1111
rect 5026 1089 5056 1111
rect 5112 1089 5142 1111
rect 5256 1089 5286 1111
rect 5342 1089 5372 1111
rect 5435 1089 5465 1111
rect 5513 1089 5543 1111
rect 5606 1089 5636 1111
rect 5692 1089 5722 1111
rect 5836 1089 5866 1111
rect 5922 1089 5952 1111
rect 6015 1089 6045 1111
rect 6093 1089 6123 1111
rect 6186 1089 6216 1111
rect 6272 1089 6302 1111
rect 6416 1089 6446 1111
rect 6502 1089 6532 1111
rect 6595 1089 6625 1111
rect 6673 1089 6703 1111
rect 6766 1089 6796 1111
rect 6852 1089 6882 1111
rect -43 1043 6925 1073
rect 100 1015 130 1043
rect 215 1005 245 1027
rect 293 1005 323 1027
rect 408 1015 438 1043
rect 100 965 130 987
rect 680 1015 710 1043
rect 795 1005 825 1027
rect 873 1005 903 1027
rect 988 1015 1018 1043
rect 215 944 245 977
rect 36 883 66 905
rect 122 883 137 917
rect 215 883 245 910
rect 293 944 323 977
rect 408 965 438 987
rect 680 965 710 987
rect 1260 1015 1290 1043
rect 1375 1005 1405 1027
rect 1453 1005 1483 1027
rect 1568 1015 1598 1043
rect 795 944 825 977
rect 293 883 323 910
rect 401 883 416 917
rect 472 883 502 905
rect 616 883 646 905
rect 702 883 717 917
rect 795 883 825 910
rect 873 944 903 977
rect 988 965 1018 987
rect 1260 965 1290 987
rect 1840 1015 1870 1043
rect 1955 1005 1985 1027
rect 2033 1005 2063 1027
rect 2148 1015 2178 1043
rect 1375 944 1405 977
rect 873 883 903 910
rect 981 883 996 917
rect 1052 883 1082 905
rect 1196 883 1226 905
rect 1282 883 1297 917
rect 1375 883 1405 910
rect 1453 944 1483 977
rect 1568 965 1598 987
rect 1840 965 1870 987
rect 2420 1015 2450 1043
rect 2535 1005 2565 1027
rect 2613 1005 2643 1027
rect 2728 1015 2758 1043
rect 1955 944 1985 977
rect 1453 883 1483 910
rect 1561 883 1576 917
rect 1632 883 1662 905
rect 1776 883 1806 905
rect 1862 883 1877 917
rect 1955 883 1985 910
rect 2033 944 2063 977
rect 2148 965 2178 987
rect 2420 965 2450 987
rect 3000 1015 3030 1043
rect 3115 1005 3145 1027
rect 3193 1005 3223 1027
rect 3308 1015 3338 1043
rect 2535 944 2565 977
rect 2033 883 2063 910
rect 2141 883 2156 917
rect 2212 883 2242 905
rect 2356 883 2386 905
rect 2442 883 2457 917
rect 2535 883 2565 910
rect 2613 944 2643 977
rect 2728 965 2758 987
rect 3000 965 3030 987
rect 3580 1015 3610 1043
rect 3695 1005 3725 1027
rect 3773 1005 3803 1027
rect 3888 1015 3918 1043
rect 3115 944 3145 977
rect 2613 883 2643 910
rect 2721 883 2736 917
rect 2792 883 2822 905
rect 2936 883 2966 905
rect 3022 883 3037 917
rect 3115 883 3145 910
rect 3193 944 3223 977
rect 3308 965 3338 987
rect 3580 965 3610 987
rect 4160 1015 4190 1043
rect 4275 1005 4305 1027
rect 4353 1005 4383 1027
rect 4468 1015 4498 1043
rect 3695 944 3725 977
rect 3193 883 3223 910
rect 3301 883 3316 917
rect 3372 883 3402 905
rect 3516 883 3546 905
rect 3602 883 3617 917
rect 3695 883 3725 910
rect 3773 944 3803 977
rect 3888 965 3918 987
rect 4160 965 4190 987
rect 4740 1015 4770 1043
rect 4855 1005 4885 1027
rect 4933 1005 4963 1027
rect 5048 1015 5078 1043
rect 4275 944 4305 977
rect 3773 883 3803 910
rect 3881 883 3896 917
rect 3952 883 3982 905
rect 4096 883 4126 905
rect 4182 883 4197 917
rect 4275 883 4305 910
rect 4353 944 4383 977
rect 4468 965 4498 987
rect 4740 965 4770 987
rect 5320 1015 5350 1043
rect 5435 1005 5465 1027
rect 5513 1005 5543 1027
rect 5628 1015 5658 1043
rect 4855 944 4885 977
rect 4353 883 4383 910
rect 4461 883 4476 917
rect 4532 883 4562 905
rect 4676 883 4706 905
rect 4762 883 4777 917
rect 4855 883 4885 910
rect 4933 944 4963 977
rect 5048 965 5078 987
rect 5320 965 5350 987
rect 5900 1015 5930 1043
rect 6015 1005 6045 1027
rect 6093 1005 6123 1027
rect 6208 1015 6238 1043
rect 5435 944 5465 977
rect 4933 883 4963 910
rect 5041 883 5056 917
rect 5112 883 5142 905
rect 5256 883 5286 905
rect 5342 883 5357 917
rect 5435 883 5465 910
rect 5513 944 5543 977
rect 5628 965 5658 987
rect 5900 965 5930 987
rect 6480 1015 6510 1043
rect 6595 1005 6625 1027
rect 6673 1005 6703 1027
rect 6788 1015 6818 1043
rect 6015 944 6045 977
rect 5513 883 5543 910
rect 5621 883 5636 917
rect 5692 883 5722 905
rect 5836 883 5866 905
rect 5922 883 5937 917
rect 6015 883 6045 910
rect 6093 944 6123 977
rect 6208 965 6238 987
rect 6480 965 6510 987
rect 6595 944 6625 977
rect 6093 883 6123 910
rect 6201 883 6216 917
rect 6272 883 6302 905
rect 6416 883 6446 905
rect 6502 883 6517 917
rect 6595 883 6625 910
rect 6673 944 6703 977
rect 6788 965 6818 987
rect 6673 883 6703 910
rect 6781 883 6796 917
rect 6852 883 6882 905
rect 122 869 152 883
rect 386 869 416 883
rect 702 869 732 883
rect 966 869 996 883
rect 1282 869 1312 883
rect 1546 869 1576 883
rect 1862 869 1892 883
rect 2126 869 2156 883
rect 2442 869 2472 883
rect 2706 869 2736 883
rect 3022 869 3052 883
rect 3286 869 3316 883
rect 3602 869 3632 883
rect 3866 869 3896 883
rect 4182 869 4212 883
rect 4446 869 4476 883
rect 4762 869 4792 883
rect 5026 869 5056 883
rect 5342 869 5372 883
rect 5606 869 5636 883
rect 5922 869 5952 883
rect 6186 869 6216 883
rect 6502 869 6532 883
rect 6766 869 6796 883
rect 36 819 66 841
rect 122 819 152 841
rect 215 819 245 841
rect 293 819 323 841
rect 386 819 416 841
rect 472 819 502 841
rect 616 819 646 841
rect 702 819 732 841
rect 795 819 825 841
rect 873 819 903 841
rect 966 819 996 841
rect 1052 819 1082 841
rect 1196 819 1226 841
rect 1282 819 1312 841
rect 1375 819 1405 841
rect 1453 819 1483 841
rect 1546 819 1576 841
rect 1632 819 1662 841
rect 1776 819 1806 841
rect 1862 819 1892 841
rect 1955 819 1985 841
rect 2033 819 2063 841
rect 2126 819 2156 841
rect 2212 819 2242 841
rect 2356 819 2386 841
rect 2442 819 2472 841
rect 2535 819 2565 841
rect 2613 819 2643 841
rect 2706 819 2736 841
rect 2792 819 2822 841
rect 2936 819 2966 841
rect 3022 819 3052 841
rect 3115 819 3145 841
rect 3193 819 3223 841
rect 3286 819 3316 841
rect 3372 819 3402 841
rect 3516 819 3546 841
rect 3602 819 3632 841
rect 3695 819 3725 841
rect 3773 819 3803 841
rect 3866 819 3896 841
rect 3952 819 3982 841
rect 4096 819 4126 841
rect 4182 819 4212 841
rect 4275 819 4305 841
rect 4353 819 4383 841
rect 4446 819 4476 841
rect 4532 819 4562 841
rect 4676 819 4706 841
rect 4762 819 4792 841
rect 4855 819 4885 841
rect 4933 819 4963 841
rect 5026 819 5056 841
rect 5112 819 5142 841
rect 5256 819 5286 841
rect 5342 819 5372 841
rect 5435 819 5465 841
rect 5513 819 5543 841
rect 5606 819 5636 841
rect 5692 819 5722 841
rect 5836 819 5866 841
rect 5922 819 5952 841
rect 6015 819 6045 841
rect 6093 819 6123 841
rect 6186 819 6216 841
rect 6272 819 6302 841
rect 6416 819 6446 841
rect 6502 819 6532 841
rect 6595 819 6625 841
rect 6673 819 6703 841
rect 6766 819 6796 841
rect 6852 819 6882 841
rect -43 773 6925 803
rect 100 745 130 773
rect 215 735 245 757
rect 293 735 323 757
rect 408 745 438 773
rect 100 695 130 717
rect 680 745 710 773
rect 795 735 825 757
rect 873 735 903 757
rect 988 745 1018 773
rect 215 674 245 707
rect 36 613 66 635
rect 122 613 137 647
rect 215 613 245 640
rect 293 674 323 707
rect 408 695 438 717
rect 680 695 710 717
rect 1260 745 1290 773
rect 1375 735 1405 757
rect 1453 735 1483 757
rect 1568 745 1598 773
rect 795 674 825 707
rect 293 613 323 640
rect 401 613 416 647
rect 472 613 502 635
rect 616 613 646 635
rect 702 613 717 647
rect 795 613 825 640
rect 873 674 903 707
rect 988 695 1018 717
rect 1260 695 1290 717
rect 1840 745 1870 773
rect 1955 735 1985 757
rect 2033 735 2063 757
rect 2148 745 2178 773
rect 1375 674 1405 707
rect 873 613 903 640
rect 981 613 996 647
rect 1052 613 1082 635
rect 1196 613 1226 635
rect 1282 613 1297 647
rect 1375 613 1405 640
rect 1453 674 1483 707
rect 1568 695 1598 717
rect 1840 695 1870 717
rect 2420 745 2450 773
rect 2535 735 2565 757
rect 2613 735 2643 757
rect 2728 745 2758 773
rect 1955 674 1985 707
rect 1453 613 1483 640
rect 1561 613 1576 647
rect 1632 613 1662 635
rect 1776 613 1806 635
rect 1862 613 1877 647
rect 1955 613 1985 640
rect 2033 674 2063 707
rect 2148 695 2178 717
rect 2420 695 2450 717
rect 3000 745 3030 773
rect 3115 735 3145 757
rect 3193 735 3223 757
rect 3308 745 3338 773
rect 2535 674 2565 707
rect 2033 613 2063 640
rect 2141 613 2156 647
rect 2212 613 2242 635
rect 2356 613 2386 635
rect 2442 613 2457 647
rect 2535 613 2565 640
rect 2613 674 2643 707
rect 2728 695 2758 717
rect 3000 695 3030 717
rect 3580 745 3610 773
rect 3695 735 3725 757
rect 3773 735 3803 757
rect 3888 745 3918 773
rect 3115 674 3145 707
rect 2613 613 2643 640
rect 2721 613 2736 647
rect 2792 613 2822 635
rect 2936 613 2966 635
rect 3022 613 3037 647
rect 3115 613 3145 640
rect 3193 674 3223 707
rect 3308 695 3338 717
rect 3580 695 3610 717
rect 4160 745 4190 773
rect 4275 735 4305 757
rect 4353 735 4383 757
rect 4468 745 4498 773
rect 3695 674 3725 707
rect 3193 613 3223 640
rect 3301 613 3316 647
rect 3372 613 3402 635
rect 3516 613 3546 635
rect 3602 613 3617 647
rect 3695 613 3725 640
rect 3773 674 3803 707
rect 3888 695 3918 717
rect 4160 695 4190 717
rect 4740 745 4770 773
rect 4855 735 4885 757
rect 4933 735 4963 757
rect 5048 745 5078 773
rect 4275 674 4305 707
rect 3773 613 3803 640
rect 3881 613 3896 647
rect 3952 613 3982 635
rect 4096 613 4126 635
rect 4182 613 4197 647
rect 4275 613 4305 640
rect 4353 674 4383 707
rect 4468 695 4498 717
rect 4740 695 4770 717
rect 5320 745 5350 773
rect 5435 735 5465 757
rect 5513 735 5543 757
rect 5628 745 5658 773
rect 4855 674 4885 707
rect 4353 613 4383 640
rect 4461 613 4476 647
rect 4532 613 4562 635
rect 4676 613 4706 635
rect 4762 613 4777 647
rect 4855 613 4885 640
rect 4933 674 4963 707
rect 5048 695 5078 717
rect 5320 695 5350 717
rect 5900 745 5930 773
rect 6015 735 6045 757
rect 6093 735 6123 757
rect 6208 745 6238 773
rect 5435 674 5465 707
rect 4933 613 4963 640
rect 5041 613 5056 647
rect 5112 613 5142 635
rect 5256 613 5286 635
rect 5342 613 5357 647
rect 5435 613 5465 640
rect 5513 674 5543 707
rect 5628 695 5658 717
rect 5900 695 5930 717
rect 6480 745 6510 773
rect 6595 735 6625 757
rect 6673 735 6703 757
rect 6788 745 6818 773
rect 6015 674 6045 707
rect 5513 613 5543 640
rect 5621 613 5636 647
rect 5692 613 5722 635
rect 5836 613 5866 635
rect 5922 613 5937 647
rect 6015 613 6045 640
rect 6093 674 6123 707
rect 6208 695 6238 717
rect 6480 695 6510 717
rect 6595 674 6625 707
rect 6093 613 6123 640
rect 6201 613 6216 647
rect 6272 613 6302 635
rect 6416 613 6446 635
rect 6502 613 6517 647
rect 6595 613 6625 640
rect 6673 674 6703 707
rect 6788 695 6818 717
rect 6673 613 6703 640
rect 6781 613 6796 647
rect 6852 613 6882 635
rect 122 599 152 613
rect 386 599 416 613
rect 702 599 732 613
rect 966 599 996 613
rect 1282 599 1312 613
rect 1546 599 1576 613
rect 1862 599 1892 613
rect 2126 599 2156 613
rect 2442 599 2472 613
rect 2706 599 2736 613
rect 3022 599 3052 613
rect 3286 599 3316 613
rect 3602 599 3632 613
rect 3866 599 3896 613
rect 4182 599 4212 613
rect 4446 599 4476 613
rect 4762 599 4792 613
rect 5026 599 5056 613
rect 5342 599 5372 613
rect 5606 599 5636 613
rect 5922 599 5952 613
rect 6186 599 6216 613
rect 6502 599 6532 613
rect 6766 599 6796 613
rect 36 549 66 571
rect 122 549 152 571
rect 215 549 245 571
rect 293 549 323 571
rect 386 549 416 571
rect 472 549 502 571
rect 616 549 646 571
rect 702 549 732 571
rect 795 549 825 571
rect 873 549 903 571
rect 966 549 996 571
rect 1052 549 1082 571
rect 1196 549 1226 571
rect 1282 549 1312 571
rect 1375 549 1405 571
rect 1453 549 1483 571
rect 1546 549 1576 571
rect 1632 549 1662 571
rect 1776 549 1806 571
rect 1862 549 1892 571
rect 1955 549 1985 571
rect 2033 549 2063 571
rect 2126 549 2156 571
rect 2212 549 2242 571
rect 2356 549 2386 571
rect 2442 549 2472 571
rect 2535 549 2565 571
rect 2613 549 2643 571
rect 2706 549 2736 571
rect 2792 549 2822 571
rect 2936 549 2966 571
rect 3022 549 3052 571
rect 3115 549 3145 571
rect 3193 549 3223 571
rect 3286 549 3316 571
rect 3372 549 3402 571
rect 3516 549 3546 571
rect 3602 549 3632 571
rect 3695 549 3725 571
rect 3773 549 3803 571
rect 3866 549 3896 571
rect 3952 549 3982 571
rect 4096 549 4126 571
rect 4182 549 4212 571
rect 4275 549 4305 571
rect 4353 549 4383 571
rect 4446 549 4476 571
rect 4532 549 4562 571
rect 4676 549 4706 571
rect 4762 549 4792 571
rect 4855 549 4885 571
rect 4933 549 4963 571
rect 5026 549 5056 571
rect 5112 549 5142 571
rect 5256 549 5286 571
rect 5342 549 5372 571
rect 5435 549 5465 571
rect 5513 549 5543 571
rect 5606 549 5636 571
rect 5692 549 5722 571
rect 5836 549 5866 571
rect 5922 549 5952 571
rect 6015 549 6045 571
rect 6093 549 6123 571
rect 6186 549 6216 571
rect 6272 549 6302 571
rect 6416 549 6446 571
rect 6502 549 6532 571
rect 6595 549 6625 571
rect 6673 549 6703 571
rect 6766 549 6796 571
rect 6852 549 6882 571
rect -43 503 6925 533
rect 100 475 130 503
rect 215 465 245 487
rect 293 465 323 487
rect 408 475 438 503
rect 100 425 130 447
rect 680 475 710 503
rect 795 465 825 487
rect 873 465 903 487
rect 988 475 1018 503
rect 215 404 245 437
rect 36 343 66 365
rect 122 343 137 377
rect 215 343 245 370
rect 293 404 323 437
rect 408 425 438 447
rect 680 425 710 447
rect 1260 475 1290 503
rect 1375 465 1405 487
rect 1453 465 1483 487
rect 1568 475 1598 503
rect 795 404 825 437
rect 293 343 323 370
rect 401 343 416 377
rect 472 343 502 365
rect 616 343 646 365
rect 702 343 717 377
rect 795 343 825 370
rect 873 404 903 437
rect 988 425 1018 447
rect 1260 425 1290 447
rect 1840 475 1870 503
rect 1955 465 1985 487
rect 2033 465 2063 487
rect 2148 475 2178 503
rect 1375 404 1405 437
rect 873 343 903 370
rect 981 343 996 377
rect 1052 343 1082 365
rect 1196 343 1226 365
rect 1282 343 1297 377
rect 1375 343 1405 370
rect 1453 404 1483 437
rect 1568 425 1598 447
rect 1840 425 1870 447
rect 2420 475 2450 503
rect 2535 465 2565 487
rect 2613 465 2643 487
rect 2728 475 2758 503
rect 1955 404 1985 437
rect 1453 343 1483 370
rect 1561 343 1576 377
rect 1632 343 1662 365
rect 1776 343 1806 365
rect 1862 343 1877 377
rect 1955 343 1985 370
rect 2033 404 2063 437
rect 2148 425 2178 447
rect 2420 425 2450 447
rect 3000 475 3030 503
rect 3115 465 3145 487
rect 3193 465 3223 487
rect 3308 475 3338 503
rect 2535 404 2565 437
rect 2033 343 2063 370
rect 2141 343 2156 377
rect 2212 343 2242 365
rect 2356 343 2386 365
rect 2442 343 2457 377
rect 2535 343 2565 370
rect 2613 404 2643 437
rect 2728 425 2758 447
rect 3000 425 3030 447
rect 3580 475 3610 503
rect 3695 465 3725 487
rect 3773 465 3803 487
rect 3888 475 3918 503
rect 3115 404 3145 437
rect 2613 343 2643 370
rect 2721 343 2736 377
rect 2792 343 2822 365
rect 2936 343 2966 365
rect 3022 343 3037 377
rect 3115 343 3145 370
rect 3193 404 3223 437
rect 3308 425 3338 447
rect 3580 425 3610 447
rect 4160 475 4190 503
rect 4275 465 4305 487
rect 4353 465 4383 487
rect 4468 475 4498 503
rect 3695 404 3725 437
rect 3193 343 3223 370
rect 3301 343 3316 377
rect 3372 343 3402 365
rect 3516 343 3546 365
rect 3602 343 3617 377
rect 3695 343 3725 370
rect 3773 404 3803 437
rect 3888 425 3918 447
rect 4160 425 4190 447
rect 4740 475 4770 503
rect 4855 465 4885 487
rect 4933 465 4963 487
rect 5048 475 5078 503
rect 4275 404 4305 437
rect 3773 343 3803 370
rect 3881 343 3896 377
rect 3952 343 3982 365
rect 4096 343 4126 365
rect 4182 343 4197 377
rect 4275 343 4305 370
rect 4353 404 4383 437
rect 4468 425 4498 447
rect 4740 425 4770 447
rect 5320 475 5350 503
rect 5435 465 5465 487
rect 5513 465 5543 487
rect 5628 475 5658 503
rect 4855 404 4885 437
rect 4353 343 4383 370
rect 4461 343 4476 377
rect 4532 343 4562 365
rect 4676 343 4706 365
rect 4762 343 4777 377
rect 4855 343 4885 370
rect 4933 404 4963 437
rect 5048 425 5078 447
rect 5320 425 5350 447
rect 5900 475 5930 503
rect 6015 465 6045 487
rect 6093 465 6123 487
rect 6208 475 6238 503
rect 5435 404 5465 437
rect 4933 343 4963 370
rect 5041 343 5056 377
rect 5112 343 5142 365
rect 5256 343 5286 365
rect 5342 343 5357 377
rect 5435 343 5465 370
rect 5513 404 5543 437
rect 5628 425 5658 447
rect 5900 425 5930 447
rect 6480 475 6510 503
rect 6595 465 6625 487
rect 6673 465 6703 487
rect 6788 475 6818 503
rect 6015 404 6045 437
rect 5513 343 5543 370
rect 5621 343 5636 377
rect 5692 343 5722 365
rect 5836 343 5866 365
rect 5922 343 5937 377
rect 6015 343 6045 370
rect 6093 404 6123 437
rect 6208 425 6238 447
rect 6480 425 6510 447
rect 6595 404 6625 437
rect 6093 343 6123 370
rect 6201 343 6216 377
rect 6272 343 6302 365
rect 6416 343 6446 365
rect 6502 343 6517 377
rect 6595 343 6625 370
rect 6673 404 6703 437
rect 6788 425 6818 447
rect 6673 343 6703 370
rect 6781 343 6796 377
rect 6852 343 6882 365
rect 122 329 152 343
rect 386 329 416 343
rect 702 329 732 343
rect 966 329 996 343
rect 1282 329 1312 343
rect 1546 329 1576 343
rect 1862 329 1892 343
rect 2126 329 2156 343
rect 2442 329 2472 343
rect 2706 329 2736 343
rect 3022 329 3052 343
rect 3286 329 3316 343
rect 3602 329 3632 343
rect 3866 329 3896 343
rect 4182 329 4212 343
rect 4446 329 4476 343
rect 4762 329 4792 343
rect 5026 329 5056 343
rect 5342 329 5372 343
rect 5606 329 5636 343
rect 5922 329 5952 343
rect 6186 329 6216 343
rect 6502 329 6532 343
rect 6766 329 6796 343
rect 36 279 66 301
rect 122 279 152 301
rect 215 279 245 301
rect 293 279 323 301
rect 386 279 416 301
rect 472 279 502 301
rect 616 279 646 301
rect 702 279 732 301
rect 795 279 825 301
rect 873 279 903 301
rect 966 279 996 301
rect 1052 279 1082 301
rect 1196 279 1226 301
rect 1282 279 1312 301
rect 1375 279 1405 301
rect 1453 279 1483 301
rect 1546 279 1576 301
rect 1632 279 1662 301
rect 1776 279 1806 301
rect 1862 279 1892 301
rect 1955 279 1985 301
rect 2033 279 2063 301
rect 2126 279 2156 301
rect 2212 279 2242 301
rect 2356 279 2386 301
rect 2442 279 2472 301
rect 2535 279 2565 301
rect 2613 279 2643 301
rect 2706 279 2736 301
rect 2792 279 2822 301
rect 2936 279 2966 301
rect 3022 279 3052 301
rect 3115 279 3145 301
rect 3193 279 3223 301
rect 3286 279 3316 301
rect 3372 279 3402 301
rect 3516 279 3546 301
rect 3602 279 3632 301
rect 3695 279 3725 301
rect 3773 279 3803 301
rect 3866 279 3896 301
rect 3952 279 3982 301
rect 4096 279 4126 301
rect 4182 279 4212 301
rect 4275 279 4305 301
rect 4353 279 4383 301
rect 4446 279 4476 301
rect 4532 279 4562 301
rect 4676 279 4706 301
rect 4762 279 4792 301
rect 4855 279 4885 301
rect 4933 279 4963 301
rect 5026 279 5056 301
rect 5112 279 5142 301
rect 5256 279 5286 301
rect 5342 279 5372 301
rect 5435 279 5465 301
rect 5513 279 5543 301
rect 5606 279 5636 301
rect 5692 279 5722 301
rect 5836 279 5866 301
rect 5922 279 5952 301
rect 6015 279 6045 301
rect 6093 279 6123 301
rect 6186 279 6216 301
rect 6272 279 6302 301
rect 6416 279 6446 301
rect 6502 279 6532 301
rect 6595 279 6625 301
rect 6673 279 6703 301
rect 6766 279 6796 301
rect 6852 279 6882 301
rect -43 233 6925 263
rect 100 205 130 233
rect 215 195 245 217
rect 293 195 323 217
rect 408 205 438 233
rect 100 155 130 177
rect 680 205 710 233
rect 795 195 825 217
rect 873 195 903 217
rect 988 205 1018 233
rect 215 134 245 167
rect 36 73 66 95
rect 122 73 137 107
rect 215 73 245 100
rect 293 134 323 167
rect 408 155 438 177
rect 680 155 710 177
rect 1260 205 1290 233
rect 1375 195 1405 217
rect 1453 195 1483 217
rect 1568 205 1598 233
rect 795 134 825 167
rect 293 73 323 100
rect 401 73 416 107
rect 472 73 502 95
rect 616 73 646 95
rect 702 73 717 107
rect 795 73 825 100
rect 873 134 903 167
rect 988 155 1018 177
rect 1260 155 1290 177
rect 1840 205 1870 233
rect 1955 195 1985 217
rect 2033 195 2063 217
rect 2148 205 2178 233
rect 1375 134 1405 167
rect 873 73 903 100
rect 981 73 996 107
rect 1052 73 1082 95
rect 1196 73 1226 95
rect 1282 73 1297 107
rect 1375 73 1405 100
rect 1453 134 1483 167
rect 1568 155 1598 177
rect 1840 155 1870 177
rect 2420 205 2450 233
rect 2535 195 2565 217
rect 2613 195 2643 217
rect 2728 205 2758 233
rect 1955 134 1985 167
rect 1453 73 1483 100
rect 1561 73 1576 107
rect 1632 73 1662 95
rect 1776 73 1806 95
rect 1862 73 1877 107
rect 1955 73 1985 100
rect 2033 134 2063 167
rect 2148 155 2178 177
rect 2420 155 2450 177
rect 3000 205 3030 233
rect 3115 195 3145 217
rect 3193 195 3223 217
rect 3308 205 3338 233
rect 2535 134 2565 167
rect 2033 73 2063 100
rect 2141 73 2156 107
rect 2212 73 2242 95
rect 2356 73 2386 95
rect 2442 73 2457 107
rect 2535 73 2565 100
rect 2613 134 2643 167
rect 2728 155 2758 177
rect 3000 155 3030 177
rect 3580 205 3610 233
rect 3695 195 3725 217
rect 3773 195 3803 217
rect 3888 205 3918 233
rect 3115 134 3145 167
rect 2613 73 2643 100
rect 2721 73 2736 107
rect 2792 73 2822 95
rect 2936 73 2966 95
rect 3022 73 3037 107
rect 3115 73 3145 100
rect 3193 134 3223 167
rect 3308 155 3338 177
rect 3580 155 3610 177
rect 4160 205 4190 233
rect 4275 195 4305 217
rect 4353 195 4383 217
rect 4468 205 4498 233
rect 3695 134 3725 167
rect 3193 73 3223 100
rect 3301 73 3316 107
rect 3372 73 3402 95
rect 3516 73 3546 95
rect 3602 73 3617 107
rect 3695 73 3725 100
rect 3773 134 3803 167
rect 3888 155 3918 177
rect 4160 155 4190 177
rect 4740 205 4770 233
rect 4855 195 4885 217
rect 4933 195 4963 217
rect 5048 205 5078 233
rect 4275 134 4305 167
rect 3773 73 3803 100
rect 3881 73 3896 107
rect 3952 73 3982 95
rect 4096 73 4126 95
rect 4182 73 4197 107
rect 4275 73 4305 100
rect 4353 134 4383 167
rect 4468 155 4498 177
rect 4740 155 4770 177
rect 5320 205 5350 233
rect 5435 195 5465 217
rect 5513 195 5543 217
rect 5628 205 5658 233
rect 4855 134 4885 167
rect 4353 73 4383 100
rect 4461 73 4476 107
rect 4532 73 4562 95
rect 4676 73 4706 95
rect 4762 73 4777 107
rect 4855 73 4885 100
rect 4933 134 4963 167
rect 5048 155 5078 177
rect 5320 155 5350 177
rect 5900 205 5930 233
rect 6015 195 6045 217
rect 6093 195 6123 217
rect 6208 205 6238 233
rect 5435 134 5465 167
rect 4933 73 4963 100
rect 5041 73 5056 107
rect 5112 73 5142 95
rect 5256 73 5286 95
rect 5342 73 5357 107
rect 5435 73 5465 100
rect 5513 134 5543 167
rect 5628 155 5658 177
rect 5900 155 5930 177
rect 6480 205 6510 233
rect 6595 195 6625 217
rect 6673 195 6703 217
rect 6788 205 6818 233
rect 6015 134 6045 167
rect 5513 73 5543 100
rect 5621 73 5636 107
rect 5692 73 5722 95
rect 5836 73 5866 95
rect 5922 73 5937 107
rect 6015 73 6045 100
rect 6093 134 6123 167
rect 6208 155 6238 177
rect 6480 155 6510 177
rect 6595 134 6625 167
rect 6093 73 6123 100
rect 6201 73 6216 107
rect 6272 73 6302 95
rect 6416 73 6446 95
rect 6502 73 6517 107
rect 6595 73 6625 100
rect 6673 134 6703 167
rect 6788 155 6818 177
rect 6673 73 6703 100
rect 6781 73 6796 107
rect 6852 73 6882 95
rect 122 59 152 73
rect 386 59 416 73
rect 702 59 732 73
rect 966 59 996 73
rect 1282 59 1312 73
rect 1546 59 1576 73
rect 1862 59 1892 73
rect 2126 59 2156 73
rect 2442 59 2472 73
rect 2706 59 2736 73
rect 3022 59 3052 73
rect 3286 59 3316 73
rect 3602 59 3632 73
rect 3866 59 3896 73
rect 4182 59 4212 73
rect 4446 59 4476 73
rect 4762 59 4792 73
rect 5026 59 5056 73
rect 5342 59 5372 73
rect 5606 59 5636 73
rect 5922 59 5952 73
rect 6186 59 6216 73
rect 6502 59 6532 73
rect 6766 59 6796 73
rect 36 9 66 31
rect 122 9 152 31
rect 215 9 245 31
rect 293 9 323 31
rect 386 9 416 31
rect 472 9 502 31
rect 616 9 646 31
rect 702 9 732 31
rect 795 9 825 31
rect 873 9 903 31
rect 966 9 996 31
rect 1052 9 1082 31
rect 1196 9 1226 31
rect 1282 9 1312 31
rect 1375 9 1405 31
rect 1453 9 1483 31
rect 1546 9 1576 31
rect 1632 9 1662 31
rect 1776 9 1806 31
rect 1862 9 1892 31
rect 1955 9 1985 31
rect 2033 9 2063 31
rect 2126 9 2156 31
rect 2212 9 2242 31
rect 2356 9 2386 31
rect 2442 9 2472 31
rect 2535 9 2565 31
rect 2613 9 2643 31
rect 2706 9 2736 31
rect 2792 9 2822 31
rect 2936 9 2966 31
rect 3022 9 3052 31
rect 3115 9 3145 31
rect 3193 9 3223 31
rect 3286 9 3316 31
rect 3372 9 3402 31
rect 3516 9 3546 31
rect 3602 9 3632 31
rect 3695 9 3725 31
rect 3773 9 3803 31
rect 3866 9 3896 31
rect 3952 9 3982 31
rect 4096 9 4126 31
rect 4182 9 4212 31
rect 4275 9 4305 31
rect 4353 9 4383 31
rect 4446 9 4476 31
rect 4532 9 4562 31
rect 4676 9 4706 31
rect 4762 9 4792 31
rect 4855 9 4885 31
rect 4933 9 4963 31
rect 5026 9 5056 31
rect 5112 9 5142 31
rect 5256 9 5286 31
rect 5342 9 5372 31
rect 5435 9 5465 31
rect 5513 9 5543 31
rect 5606 9 5636 31
rect 5692 9 5722 31
rect 5836 9 5866 31
rect 5922 9 5952 31
rect 6015 9 6045 31
rect 6093 9 6123 31
rect 6186 9 6216 31
rect 6272 9 6302 31
rect 6416 9 6446 31
rect 6502 9 6532 31
rect 6595 9 6625 31
rect 6673 9 6703 31
rect 6766 9 6796 31
rect 6852 9 6882 31
<< polycont >>
rect -91 4283 -43 4313
rect 36 4145 66 4179
rect 137 4123 167 4157
rect 215 4150 245 4184
rect 293 4150 323 4184
rect 371 4123 401 4157
rect 472 4145 502 4179
rect 616 4145 646 4179
rect 717 4123 747 4157
rect 795 4150 825 4184
rect 873 4150 903 4184
rect 951 4123 981 4157
rect 1052 4145 1082 4179
rect 1196 4145 1226 4179
rect 1297 4123 1327 4157
rect 1375 4150 1405 4184
rect 1453 4150 1483 4184
rect 1531 4123 1561 4157
rect 1632 4145 1662 4179
rect 1776 4145 1806 4179
rect 1877 4123 1907 4157
rect 1955 4150 1985 4184
rect 2033 4150 2063 4184
rect 2111 4123 2141 4157
rect 2212 4145 2242 4179
rect 2356 4145 2386 4179
rect 2457 4123 2487 4157
rect 2535 4150 2565 4184
rect 2613 4150 2643 4184
rect 2691 4123 2721 4157
rect 2792 4145 2822 4179
rect 2936 4145 2966 4179
rect 3037 4123 3067 4157
rect 3115 4150 3145 4184
rect 3193 4150 3223 4184
rect 3271 4123 3301 4157
rect 3372 4145 3402 4179
rect 3516 4145 3546 4179
rect 3617 4123 3647 4157
rect 3695 4150 3725 4184
rect 3773 4150 3803 4184
rect 3851 4123 3881 4157
rect 3952 4145 3982 4179
rect 4096 4145 4126 4179
rect 4197 4123 4227 4157
rect 4275 4150 4305 4184
rect 4353 4150 4383 4184
rect 4431 4123 4461 4157
rect 4532 4145 4562 4179
rect 4676 4145 4706 4179
rect 4777 4123 4807 4157
rect 4855 4150 4885 4184
rect 4933 4150 4963 4184
rect 5011 4123 5041 4157
rect 5112 4145 5142 4179
rect 5256 4145 5286 4179
rect 5357 4123 5387 4157
rect 5435 4150 5465 4184
rect 5513 4150 5543 4184
rect 5591 4123 5621 4157
rect 5692 4145 5722 4179
rect 5836 4145 5866 4179
rect 5937 4123 5967 4157
rect 6015 4150 6045 4184
rect 6093 4150 6123 4184
rect 6171 4123 6201 4157
rect 6272 4145 6302 4179
rect 6416 4145 6446 4179
rect 6517 4123 6547 4157
rect 6595 4150 6625 4184
rect 6673 4150 6703 4184
rect 6751 4123 6781 4157
rect 6852 4145 6882 4179
rect -91 4013 -43 4043
rect 36 3875 66 3909
rect 137 3853 167 3887
rect 215 3880 245 3914
rect 293 3880 323 3914
rect 371 3853 401 3887
rect 472 3875 502 3909
rect 616 3875 646 3909
rect 717 3853 747 3887
rect 795 3880 825 3914
rect 873 3880 903 3914
rect 951 3853 981 3887
rect 1052 3875 1082 3909
rect 1196 3875 1226 3909
rect 1297 3853 1327 3887
rect 1375 3880 1405 3914
rect 1453 3880 1483 3914
rect 1531 3853 1561 3887
rect 1632 3875 1662 3909
rect 1776 3875 1806 3909
rect 1877 3853 1907 3887
rect 1955 3880 1985 3914
rect 2033 3880 2063 3914
rect 2111 3853 2141 3887
rect 2212 3875 2242 3909
rect 2356 3875 2386 3909
rect 2457 3853 2487 3887
rect 2535 3880 2565 3914
rect 2613 3880 2643 3914
rect 2691 3853 2721 3887
rect 2792 3875 2822 3909
rect 2936 3875 2966 3909
rect 3037 3853 3067 3887
rect 3115 3880 3145 3914
rect 3193 3880 3223 3914
rect 3271 3853 3301 3887
rect 3372 3875 3402 3909
rect 3516 3875 3546 3909
rect 3617 3853 3647 3887
rect 3695 3880 3725 3914
rect 3773 3880 3803 3914
rect 3851 3853 3881 3887
rect 3952 3875 3982 3909
rect 4096 3875 4126 3909
rect 4197 3853 4227 3887
rect 4275 3880 4305 3914
rect 4353 3880 4383 3914
rect 4431 3853 4461 3887
rect 4532 3875 4562 3909
rect 4676 3875 4706 3909
rect 4777 3853 4807 3887
rect 4855 3880 4885 3914
rect 4933 3880 4963 3914
rect 5011 3853 5041 3887
rect 5112 3875 5142 3909
rect 5256 3875 5286 3909
rect 5357 3853 5387 3887
rect 5435 3880 5465 3914
rect 5513 3880 5543 3914
rect 5591 3853 5621 3887
rect 5692 3875 5722 3909
rect 5836 3875 5866 3909
rect 5937 3853 5967 3887
rect 6015 3880 6045 3914
rect 6093 3880 6123 3914
rect 6171 3853 6201 3887
rect 6272 3875 6302 3909
rect 6416 3875 6446 3909
rect 6517 3853 6547 3887
rect 6595 3880 6625 3914
rect 6673 3880 6703 3914
rect 6751 3853 6781 3887
rect 6852 3875 6882 3909
rect -91 3743 -43 3773
rect 36 3605 66 3639
rect 137 3583 167 3617
rect 215 3610 245 3644
rect 293 3610 323 3644
rect 371 3583 401 3617
rect 472 3605 502 3639
rect 616 3605 646 3639
rect 717 3583 747 3617
rect 795 3610 825 3644
rect 873 3610 903 3644
rect 951 3583 981 3617
rect 1052 3605 1082 3639
rect 1196 3605 1226 3639
rect 1297 3583 1327 3617
rect 1375 3610 1405 3644
rect 1453 3610 1483 3644
rect 1531 3583 1561 3617
rect 1632 3605 1662 3639
rect 1776 3605 1806 3639
rect 1877 3583 1907 3617
rect 1955 3610 1985 3644
rect 2033 3610 2063 3644
rect 2111 3583 2141 3617
rect 2212 3605 2242 3639
rect 2356 3605 2386 3639
rect 2457 3583 2487 3617
rect 2535 3610 2565 3644
rect 2613 3610 2643 3644
rect 2691 3583 2721 3617
rect 2792 3605 2822 3639
rect 2936 3605 2966 3639
rect 3037 3583 3067 3617
rect 3115 3610 3145 3644
rect 3193 3610 3223 3644
rect 3271 3583 3301 3617
rect 3372 3605 3402 3639
rect 3516 3605 3546 3639
rect 3617 3583 3647 3617
rect 3695 3610 3725 3644
rect 3773 3610 3803 3644
rect 3851 3583 3881 3617
rect 3952 3605 3982 3639
rect 4096 3605 4126 3639
rect 4197 3583 4227 3617
rect 4275 3610 4305 3644
rect 4353 3610 4383 3644
rect 4431 3583 4461 3617
rect 4532 3605 4562 3639
rect 4676 3605 4706 3639
rect 4777 3583 4807 3617
rect 4855 3610 4885 3644
rect 4933 3610 4963 3644
rect 5011 3583 5041 3617
rect 5112 3605 5142 3639
rect 5256 3605 5286 3639
rect 5357 3583 5387 3617
rect 5435 3610 5465 3644
rect 5513 3610 5543 3644
rect 5591 3583 5621 3617
rect 5692 3605 5722 3639
rect 5836 3605 5866 3639
rect 5937 3583 5967 3617
rect 6015 3610 6045 3644
rect 6093 3610 6123 3644
rect 6171 3583 6201 3617
rect 6272 3605 6302 3639
rect 6416 3605 6446 3639
rect 6517 3583 6547 3617
rect 6595 3610 6625 3644
rect 6673 3610 6703 3644
rect 6751 3583 6781 3617
rect 6852 3605 6882 3639
rect -91 3473 -43 3503
rect 36 3335 66 3369
rect 137 3313 167 3347
rect 215 3340 245 3374
rect 293 3340 323 3374
rect 371 3313 401 3347
rect 472 3335 502 3369
rect 616 3335 646 3369
rect 717 3313 747 3347
rect 795 3340 825 3374
rect 873 3340 903 3374
rect 951 3313 981 3347
rect 1052 3335 1082 3369
rect 1196 3335 1226 3369
rect 1297 3313 1327 3347
rect 1375 3340 1405 3374
rect 1453 3340 1483 3374
rect 1531 3313 1561 3347
rect 1632 3335 1662 3369
rect 1776 3335 1806 3369
rect 1877 3313 1907 3347
rect 1955 3340 1985 3374
rect 2033 3340 2063 3374
rect 2111 3313 2141 3347
rect 2212 3335 2242 3369
rect 2356 3335 2386 3369
rect 2457 3313 2487 3347
rect 2535 3340 2565 3374
rect 2613 3340 2643 3374
rect 2691 3313 2721 3347
rect 2792 3335 2822 3369
rect 2936 3335 2966 3369
rect 3037 3313 3067 3347
rect 3115 3340 3145 3374
rect 3193 3340 3223 3374
rect 3271 3313 3301 3347
rect 3372 3335 3402 3369
rect 3516 3335 3546 3369
rect 3617 3313 3647 3347
rect 3695 3340 3725 3374
rect 3773 3340 3803 3374
rect 3851 3313 3881 3347
rect 3952 3335 3982 3369
rect 4096 3335 4126 3369
rect 4197 3313 4227 3347
rect 4275 3340 4305 3374
rect 4353 3340 4383 3374
rect 4431 3313 4461 3347
rect 4532 3335 4562 3369
rect 4676 3335 4706 3369
rect 4777 3313 4807 3347
rect 4855 3340 4885 3374
rect 4933 3340 4963 3374
rect 5011 3313 5041 3347
rect 5112 3335 5142 3369
rect 5256 3335 5286 3369
rect 5357 3313 5387 3347
rect 5435 3340 5465 3374
rect 5513 3340 5543 3374
rect 5591 3313 5621 3347
rect 5692 3335 5722 3369
rect 5836 3335 5866 3369
rect 5937 3313 5967 3347
rect 6015 3340 6045 3374
rect 6093 3340 6123 3374
rect 6171 3313 6201 3347
rect 6272 3335 6302 3369
rect 6416 3335 6446 3369
rect 6517 3313 6547 3347
rect 6595 3340 6625 3374
rect 6673 3340 6703 3374
rect 6751 3313 6781 3347
rect 6852 3335 6882 3369
rect -91 3203 -43 3233
rect 36 3065 66 3099
rect 137 3043 167 3077
rect 215 3070 245 3104
rect 293 3070 323 3104
rect 371 3043 401 3077
rect 472 3065 502 3099
rect 616 3065 646 3099
rect 717 3043 747 3077
rect 795 3070 825 3104
rect 873 3070 903 3104
rect 951 3043 981 3077
rect 1052 3065 1082 3099
rect 1196 3065 1226 3099
rect 1297 3043 1327 3077
rect 1375 3070 1405 3104
rect 1453 3070 1483 3104
rect 1531 3043 1561 3077
rect 1632 3065 1662 3099
rect 1776 3065 1806 3099
rect 1877 3043 1907 3077
rect 1955 3070 1985 3104
rect 2033 3070 2063 3104
rect 2111 3043 2141 3077
rect 2212 3065 2242 3099
rect 2356 3065 2386 3099
rect 2457 3043 2487 3077
rect 2535 3070 2565 3104
rect 2613 3070 2643 3104
rect 2691 3043 2721 3077
rect 2792 3065 2822 3099
rect 2936 3065 2966 3099
rect 3037 3043 3067 3077
rect 3115 3070 3145 3104
rect 3193 3070 3223 3104
rect 3271 3043 3301 3077
rect 3372 3065 3402 3099
rect 3516 3065 3546 3099
rect 3617 3043 3647 3077
rect 3695 3070 3725 3104
rect 3773 3070 3803 3104
rect 3851 3043 3881 3077
rect 3952 3065 3982 3099
rect 4096 3065 4126 3099
rect 4197 3043 4227 3077
rect 4275 3070 4305 3104
rect 4353 3070 4383 3104
rect 4431 3043 4461 3077
rect 4532 3065 4562 3099
rect 4676 3065 4706 3099
rect 4777 3043 4807 3077
rect 4855 3070 4885 3104
rect 4933 3070 4963 3104
rect 5011 3043 5041 3077
rect 5112 3065 5142 3099
rect 5256 3065 5286 3099
rect 5357 3043 5387 3077
rect 5435 3070 5465 3104
rect 5513 3070 5543 3104
rect 5591 3043 5621 3077
rect 5692 3065 5722 3099
rect 5836 3065 5866 3099
rect 5937 3043 5967 3077
rect 6015 3070 6045 3104
rect 6093 3070 6123 3104
rect 6171 3043 6201 3077
rect 6272 3065 6302 3099
rect 6416 3065 6446 3099
rect 6517 3043 6547 3077
rect 6595 3070 6625 3104
rect 6673 3070 6703 3104
rect 6751 3043 6781 3077
rect 6852 3065 6882 3099
rect -91 2933 -43 2963
rect 36 2795 66 2829
rect 137 2773 167 2807
rect 215 2800 245 2834
rect 293 2800 323 2834
rect 371 2773 401 2807
rect 472 2795 502 2829
rect 616 2795 646 2829
rect 717 2773 747 2807
rect 795 2800 825 2834
rect 873 2800 903 2834
rect 951 2773 981 2807
rect 1052 2795 1082 2829
rect 1196 2795 1226 2829
rect 1297 2773 1327 2807
rect 1375 2800 1405 2834
rect 1453 2800 1483 2834
rect 1531 2773 1561 2807
rect 1632 2795 1662 2829
rect 1776 2795 1806 2829
rect 1877 2773 1907 2807
rect 1955 2800 1985 2834
rect 2033 2800 2063 2834
rect 2111 2773 2141 2807
rect 2212 2795 2242 2829
rect 2356 2795 2386 2829
rect 2457 2773 2487 2807
rect 2535 2800 2565 2834
rect 2613 2800 2643 2834
rect 2691 2773 2721 2807
rect 2792 2795 2822 2829
rect 2936 2795 2966 2829
rect 3037 2773 3067 2807
rect 3115 2800 3145 2834
rect 3193 2800 3223 2834
rect 3271 2773 3301 2807
rect 3372 2795 3402 2829
rect 3516 2795 3546 2829
rect 3617 2773 3647 2807
rect 3695 2800 3725 2834
rect 3773 2800 3803 2834
rect 3851 2773 3881 2807
rect 3952 2795 3982 2829
rect 4096 2795 4126 2829
rect 4197 2773 4227 2807
rect 4275 2800 4305 2834
rect 4353 2800 4383 2834
rect 4431 2773 4461 2807
rect 4532 2795 4562 2829
rect 4676 2795 4706 2829
rect 4777 2773 4807 2807
rect 4855 2800 4885 2834
rect 4933 2800 4963 2834
rect 5011 2773 5041 2807
rect 5112 2795 5142 2829
rect 5256 2795 5286 2829
rect 5357 2773 5387 2807
rect 5435 2800 5465 2834
rect 5513 2800 5543 2834
rect 5591 2773 5621 2807
rect 5692 2795 5722 2829
rect 5836 2795 5866 2829
rect 5937 2773 5967 2807
rect 6015 2800 6045 2834
rect 6093 2800 6123 2834
rect 6171 2773 6201 2807
rect 6272 2795 6302 2829
rect 6416 2795 6446 2829
rect 6517 2773 6547 2807
rect 6595 2800 6625 2834
rect 6673 2800 6703 2834
rect 6751 2773 6781 2807
rect 6852 2795 6882 2829
rect -91 2663 -43 2693
rect 36 2525 66 2559
rect 137 2503 167 2537
rect 215 2530 245 2564
rect 293 2530 323 2564
rect 371 2503 401 2537
rect 472 2525 502 2559
rect 616 2525 646 2559
rect 717 2503 747 2537
rect 795 2530 825 2564
rect 873 2530 903 2564
rect 951 2503 981 2537
rect 1052 2525 1082 2559
rect 1196 2525 1226 2559
rect 1297 2503 1327 2537
rect 1375 2530 1405 2564
rect 1453 2530 1483 2564
rect 1531 2503 1561 2537
rect 1632 2525 1662 2559
rect 1776 2525 1806 2559
rect 1877 2503 1907 2537
rect 1955 2530 1985 2564
rect 2033 2530 2063 2564
rect 2111 2503 2141 2537
rect 2212 2525 2242 2559
rect 2356 2525 2386 2559
rect 2457 2503 2487 2537
rect 2535 2530 2565 2564
rect 2613 2530 2643 2564
rect 2691 2503 2721 2537
rect 2792 2525 2822 2559
rect 2936 2525 2966 2559
rect 3037 2503 3067 2537
rect 3115 2530 3145 2564
rect 3193 2530 3223 2564
rect 3271 2503 3301 2537
rect 3372 2525 3402 2559
rect 3516 2525 3546 2559
rect 3617 2503 3647 2537
rect 3695 2530 3725 2564
rect 3773 2530 3803 2564
rect 3851 2503 3881 2537
rect 3952 2525 3982 2559
rect 4096 2525 4126 2559
rect 4197 2503 4227 2537
rect 4275 2530 4305 2564
rect 4353 2530 4383 2564
rect 4431 2503 4461 2537
rect 4532 2525 4562 2559
rect 4676 2525 4706 2559
rect 4777 2503 4807 2537
rect 4855 2530 4885 2564
rect 4933 2530 4963 2564
rect 5011 2503 5041 2537
rect 5112 2525 5142 2559
rect 5256 2525 5286 2559
rect 5357 2503 5387 2537
rect 5435 2530 5465 2564
rect 5513 2530 5543 2564
rect 5591 2503 5621 2537
rect 5692 2525 5722 2559
rect 5836 2525 5866 2559
rect 5937 2503 5967 2537
rect 6015 2530 6045 2564
rect 6093 2530 6123 2564
rect 6171 2503 6201 2537
rect 6272 2525 6302 2559
rect 6416 2525 6446 2559
rect 6517 2503 6547 2537
rect 6595 2530 6625 2564
rect 6673 2530 6703 2564
rect 6751 2503 6781 2537
rect 6852 2525 6882 2559
rect -91 2393 -43 2423
rect 36 2255 66 2289
rect 137 2233 167 2267
rect 215 2260 245 2294
rect 293 2260 323 2294
rect 371 2233 401 2267
rect 472 2255 502 2289
rect 616 2255 646 2289
rect 717 2233 747 2267
rect 795 2260 825 2294
rect 873 2260 903 2294
rect 951 2233 981 2267
rect 1052 2255 1082 2289
rect 1196 2255 1226 2289
rect 1297 2233 1327 2267
rect 1375 2260 1405 2294
rect 1453 2260 1483 2294
rect 1531 2233 1561 2267
rect 1632 2255 1662 2289
rect 1776 2255 1806 2289
rect 1877 2233 1907 2267
rect 1955 2260 1985 2294
rect 2033 2260 2063 2294
rect 2111 2233 2141 2267
rect 2212 2255 2242 2289
rect 2356 2255 2386 2289
rect 2457 2233 2487 2267
rect 2535 2260 2565 2294
rect 2613 2260 2643 2294
rect 2691 2233 2721 2267
rect 2792 2255 2822 2289
rect 2936 2255 2966 2289
rect 3037 2233 3067 2267
rect 3115 2260 3145 2294
rect 3193 2260 3223 2294
rect 3271 2233 3301 2267
rect 3372 2255 3402 2289
rect 3516 2255 3546 2289
rect 3617 2233 3647 2267
rect 3695 2260 3725 2294
rect 3773 2260 3803 2294
rect 3851 2233 3881 2267
rect 3952 2255 3982 2289
rect 4096 2255 4126 2289
rect 4197 2233 4227 2267
rect 4275 2260 4305 2294
rect 4353 2260 4383 2294
rect 4431 2233 4461 2267
rect 4532 2255 4562 2289
rect 4676 2255 4706 2289
rect 4777 2233 4807 2267
rect 4855 2260 4885 2294
rect 4933 2260 4963 2294
rect 5011 2233 5041 2267
rect 5112 2255 5142 2289
rect 5256 2255 5286 2289
rect 5357 2233 5387 2267
rect 5435 2260 5465 2294
rect 5513 2260 5543 2294
rect 5591 2233 5621 2267
rect 5692 2255 5722 2289
rect 5836 2255 5866 2289
rect 5937 2233 5967 2267
rect 6015 2260 6045 2294
rect 6093 2260 6123 2294
rect 6171 2233 6201 2267
rect 6272 2255 6302 2289
rect 6416 2255 6446 2289
rect 6517 2233 6547 2267
rect 6595 2260 6625 2294
rect 6673 2260 6703 2294
rect 6751 2233 6781 2267
rect 6852 2255 6882 2289
rect -91 2123 -43 2153
rect 36 1985 66 2019
rect 137 1963 167 1997
rect 215 1990 245 2024
rect 293 1990 323 2024
rect 371 1963 401 1997
rect 472 1985 502 2019
rect 616 1985 646 2019
rect 717 1963 747 1997
rect 795 1990 825 2024
rect 873 1990 903 2024
rect 951 1963 981 1997
rect 1052 1985 1082 2019
rect 1196 1985 1226 2019
rect 1297 1963 1327 1997
rect 1375 1990 1405 2024
rect 1453 1990 1483 2024
rect 1531 1963 1561 1997
rect 1632 1985 1662 2019
rect 1776 1985 1806 2019
rect 1877 1963 1907 1997
rect 1955 1990 1985 2024
rect 2033 1990 2063 2024
rect 2111 1963 2141 1997
rect 2212 1985 2242 2019
rect 2356 1985 2386 2019
rect 2457 1963 2487 1997
rect 2535 1990 2565 2024
rect 2613 1990 2643 2024
rect 2691 1963 2721 1997
rect 2792 1985 2822 2019
rect 2936 1985 2966 2019
rect 3037 1963 3067 1997
rect 3115 1990 3145 2024
rect 3193 1990 3223 2024
rect 3271 1963 3301 1997
rect 3372 1985 3402 2019
rect 3516 1985 3546 2019
rect 3617 1963 3647 1997
rect 3695 1990 3725 2024
rect 3773 1990 3803 2024
rect 3851 1963 3881 1997
rect 3952 1985 3982 2019
rect 4096 1985 4126 2019
rect 4197 1963 4227 1997
rect 4275 1990 4305 2024
rect 4353 1990 4383 2024
rect 4431 1963 4461 1997
rect 4532 1985 4562 2019
rect 4676 1985 4706 2019
rect 4777 1963 4807 1997
rect 4855 1990 4885 2024
rect 4933 1990 4963 2024
rect 5011 1963 5041 1997
rect 5112 1985 5142 2019
rect 5256 1985 5286 2019
rect 5357 1963 5387 1997
rect 5435 1990 5465 2024
rect 5513 1990 5543 2024
rect 5591 1963 5621 1997
rect 5692 1985 5722 2019
rect 5836 1985 5866 2019
rect 5937 1963 5967 1997
rect 6015 1990 6045 2024
rect 6093 1990 6123 2024
rect 6171 1963 6201 1997
rect 6272 1985 6302 2019
rect 6416 1985 6446 2019
rect 6517 1963 6547 1997
rect 6595 1990 6625 2024
rect 6673 1990 6703 2024
rect 6751 1963 6781 1997
rect 6852 1985 6882 2019
rect -91 1853 -43 1883
rect 36 1715 66 1749
rect 137 1693 167 1727
rect 215 1720 245 1754
rect 293 1720 323 1754
rect 371 1693 401 1727
rect 472 1715 502 1749
rect 616 1715 646 1749
rect 717 1693 747 1727
rect 795 1720 825 1754
rect 873 1720 903 1754
rect 951 1693 981 1727
rect 1052 1715 1082 1749
rect 1196 1715 1226 1749
rect 1297 1693 1327 1727
rect 1375 1720 1405 1754
rect 1453 1720 1483 1754
rect 1531 1693 1561 1727
rect 1632 1715 1662 1749
rect 1776 1715 1806 1749
rect 1877 1693 1907 1727
rect 1955 1720 1985 1754
rect 2033 1720 2063 1754
rect 2111 1693 2141 1727
rect 2212 1715 2242 1749
rect 2356 1715 2386 1749
rect 2457 1693 2487 1727
rect 2535 1720 2565 1754
rect 2613 1720 2643 1754
rect 2691 1693 2721 1727
rect 2792 1715 2822 1749
rect 2936 1715 2966 1749
rect 3037 1693 3067 1727
rect 3115 1720 3145 1754
rect 3193 1720 3223 1754
rect 3271 1693 3301 1727
rect 3372 1715 3402 1749
rect 3516 1715 3546 1749
rect 3617 1693 3647 1727
rect 3695 1720 3725 1754
rect 3773 1720 3803 1754
rect 3851 1693 3881 1727
rect 3952 1715 3982 1749
rect 4096 1715 4126 1749
rect 4197 1693 4227 1727
rect 4275 1720 4305 1754
rect 4353 1720 4383 1754
rect 4431 1693 4461 1727
rect 4532 1715 4562 1749
rect 4676 1715 4706 1749
rect 4777 1693 4807 1727
rect 4855 1720 4885 1754
rect 4933 1720 4963 1754
rect 5011 1693 5041 1727
rect 5112 1715 5142 1749
rect 5256 1715 5286 1749
rect 5357 1693 5387 1727
rect 5435 1720 5465 1754
rect 5513 1720 5543 1754
rect 5591 1693 5621 1727
rect 5692 1715 5722 1749
rect 5836 1715 5866 1749
rect 5937 1693 5967 1727
rect 6015 1720 6045 1754
rect 6093 1720 6123 1754
rect 6171 1693 6201 1727
rect 6272 1715 6302 1749
rect 6416 1715 6446 1749
rect 6517 1693 6547 1727
rect 6595 1720 6625 1754
rect 6673 1720 6703 1754
rect 6751 1693 6781 1727
rect 6852 1715 6882 1749
rect -91 1583 -43 1613
rect 36 1445 66 1479
rect 137 1423 167 1457
rect 215 1450 245 1484
rect 293 1450 323 1484
rect 371 1423 401 1457
rect 472 1445 502 1479
rect 616 1445 646 1479
rect 717 1423 747 1457
rect 795 1450 825 1484
rect 873 1450 903 1484
rect 951 1423 981 1457
rect 1052 1445 1082 1479
rect 1196 1445 1226 1479
rect 1297 1423 1327 1457
rect 1375 1450 1405 1484
rect 1453 1450 1483 1484
rect 1531 1423 1561 1457
rect 1632 1445 1662 1479
rect 1776 1445 1806 1479
rect 1877 1423 1907 1457
rect 1955 1450 1985 1484
rect 2033 1450 2063 1484
rect 2111 1423 2141 1457
rect 2212 1445 2242 1479
rect 2356 1445 2386 1479
rect 2457 1423 2487 1457
rect 2535 1450 2565 1484
rect 2613 1450 2643 1484
rect 2691 1423 2721 1457
rect 2792 1445 2822 1479
rect 2936 1445 2966 1479
rect 3037 1423 3067 1457
rect 3115 1450 3145 1484
rect 3193 1450 3223 1484
rect 3271 1423 3301 1457
rect 3372 1445 3402 1479
rect 3516 1445 3546 1479
rect 3617 1423 3647 1457
rect 3695 1450 3725 1484
rect 3773 1450 3803 1484
rect 3851 1423 3881 1457
rect 3952 1445 3982 1479
rect 4096 1445 4126 1479
rect 4197 1423 4227 1457
rect 4275 1450 4305 1484
rect 4353 1450 4383 1484
rect 4431 1423 4461 1457
rect 4532 1445 4562 1479
rect 4676 1445 4706 1479
rect 4777 1423 4807 1457
rect 4855 1450 4885 1484
rect 4933 1450 4963 1484
rect 5011 1423 5041 1457
rect 5112 1445 5142 1479
rect 5256 1445 5286 1479
rect 5357 1423 5387 1457
rect 5435 1450 5465 1484
rect 5513 1450 5543 1484
rect 5591 1423 5621 1457
rect 5692 1445 5722 1479
rect 5836 1445 5866 1479
rect 5937 1423 5967 1457
rect 6015 1450 6045 1484
rect 6093 1450 6123 1484
rect 6171 1423 6201 1457
rect 6272 1445 6302 1479
rect 6416 1445 6446 1479
rect 6517 1423 6547 1457
rect 6595 1450 6625 1484
rect 6673 1450 6703 1484
rect 6751 1423 6781 1457
rect 6852 1445 6882 1479
rect -91 1313 -43 1343
rect 36 1175 66 1209
rect 137 1153 167 1187
rect 215 1180 245 1214
rect 293 1180 323 1214
rect 371 1153 401 1187
rect 472 1175 502 1209
rect 616 1175 646 1209
rect 717 1153 747 1187
rect 795 1180 825 1214
rect 873 1180 903 1214
rect 951 1153 981 1187
rect 1052 1175 1082 1209
rect 1196 1175 1226 1209
rect 1297 1153 1327 1187
rect 1375 1180 1405 1214
rect 1453 1180 1483 1214
rect 1531 1153 1561 1187
rect 1632 1175 1662 1209
rect 1776 1175 1806 1209
rect 1877 1153 1907 1187
rect 1955 1180 1985 1214
rect 2033 1180 2063 1214
rect 2111 1153 2141 1187
rect 2212 1175 2242 1209
rect 2356 1175 2386 1209
rect 2457 1153 2487 1187
rect 2535 1180 2565 1214
rect 2613 1180 2643 1214
rect 2691 1153 2721 1187
rect 2792 1175 2822 1209
rect 2936 1175 2966 1209
rect 3037 1153 3067 1187
rect 3115 1180 3145 1214
rect 3193 1180 3223 1214
rect 3271 1153 3301 1187
rect 3372 1175 3402 1209
rect 3516 1175 3546 1209
rect 3617 1153 3647 1187
rect 3695 1180 3725 1214
rect 3773 1180 3803 1214
rect 3851 1153 3881 1187
rect 3952 1175 3982 1209
rect 4096 1175 4126 1209
rect 4197 1153 4227 1187
rect 4275 1180 4305 1214
rect 4353 1180 4383 1214
rect 4431 1153 4461 1187
rect 4532 1175 4562 1209
rect 4676 1175 4706 1209
rect 4777 1153 4807 1187
rect 4855 1180 4885 1214
rect 4933 1180 4963 1214
rect 5011 1153 5041 1187
rect 5112 1175 5142 1209
rect 5256 1175 5286 1209
rect 5357 1153 5387 1187
rect 5435 1180 5465 1214
rect 5513 1180 5543 1214
rect 5591 1153 5621 1187
rect 5692 1175 5722 1209
rect 5836 1175 5866 1209
rect 5937 1153 5967 1187
rect 6015 1180 6045 1214
rect 6093 1180 6123 1214
rect 6171 1153 6201 1187
rect 6272 1175 6302 1209
rect 6416 1175 6446 1209
rect 6517 1153 6547 1187
rect 6595 1180 6625 1214
rect 6673 1180 6703 1214
rect 6751 1153 6781 1187
rect 6852 1175 6882 1209
rect -91 1043 -43 1073
rect 36 905 66 939
rect 137 883 167 917
rect 215 910 245 944
rect 293 910 323 944
rect 371 883 401 917
rect 472 905 502 939
rect 616 905 646 939
rect 717 883 747 917
rect 795 910 825 944
rect 873 910 903 944
rect 951 883 981 917
rect 1052 905 1082 939
rect 1196 905 1226 939
rect 1297 883 1327 917
rect 1375 910 1405 944
rect 1453 910 1483 944
rect 1531 883 1561 917
rect 1632 905 1662 939
rect 1776 905 1806 939
rect 1877 883 1907 917
rect 1955 910 1985 944
rect 2033 910 2063 944
rect 2111 883 2141 917
rect 2212 905 2242 939
rect 2356 905 2386 939
rect 2457 883 2487 917
rect 2535 910 2565 944
rect 2613 910 2643 944
rect 2691 883 2721 917
rect 2792 905 2822 939
rect 2936 905 2966 939
rect 3037 883 3067 917
rect 3115 910 3145 944
rect 3193 910 3223 944
rect 3271 883 3301 917
rect 3372 905 3402 939
rect 3516 905 3546 939
rect 3617 883 3647 917
rect 3695 910 3725 944
rect 3773 910 3803 944
rect 3851 883 3881 917
rect 3952 905 3982 939
rect 4096 905 4126 939
rect 4197 883 4227 917
rect 4275 910 4305 944
rect 4353 910 4383 944
rect 4431 883 4461 917
rect 4532 905 4562 939
rect 4676 905 4706 939
rect 4777 883 4807 917
rect 4855 910 4885 944
rect 4933 910 4963 944
rect 5011 883 5041 917
rect 5112 905 5142 939
rect 5256 905 5286 939
rect 5357 883 5387 917
rect 5435 910 5465 944
rect 5513 910 5543 944
rect 5591 883 5621 917
rect 5692 905 5722 939
rect 5836 905 5866 939
rect 5937 883 5967 917
rect 6015 910 6045 944
rect 6093 910 6123 944
rect 6171 883 6201 917
rect 6272 905 6302 939
rect 6416 905 6446 939
rect 6517 883 6547 917
rect 6595 910 6625 944
rect 6673 910 6703 944
rect 6751 883 6781 917
rect 6852 905 6882 939
rect -91 773 -43 803
rect 36 635 66 669
rect 137 613 167 647
rect 215 640 245 674
rect 293 640 323 674
rect 371 613 401 647
rect 472 635 502 669
rect 616 635 646 669
rect 717 613 747 647
rect 795 640 825 674
rect 873 640 903 674
rect 951 613 981 647
rect 1052 635 1082 669
rect 1196 635 1226 669
rect 1297 613 1327 647
rect 1375 640 1405 674
rect 1453 640 1483 674
rect 1531 613 1561 647
rect 1632 635 1662 669
rect 1776 635 1806 669
rect 1877 613 1907 647
rect 1955 640 1985 674
rect 2033 640 2063 674
rect 2111 613 2141 647
rect 2212 635 2242 669
rect 2356 635 2386 669
rect 2457 613 2487 647
rect 2535 640 2565 674
rect 2613 640 2643 674
rect 2691 613 2721 647
rect 2792 635 2822 669
rect 2936 635 2966 669
rect 3037 613 3067 647
rect 3115 640 3145 674
rect 3193 640 3223 674
rect 3271 613 3301 647
rect 3372 635 3402 669
rect 3516 635 3546 669
rect 3617 613 3647 647
rect 3695 640 3725 674
rect 3773 640 3803 674
rect 3851 613 3881 647
rect 3952 635 3982 669
rect 4096 635 4126 669
rect 4197 613 4227 647
rect 4275 640 4305 674
rect 4353 640 4383 674
rect 4431 613 4461 647
rect 4532 635 4562 669
rect 4676 635 4706 669
rect 4777 613 4807 647
rect 4855 640 4885 674
rect 4933 640 4963 674
rect 5011 613 5041 647
rect 5112 635 5142 669
rect 5256 635 5286 669
rect 5357 613 5387 647
rect 5435 640 5465 674
rect 5513 640 5543 674
rect 5591 613 5621 647
rect 5692 635 5722 669
rect 5836 635 5866 669
rect 5937 613 5967 647
rect 6015 640 6045 674
rect 6093 640 6123 674
rect 6171 613 6201 647
rect 6272 635 6302 669
rect 6416 635 6446 669
rect 6517 613 6547 647
rect 6595 640 6625 674
rect 6673 640 6703 674
rect 6751 613 6781 647
rect 6852 635 6882 669
rect -91 503 -43 533
rect 36 365 66 399
rect 137 343 167 377
rect 215 370 245 404
rect 293 370 323 404
rect 371 343 401 377
rect 472 365 502 399
rect 616 365 646 399
rect 717 343 747 377
rect 795 370 825 404
rect 873 370 903 404
rect 951 343 981 377
rect 1052 365 1082 399
rect 1196 365 1226 399
rect 1297 343 1327 377
rect 1375 370 1405 404
rect 1453 370 1483 404
rect 1531 343 1561 377
rect 1632 365 1662 399
rect 1776 365 1806 399
rect 1877 343 1907 377
rect 1955 370 1985 404
rect 2033 370 2063 404
rect 2111 343 2141 377
rect 2212 365 2242 399
rect 2356 365 2386 399
rect 2457 343 2487 377
rect 2535 370 2565 404
rect 2613 370 2643 404
rect 2691 343 2721 377
rect 2792 365 2822 399
rect 2936 365 2966 399
rect 3037 343 3067 377
rect 3115 370 3145 404
rect 3193 370 3223 404
rect 3271 343 3301 377
rect 3372 365 3402 399
rect 3516 365 3546 399
rect 3617 343 3647 377
rect 3695 370 3725 404
rect 3773 370 3803 404
rect 3851 343 3881 377
rect 3952 365 3982 399
rect 4096 365 4126 399
rect 4197 343 4227 377
rect 4275 370 4305 404
rect 4353 370 4383 404
rect 4431 343 4461 377
rect 4532 365 4562 399
rect 4676 365 4706 399
rect 4777 343 4807 377
rect 4855 370 4885 404
rect 4933 370 4963 404
rect 5011 343 5041 377
rect 5112 365 5142 399
rect 5256 365 5286 399
rect 5357 343 5387 377
rect 5435 370 5465 404
rect 5513 370 5543 404
rect 5591 343 5621 377
rect 5692 365 5722 399
rect 5836 365 5866 399
rect 5937 343 5967 377
rect 6015 370 6045 404
rect 6093 370 6123 404
rect 6171 343 6201 377
rect 6272 365 6302 399
rect 6416 365 6446 399
rect 6517 343 6547 377
rect 6595 370 6625 404
rect 6673 370 6703 404
rect 6751 343 6781 377
rect 6852 365 6882 399
rect -91 233 -43 263
rect 36 95 66 129
rect 137 73 167 107
rect 215 100 245 134
rect 293 100 323 134
rect 371 73 401 107
rect 472 95 502 129
rect 616 95 646 129
rect 717 73 747 107
rect 795 100 825 134
rect 873 100 903 134
rect 951 73 981 107
rect 1052 95 1082 129
rect 1196 95 1226 129
rect 1297 73 1327 107
rect 1375 100 1405 134
rect 1453 100 1483 134
rect 1531 73 1561 107
rect 1632 95 1662 129
rect 1776 95 1806 129
rect 1877 73 1907 107
rect 1955 100 1985 134
rect 2033 100 2063 134
rect 2111 73 2141 107
rect 2212 95 2242 129
rect 2356 95 2386 129
rect 2457 73 2487 107
rect 2535 100 2565 134
rect 2613 100 2643 134
rect 2691 73 2721 107
rect 2792 95 2822 129
rect 2936 95 2966 129
rect 3037 73 3067 107
rect 3115 100 3145 134
rect 3193 100 3223 134
rect 3271 73 3301 107
rect 3372 95 3402 129
rect 3516 95 3546 129
rect 3617 73 3647 107
rect 3695 100 3725 134
rect 3773 100 3803 134
rect 3851 73 3881 107
rect 3952 95 3982 129
rect 4096 95 4126 129
rect 4197 73 4227 107
rect 4275 100 4305 134
rect 4353 100 4383 134
rect 4431 73 4461 107
rect 4532 95 4562 129
rect 4676 95 4706 129
rect 4777 73 4807 107
rect 4855 100 4885 134
rect 4933 100 4963 134
rect 5011 73 5041 107
rect 5112 95 5142 129
rect 5256 95 5286 129
rect 5357 73 5387 107
rect 5435 100 5465 134
rect 5513 100 5543 134
rect 5591 73 5621 107
rect 5692 95 5722 129
rect 5836 95 5866 129
rect 5937 73 5967 107
rect 6015 100 6045 134
rect 6093 100 6123 134
rect 6171 73 6201 107
rect 6272 95 6302 129
rect 6416 95 6446 129
rect 6517 73 6547 107
rect 6595 100 6625 134
rect 6673 100 6703 134
rect 6751 73 6781 107
rect 6852 95 6882 129
<< corelocali >>
rect -7 4123 8 4361
tri 73 4277 95 4299 se
rect 95 4292 110 4361
tri 95 4277 110 4292 nw
rect 429 4292 444 4362
tri 67 4271 73 4277 se
rect 73 4271 82 4277
rect 67 4255 82 4271
tri 82 4264 95 4277 nw
rect 236 4269 253 4283
rect 285 4269 302 4283
tri 429 4277 444 4292 ne
tri 444 4277 466 4299 sw
rect 67 4219 82 4227
rect 148 4255 208 4269
rect 163 4245 208 4255
rect 163 4227 191 4245
tri 67 4204 82 4219 ne
tri 82 4204 104 4226 sw
rect 148 4217 191 4227
rect 206 4241 208 4245
rect 330 4255 390 4269
tri 444 4264 457 4277 ne
rect 457 4271 466 4277
tri 466 4271 472 4277 sw
rect 330 4245 375 4255
rect 206 4217 280 4241
rect 148 4213 280 4217
tri 280 4213 308 4241 sw
rect 330 4231 332 4245
tri 330 4229 332 4231 ne
rect 344 4227 375 4245
rect 344 4217 390 4227
rect 457 4256 472 4271
tri 82 4192 94 4204 ne
rect 94 4199 104 4204
tri 104 4199 109 4204 sw
rect -7 3853 8 4081
rect 94 4043 109 4199
rect 148 4157 176 4213
tri 268 4195 286 4213 ne
rect 286 4193 308 4213
tri 308 4193 328 4213 sw
tri 344 4199 362 4217 ne
rect 167 4123 176 4157
rect 210 4184 252 4185
rect 210 4150 215 4184
rect 245 4150 252 4184
rect 210 4141 252 4150
rect 286 4184 328 4193
rect 286 4150 293 4184
rect 323 4150 328 4184
rect 286 4145 328 4150
rect 362 4157 390 4217
tri 435 4204 457 4226 se
rect 457 4219 472 4227
tri 457 4204 472 4219 nw
tri 429 4198 435 4204 se
rect 435 4198 444 4204
rect 148 4113 176 4123
tri 176 4113 200 4137 sw
rect 148 4081 190 4113
tri 207 4105 208 4106 sw
rect 207 4081 208 4105
tri 210 4104 247 4141 ne
rect 247 4113 252 4141
tri 252 4113 278 4139 sw
rect 362 4123 371 4157
rect 362 4113 390 4123
rect 247 4104 331 4113
tri 247 4085 266 4104 ne
rect 266 4085 331 4104
rect 148 4059 208 4081
rect 330 4081 331 4085
rect 348 4081 390 4113
rect 330 4059 390 4081
rect 236 4043 253 4057
rect 285 4043 302 4057
tri 73 4007 95 4029 se
rect 95 4022 110 4043
tri 95 4007 110 4022 nw
rect 429 4022 444 4198
tri 444 4191 457 4204 nw
rect 530 4123 545 4361
tri 67 4001 73 4007 se
rect 73 4001 82 4007
rect 67 3985 82 4001
tri 82 3994 95 4007 nw
rect 236 3999 253 4013
rect 285 3999 302 4013
tri 429 4007 444 4022 ne
tri 444 4007 466 4029 sw
rect 67 3949 82 3957
rect 148 3985 208 3999
rect 163 3975 208 3985
rect 163 3957 191 3975
tri 67 3934 82 3949 ne
tri 82 3934 104 3956 sw
rect 148 3947 191 3957
rect 206 3971 208 3975
rect 330 3985 390 3999
tri 444 3994 457 4007 ne
rect 457 4001 466 4007
tri 466 4001 472 4007 sw
rect 330 3975 375 3985
rect 206 3947 280 3971
rect 148 3943 280 3947
tri 280 3943 308 3971 sw
rect 330 3961 332 3975
tri 330 3959 332 3961 ne
rect 344 3957 375 3975
rect 344 3947 390 3957
rect 457 3986 472 4001
tri 82 3922 94 3934 ne
rect 94 3929 104 3934
tri 104 3929 109 3934 sw
rect -7 3583 8 3811
rect 94 3821 109 3929
rect 148 3887 176 3943
tri 268 3925 286 3943 ne
rect 286 3923 308 3943
tri 308 3923 328 3943 sw
tri 344 3929 362 3947 ne
rect 167 3853 176 3887
rect 210 3914 252 3915
rect 210 3880 215 3914
rect 245 3880 252 3914
rect 210 3871 252 3880
rect 286 3914 328 3923
rect 286 3880 293 3914
rect 323 3880 328 3914
rect 286 3875 328 3880
rect 362 3887 390 3947
tri 435 3934 457 3956 se
rect 457 3949 472 3957
tri 457 3934 472 3949 nw
tri 429 3928 435 3934 se
rect 435 3928 444 3934
rect 148 3843 176 3853
tri 176 3843 200 3867 sw
rect 94 3773 110 3821
rect 148 3811 190 3843
tri 207 3835 208 3836 sw
rect 207 3811 208 3835
tri 210 3834 247 3871 ne
rect 247 3843 252 3871
tri 252 3843 278 3869 sw
rect 362 3853 371 3887
rect 362 3843 390 3853
rect 247 3834 331 3843
tri 247 3815 266 3834 ne
rect 266 3815 331 3834
rect 148 3789 208 3811
rect 330 3811 331 3815
rect 348 3811 390 3843
rect 330 3789 390 3811
rect 236 3773 253 3787
rect 285 3773 302 3787
tri 73 3737 95 3759 se
rect 95 3752 110 3773
tri 95 3737 110 3752 nw
rect 429 3752 444 3928
tri 444 3921 457 3934 nw
rect 530 3853 545 4081
tri 67 3731 73 3737 se
rect 73 3731 82 3737
rect 67 3715 82 3731
tri 82 3724 95 3737 nw
rect 236 3729 253 3743
rect 285 3729 302 3743
tri 429 3737 444 3752 ne
tri 444 3737 466 3759 sw
rect 67 3679 82 3687
rect 148 3715 208 3729
rect 163 3705 208 3715
rect 163 3687 191 3705
tri 67 3664 82 3679 ne
tri 82 3664 104 3686 sw
rect 148 3677 191 3687
rect 206 3701 208 3705
rect 330 3715 390 3729
tri 444 3724 457 3737 ne
rect 457 3731 466 3737
tri 466 3731 472 3737 sw
rect 330 3705 375 3715
rect 206 3677 280 3701
rect 148 3673 280 3677
tri 280 3673 308 3701 sw
rect 330 3691 332 3705
tri 330 3689 332 3691 ne
rect 344 3687 375 3705
rect 344 3677 390 3687
rect 457 3716 472 3731
tri 82 3652 94 3664 ne
rect 94 3659 104 3664
tri 104 3659 109 3664 sw
rect -7 3313 8 3541
rect 94 3503 109 3659
rect 148 3617 176 3673
tri 268 3655 286 3673 ne
rect 286 3653 308 3673
tri 308 3653 328 3673 sw
tri 344 3659 362 3677 ne
rect 167 3583 176 3617
rect 210 3644 252 3645
rect 210 3610 215 3644
rect 245 3610 252 3644
rect 210 3601 252 3610
rect 286 3644 328 3653
rect 286 3610 293 3644
rect 323 3610 328 3644
rect 286 3605 328 3610
rect 362 3617 390 3677
tri 435 3664 457 3686 se
rect 457 3679 472 3687
tri 457 3664 472 3679 nw
tri 429 3658 435 3664 se
rect 435 3658 444 3664
rect 148 3573 176 3583
tri 176 3573 200 3597 sw
rect 148 3541 190 3573
tri 207 3565 208 3566 sw
rect 207 3541 208 3565
tri 210 3564 247 3601 ne
rect 247 3573 252 3601
tri 252 3573 278 3599 sw
rect 362 3583 371 3617
rect 362 3573 390 3583
rect 247 3564 331 3573
tri 247 3545 266 3564 ne
rect 266 3545 331 3564
rect 148 3519 208 3541
rect 330 3541 331 3545
rect 348 3541 390 3573
rect 330 3519 390 3541
rect 236 3503 253 3517
rect 285 3503 302 3517
tri 73 3467 95 3489 se
rect 95 3482 110 3503
tri 95 3467 110 3482 nw
rect 429 3482 444 3658
tri 444 3651 457 3664 nw
rect 530 3583 545 3811
tri 67 3461 73 3467 se
rect 73 3461 82 3467
rect 67 3445 82 3461
tri 82 3454 95 3467 nw
rect 236 3459 253 3473
rect 285 3459 302 3473
tri 429 3467 444 3482 ne
tri 444 3467 466 3489 sw
rect 67 3409 82 3417
rect 148 3445 208 3459
rect 163 3435 208 3445
rect 163 3417 191 3435
tri 67 3394 82 3409 ne
tri 82 3394 104 3416 sw
rect 148 3407 191 3417
rect 206 3431 208 3435
rect 330 3445 390 3459
tri 444 3454 457 3467 ne
rect 457 3461 466 3467
tri 466 3461 472 3467 sw
rect 330 3435 375 3445
rect 206 3407 280 3431
rect 148 3403 280 3407
tri 280 3403 308 3431 sw
rect 330 3421 332 3435
tri 330 3419 332 3421 ne
rect 344 3417 375 3435
rect 344 3407 390 3417
rect 457 3446 472 3461
tri 82 3382 94 3394 ne
rect 94 3389 104 3394
tri 104 3389 109 3394 sw
rect -7 3043 8 3271
rect 94 3281 109 3389
rect 148 3347 176 3403
tri 268 3385 286 3403 ne
rect 286 3383 308 3403
tri 308 3383 328 3403 sw
tri 344 3389 362 3407 ne
rect 167 3313 176 3347
rect 210 3374 252 3375
rect 210 3340 215 3374
rect 245 3340 252 3374
rect 210 3331 252 3340
rect 286 3374 328 3383
rect 286 3340 293 3374
rect 323 3340 328 3374
rect 286 3335 328 3340
rect 362 3347 390 3407
tri 435 3394 457 3416 se
rect 457 3409 472 3417
tri 457 3394 472 3409 nw
tri 429 3388 435 3394 se
rect 435 3388 444 3394
rect 148 3303 176 3313
tri 176 3303 200 3327 sw
rect 94 3233 110 3281
rect 148 3271 190 3303
tri 207 3295 208 3296 sw
rect 207 3271 208 3295
tri 210 3294 247 3331 ne
rect 247 3303 252 3331
tri 252 3303 278 3329 sw
rect 362 3313 371 3347
rect 362 3303 390 3313
rect 247 3294 331 3303
tri 247 3275 266 3294 ne
rect 266 3275 331 3294
rect 148 3249 208 3271
rect 330 3271 331 3275
rect 348 3271 390 3303
rect 330 3249 390 3271
rect 236 3233 253 3247
rect 285 3233 302 3247
tri 73 3197 95 3219 se
rect 95 3212 110 3233
tri 95 3197 110 3212 nw
rect 429 3212 444 3388
tri 444 3381 457 3394 nw
rect 530 3313 545 3541
tri 67 3191 73 3197 se
rect 73 3191 82 3197
rect 67 3175 82 3191
tri 82 3184 95 3197 nw
rect 236 3189 253 3203
rect 285 3189 302 3203
tri 429 3197 444 3212 ne
tri 444 3197 466 3219 sw
rect 67 3139 82 3147
rect 148 3175 208 3189
rect 163 3165 208 3175
rect 163 3147 191 3165
tri 67 3124 82 3139 ne
tri 82 3124 104 3146 sw
rect 148 3137 191 3147
rect 206 3161 208 3165
rect 330 3175 390 3189
tri 444 3184 457 3197 ne
rect 457 3191 466 3197
tri 466 3191 472 3197 sw
rect 330 3165 375 3175
rect 206 3137 280 3161
rect 148 3133 280 3137
tri 280 3133 308 3161 sw
rect 330 3151 332 3165
tri 330 3149 332 3151 ne
rect 344 3147 375 3165
rect 344 3137 390 3147
rect 457 3176 472 3191
tri 82 3112 94 3124 ne
rect 94 3119 104 3124
tri 104 3119 109 3124 sw
rect -7 2773 8 3001
rect 94 2963 109 3119
rect 148 3077 176 3133
tri 268 3115 286 3133 ne
rect 286 3113 308 3133
tri 308 3113 328 3133 sw
tri 344 3119 362 3137 ne
rect 167 3043 176 3077
rect 210 3104 252 3105
rect 210 3070 215 3104
rect 245 3070 252 3104
rect 210 3061 252 3070
rect 286 3104 328 3113
rect 286 3070 293 3104
rect 323 3070 328 3104
rect 286 3065 328 3070
rect 362 3077 390 3137
tri 435 3124 457 3146 se
rect 457 3139 472 3147
tri 457 3124 472 3139 nw
tri 429 3118 435 3124 se
rect 435 3118 444 3124
rect 148 3033 176 3043
tri 176 3033 200 3057 sw
rect 148 3001 190 3033
tri 207 3025 208 3026 sw
rect 207 3001 208 3025
tri 210 3024 247 3061 ne
rect 247 3033 252 3061
tri 252 3033 278 3059 sw
rect 362 3043 371 3077
rect 362 3033 390 3043
rect 247 3024 331 3033
tri 247 3005 266 3024 ne
rect 266 3005 331 3024
rect 148 2979 208 3001
rect 330 3001 331 3005
rect 348 3001 390 3033
rect 330 2979 390 3001
rect 236 2963 253 2977
rect 285 2963 302 2977
tri 73 2927 95 2949 se
rect 95 2942 110 2963
tri 95 2927 110 2942 nw
rect 429 2942 444 3118
tri 444 3111 457 3124 nw
rect 530 3043 545 3271
tri 67 2921 73 2927 se
rect 73 2921 82 2927
rect 67 2905 82 2921
tri 82 2914 95 2927 nw
rect 236 2919 253 2933
rect 285 2919 302 2933
tri 429 2927 444 2942 ne
tri 444 2927 466 2949 sw
rect 67 2869 82 2877
rect 148 2905 208 2919
rect 163 2895 208 2905
rect 163 2877 191 2895
tri 67 2854 82 2869 ne
tri 82 2854 104 2876 sw
rect 148 2867 191 2877
rect 206 2891 208 2895
rect 330 2905 390 2919
tri 444 2914 457 2927 ne
rect 457 2921 466 2927
tri 466 2921 472 2927 sw
rect 330 2895 375 2905
rect 206 2867 280 2891
rect 148 2863 280 2867
tri 280 2863 308 2891 sw
rect 330 2881 332 2895
tri 330 2879 332 2881 ne
rect 344 2877 375 2895
rect 344 2867 390 2877
rect 457 2906 472 2921
tri 82 2842 94 2854 ne
rect 94 2849 104 2854
tri 104 2849 109 2854 sw
rect -7 2503 8 2731
rect 94 2741 109 2849
rect 148 2807 176 2863
tri 268 2845 286 2863 ne
rect 286 2843 308 2863
tri 308 2843 328 2863 sw
tri 344 2849 362 2867 ne
rect 167 2773 176 2807
rect 210 2834 252 2835
rect 210 2800 215 2834
rect 245 2800 252 2834
rect 210 2791 252 2800
rect 286 2834 328 2843
rect 286 2800 293 2834
rect 323 2800 328 2834
rect 286 2795 328 2800
rect 362 2807 390 2867
tri 435 2854 457 2876 se
rect 457 2869 472 2877
tri 457 2854 472 2869 nw
tri 429 2848 435 2854 se
rect 435 2848 444 2854
rect 148 2763 176 2773
tri 176 2763 200 2787 sw
rect 94 2693 110 2741
rect 148 2731 190 2763
tri 207 2755 208 2756 sw
rect 207 2731 208 2755
tri 210 2754 247 2791 ne
rect 247 2763 252 2791
tri 252 2763 278 2789 sw
rect 362 2773 371 2807
rect 362 2763 390 2773
rect 247 2754 331 2763
tri 247 2735 266 2754 ne
rect 266 2735 331 2754
rect 148 2709 208 2731
rect 330 2731 331 2735
rect 348 2731 390 2763
rect 330 2709 390 2731
rect 236 2693 253 2707
rect 285 2693 302 2707
tri 73 2657 95 2679 se
rect 95 2672 110 2693
tri 95 2657 110 2672 nw
rect 429 2672 444 2848
tri 444 2841 457 2854 nw
rect 530 2773 545 3001
tri 67 2651 73 2657 se
rect 73 2651 82 2657
rect 67 2635 82 2651
tri 82 2644 95 2657 nw
rect 236 2649 253 2663
rect 285 2649 302 2663
tri 429 2657 444 2672 ne
tri 444 2657 466 2679 sw
rect 67 2599 82 2607
rect 148 2635 208 2649
rect 163 2625 208 2635
rect 163 2607 191 2625
tri 67 2584 82 2599 ne
tri 82 2584 104 2606 sw
rect 148 2597 191 2607
rect 206 2621 208 2625
rect 330 2635 390 2649
tri 444 2644 457 2657 ne
rect 457 2651 466 2657
tri 466 2651 472 2657 sw
rect 330 2625 375 2635
rect 206 2597 280 2621
rect 148 2593 280 2597
tri 280 2593 308 2621 sw
rect 330 2611 332 2625
tri 330 2609 332 2611 ne
rect 344 2607 375 2625
rect 344 2597 390 2607
rect 457 2636 472 2651
tri 82 2572 94 2584 ne
rect 94 2579 104 2584
tri 104 2579 109 2584 sw
rect -7 2233 8 2461
rect 94 2423 109 2579
rect 148 2537 176 2593
tri 268 2575 286 2593 ne
rect 286 2573 308 2593
tri 308 2573 328 2593 sw
tri 344 2579 362 2597 ne
rect 167 2503 176 2537
rect 210 2564 252 2565
rect 210 2530 215 2564
rect 245 2530 252 2564
rect 210 2521 252 2530
rect 286 2564 328 2573
rect 286 2530 293 2564
rect 323 2530 328 2564
rect 286 2525 328 2530
rect 362 2537 390 2597
tri 435 2584 457 2606 se
rect 457 2599 472 2607
tri 457 2584 472 2599 nw
tri 429 2578 435 2584 se
rect 435 2578 444 2584
rect 148 2493 176 2503
tri 176 2493 200 2517 sw
rect 148 2461 190 2493
tri 207 2485 208 2486 sw
rect 207 2461 208 2485
tri 210 2484 247 2521 ne
rect 247 2493 252 2521
tri 252 2493 278 2519 sw
rect 362 2503 371 2537
rect 362 2493 390 2503
rect 247 2484 331 2493
tri 247 2465 266 2484 ne
rect 266 2465 331 2484
rect 148 2439 208 2461
rect 330 2461 331 2465
rect 348 2461 390 2493
rect 330 2439 390 2461
rect 236 2423 253 2437
rect 285 2423 302 2437
tri 73 2387 95 2409 se
rect 95 2402 110 2423
tri 95 2387 110 2402 nw
rect 429 2402 444 2578
tri 444 2571 457 2584 nw
rect 530 2503 545 2731
tri 67 2381 73 2387 se
rect 73 2381 82 2387
rect 67 2365 82 2381
tri 82 2374 95 2387 nw
rect 236 2379 253 2393
rect 285 2379 302 2393
tri 429 2387 444 2402 ne
tri 444 2387 466 2409 sw
rect 67 2329 82 2337
rect 148 2365 208 2379
rect 163 2355 208 2365
rect 163 2337 191 2355
tri 67 2314 82 2329 ne
tri 82 2314 104 2336 sw
rect 148 2327 191 2337
rect 206 2351 208 2355
rect 330 2365 390 2379
tri 444 2374 457 2387 ne
rect 457 2381 466 2387
tri 466 2381 472 2387 sw
rect 330 2355 375 2365
rect 206 2327 280 2351
rect 148 2323 280 2327
tri 280 2323 308 2351 sw
rect 330 2341 332 2355
tri 330 2339 332 2341 ne
rect 344 2337 375 2355
rect 344 2327 390 2337
rect 457 2366 472 2381
tri 82 2302 94 2314 ne
rect 94 2309 104 2314
tri 104 2309 109 2314 sw
rect -7 1963 8 2191
rect 94 2201 109 2309
rect 148 2267 176 2323
tri 268 2305 286 2323 ne
rect 286 2303 308 2323
tri 308 2303 328 2323 sw
tri 344 2309 362 2327 ne
rect 167 2233 176 2267
rect 210 2294 252 2295
rect 210 2260 215 2294
rect 245 2260 252 2294
rect 210 2251 252 2260
rect 286 2294 328 2303
rect 286 2260 293 2294
rect 323 2260 328 2294
rect 286 2255 328 2260
rect 362 2267 390 2327
tri 435 2314 457 2336 se
rect 457 2329 472 2337
tri 457 2314 472 2329 nw
tri 429 2308 435 2314 se
rect 435 2308 444 2314
rect 148 2223 176 2233
tri 176 2223 200 2247 sw
rect 94 2153 110 2201
rect 148 2191 190 2223
tri 207 2215 208 2216 sw
rect 207 2191 208 2215
tri 210 2214 247 2251 ne
rect 247 2223 252 2251
tri 252 2223 278 2249 sw
rect 362 2233 371 2267
rect 362 2223 390 2233
rect 247 2214 331 2223
tri 247 2195 266 2214 ne
rect 266 2195 331 2214
rect 148 2169 208 2191
rect 330 2191 331 2195
rect 348 2191 390 2223
rect 330 2169 390 2191
rect 236 2153 253 2167
rect 285 2153 302 2167
tri 73 2117 95 2139 se
rect 95 2132 110 2153
tri 95 2117 110 2132 nw
rect 429 2132 444 2308
tri 444 2301 457 2314 nw
rect 530 2233 545 2461
tri 67 2111 73 2117 se
rect 73 2111 82 2117
rect 67 2095 82 2111
tri 82 2104 95 2117 nw
rect 236 2109 253 2123
rect 285 2109 302 2123
tri 429 2117 444 2132 ne
tri 444 2117 466 2139 sw
rect 67 2059 82 2067
rect 148 2095 208 2109
rect 163 2085 208 2095
rect 163 2067 191 2085
tri 67 2044 82 2059 ne
tri 82 2044 104 2066 sw
rect 148 2057 191 2067
rect 206 2081 208 2085
rect 330 2095 390 2109
tri 444 2104 457 2117 ne
rect 457 2111 466 2117
tri 466 2111 472 2117 sw
rect 330 2085 375 2095
rect 206 2057 280 2081
rect 148 2053 280 2057
tri 280 2053 308 2081 sw
rect 330 2071 332 2085
tri 330 2069 332 2071 ne
rect 344 2067 375 2085
rect 344 2057 390 2067
rect 457 2096 472 2111
tri 82 2032 94 2044 ne
rect 94 2039 104 2044
tri 104 2039 109 2044 sw
rect -7 1693 8 1921
rect 94 1883 109 2039
rect 148 1997 176 2053
tri 268 2035 286 2053 ne
rect 286 2033 308 2053
tri 308 2033 328 2053 sw
tri 344 2039 362 2057 ne
rect 167 1963 176 1997
rect 210 2024 252 2025
rect 210 1990 215 2024
rect 245 1990 252 2024
rect 210 1981 252 1990
rect 286 2024 328 2033
rect 286 1990 293 2024
rect 323 1990 328 2024
rect 286 1985 328 1990
rect 362 1997 390 2057
tri 435 2044 457 2066 se
rect 457 2059 472 2067
tri 457 2044 472 2059 nw
tri 429 2038 435 2044 se
rect 435 2038 444 2044
rect 148 1953 176 1963
tri 176 1953 200 1977 sw
rect 148 1921 190 1953
tri 207 1945 208 1946 sw
rect 207 1921 208 1945
tri 210 1944 247 1981 ne
rect 247 1953 252 1981
tri 252 1953 278 1979 sw
rect 362 1963 371 1997
rect 362 1953 390 1963
rect 247 1944 331 1953
tri 247 1925 266 1944 ne
rect 266 1925 331 1944
rect 148 1899 208 1921
rect 330 1921 331 1925
rect 348 1921 390 1953
rect 330 1899 390 1921
rect 236 1883 253 1897
rect 285 1883 302 1897
tri 73 1847 95 1869 se
rect 95 1862 110 1883
tri 95 1847 110 1862 nw
rect 429 1862 444 2038
tri 444 2031 457 2044 nw
rect 530 1963 545 2191
tri 67 1841 73 1847 se
rect 73 1841 82 1847
rect 67 1825 82 1841
tri 82 1834 95 1847 nw
rect 236 1839 253 1853
rect 285 1839 302 1853
tri 429 1847 444 1862 ne
tri 444 1847 466 1869 sw
rect 67 1789 82 1797
rect 148 1825 208 1839
rect 163 1815 208 1825
rect 163 1797 191 1815
tri 67 1774 82 1789 ne
tri 82 1774 104 1796 sw
rect 148 1787 191 1797
rect 206 1811 208 1815
rect 330 1825 390 1839
tri 444 1834 457 1847 ne
rect 457 1841 466 1847
tri 466 1841 472 1847 sw
rect 330 1815 375 1825
rect 206 1787 280 1811
rect 148 1783 280 1787
tri 280 1783 308 1811 sw
rect 330 1801 332 1815
tri 330 1799 332 1801 ne
rect 344 1797 375 1815
rect 344 1787 390 1797
rect 457 1826 472 1841
tri 82 1762 94 1774 ne
rect 94 1769 104 1774
tri 104 1769 109 1774 sw
rect -7 1423 8 1651
rect 94 1661 109 1769
rect 148 1727 176 1783
tri 268 1765 286 1783 ne
rect 286 1763 308 1783
tri 308 1763 328 1783 sw
tri 344 1769 362 1787 ne
rect 167 1693 176 1727
rect 210 1754 252 1755
rect 210 1720 215 1754
rect 245 1720 252 1754
rect 210 1711 252 1720
rect 286 1754 328 1763
rect 286 1720 293 1754
rect 323 1720 328 1754
rect 286 1715 328 1720
rect 362 1727 390 1787
tri 435 1774 457 1796 se
rect 457 1789 472 1797
tri 457 1774 472 1789 nw
tri 429 1768 435 1774 se
rect 435 1768 444 1774
rect 148 1683 176 1693
tri 176 1683 200 1707 sw
rect 94 1613 110 1661
rect 148 1651 190 1683
tri 207 1675 208 1676 sw
rect 207 1651 208 1675
tri 210 1674 247 1711 ne
rect 247 1683 252 1711
tri 252 1683 278 1709 sw
rect 362 1693 371 1727
rect 362 1683 390 1693
rect 247 1674 331 1683
tri 247 1655 266 1674 ne
rect 266 1655 331 1674
rect 148 1629 208 1651
rect 330 1651 331 1655
rect 348 1651 390 1683
rect 330 1629 390 1651
rect 236 1613 253 1627
rect 285 1613 302 1627
tri 73 1577 95 1599 se
rect 95 1592 110 1613
tri 95 1577 110 1592 nw
rect 429 1592 444 1768
tri 444 1761 457 1774 nw
rect 530 1693 545 1921
tri 67 1571 73 1577 se
rect 73 1571 82 1577
rect 67 1555 82 1571
tri 82 1564 95 1577 nw
rect 236 1569 253 1583
rect 285 1569 302 1583
tri 429 1577 444 1592 ne
tri 444 1577 466 1599 sw
rect 67 1519 82 1527
rect 148 1555 208 1569
rect 163 1545 208 1555
rect 163 1527 191 1545
tri 67 1504 82 1519 ne
tri 82 1504 104 1526 sw
rect 148 1517 191 1527
rect 206 1541 208 1545
rect 330 1555 390 1569
tri 444 1564 457 1577 ne
rect 457 1571 466 1577
tri 466 1571 472 1577 sw
rect 330 1545 375 1555
rect 206 1517 280 1541
rect 148 1513 280 1517
tri 280 1513 308 1541 sw
rect 330 1531 332 1545
tri 330 1529 332 1531 ne
rect 344 1527 375 1545
rect 344 1517 390 1527
rect 457 1556 472 1571
tri 82 1492 94 1504 ne
rect 94 1499 104 1504
tri 104 1499 109 1504 sw
rect -7 1153 8 1381
rect 94 1343 109 1499
rect 148 1457 176 1513
tri 268 1495 286 1513 ne
rect 286 1493 308 1513
tri 308 1493 328 1513 sw
tri 344 1499 362 1517 ne
rect 167 1423 176 1457
rect 210 1484 252 1485
rect 210 1450 215 1484
rect 245 1450 252 1484
rect 210 1441 252 1450
rect 286 1484 328 1493
rect 286 1450 293 1484
rect 323 1450 328 1484
rect 286 1445 328 1450
rect 362 1457 390 1517
tri 435 1504 457 1526 se
rect 457 1519 472 1527
tri 457 1504 472 1519 nw
tri 429 1498 435 1504 se
rect 435 1498 444 1504
rect 148 1413 176 1423
tri 176 1413 200 1437 sw
rect 148 1381 190 1413
tri 207 1405 208 1406 sw
rect 207 1381 208 1405
tri 210 1404 247 1441 ne
rect 247 1413 252 1441
tri 252 1413 278 1439 sw
rect 362 1423 371 1457
rect 362 1413 390 1423
rect 247 1404 331 1413
tri 247 1385 266 1404 ne
rect 266 1385 331 1404
rect 148 1359 208 1381
rect 330 1381 331 1385
rect 348 1381 390 1413
rect 330 1359 390 1381
rect 236 1343 253 1357
rect 285 1343 302 1357
tri 73 1307 95 1329 se
rect 95 1322 110 1343
tri 95 1307 110 1322 nw
rect 429 1322 444 1498
tri 444 1491 457 1504 nw
rect 530 1423 545 1651
tri 67 1301 73 1307 se
rect 73 1301 82 1307
rect 67 1285 82 1301
tri 82 1294 95 1307 nw
rect 236 1299 253 1313
rect 285 1299 302 1313
tri 429 1307 444 1322 ne
tri 444 1307 466 1329 sw
rect 67 1249 82 1257
rect 148 1285 208 1299
rect 163 1275 208 1285
rect 163 1257 191 1275
tri 67 1234 82 1249 ne
tri 82 1234 104 1256 sw
rect 148 1247 191 1257
rect 206 1271 208 1275
rect 330 1285 390 1299
tri 444 1294 457 1307 ne
rect 457 1301 466 1307
tri 466 1301 472 1307 sw
rect 330 1275 375 1285
rect 206 1247 280 1271
rect 148 1243 280 1247
tri 280 1243 308 1271 sw
rect 330 1261 332 1275
tri 330 1259 332 1261 ne
rect 344 1257 375 1275
rect 344 1247 390 1257
rect 457 1286 472 1301
tri 82 1222 94 1234 ne
rect 94 1229 104 1234
tri 104 1229 109 1234 sw
rect -7 883 8 1111
rect 94 1121 109 1229
rect 148 1187 176 1243
tri 268 1225 286 1243 ne
rect 286 1223 308 1243
tri 308 1223 328 1243 sw
tri 344 1229 362 1247 ne
rect 167 1153 176 1187
rect 210 1214 252 1215
rect 210 1180 215 1214
rect 245 1180 252 1214
rect 210 1171 252 1180
rect 286 1214 328 1223
rect 286 1180 293 1214
rect 323 1180 328 1214
rect 286 1175 328 1180
rect 362 1187 390 1247
tri 435 1234 457 1256 se
rect 457 1249 472 1257
tri 457 1234 472 1249 nw
tri 429 1228 435 1234 se
rect 435 1228 444 1234
rect 148 1143 176 1153
tri 176 1143 200 1167 sw
rect 94 1073 110 1121
rect 148 1111 190 1143
tri 207 1135 208 1136 sw
rect 207 1111 208 1135
tri 210 1134 247 1171 ne
rect 247 1143 252 1171
tri 252 1143 278 1169 sw
rect 362 1153 371 1187
rect 362 1143 390 1153
rect 247 1134 331 1143
tri 247 1115 266 1134 ne
rect 266 1115 331 1134
rect 148 1089 208 1111
rect 330 1111 331 1115
rect 348 1111 390 1143
rect 330 1089 390 1111
rect 236 1073 253 1087
rect 285 1073 302 1087
tri 73 1037 95 1059 se
rect 95 1052 110 1073
tri 95 1037 110 1052 nw
rect 429 1052 444 1228
tri 444 1221 457 1234 nw
rect 530 1153 545 1381
tri 67 1031 73 1037 se
rect 73 1031 82 1037
rect 67 1015 82 1031
tri 82 1024 95 1037 nw
rect 236 1029 253 1043
rect 285 1029 302 1043
tri 429 1037 444 1052 ne
tri 444 1037 466 1059 sw
rect 67 979 82 987
rect 148 1015 208 1029
rect 163 1005 208 1015
rect 163 987 191 1005
tri 67 964 82 979 ne
tri 82 964 104 986 sw
rect 148 977 191 987
rect 206 1001 208 1005
rect 330 1015 390 1029
tri 444 1024 457 1037 ne
rect 457 1031 466 1037
tri 466 1031 472 1037 sw
rect 330 1005 375 1015
rect 206 977 280 1001
rect 148 973 280 977
tri 280 973 308 1001 sw
rect 330 991 332 1005
tri 330 989 332 991 ne
rect 344 987 375 1005
rect 344 977 390 987
rect 457 1016 472 1031
tri 82 952 94 964 ne
rect 94 959 104 964
tri 104 959 109 964 sw
rect -7 613 8 841
rect 94 803 109 959
rect 148 917 176 973
tri 268 955 286 973 ne
rect 286 953 308 973
tri 308 953 328 973 sw
tri 344 959 362 977 ne
rect 167 883 176 917
rect 210 944 252 945
rect 210 910 215 944
rect 245 910 252 944
rect 210 901 252 910
rect 286 944 328 953
rect 286 910 293 944
rect 323 910 328 944
rect 286 905 328 910
rect 362 917 390 977
tri 435 964 457 986 se
rect 457 979 472 987
tri 457 964 472 979 nw
tri 429 958 435 964 se
rect 435 958 444 964
rect 148 873 176 883
tri 176 873 200 897 sw
rect 148 841 190 873
tri 207 865 208 866 sw
rect 207 841 208 865
tri 210 864 247 901 ne
rect 247 873 252 901
tri 252 873 278 899 sw
rect 362 883 371 917
rect 362 873 390 883
rect 247 864 331 873
tri 247 845 266 864 ne
rect 266 845 331 864
rect 148 819 208 841
rect 330 841 331 845
rect 348 841 390 873
rect 330 819 390 841
rect 236 803 253 817
rect 285 803 302 817
tri 73 767 95 789 se
rect 95 782 110 803
tri 95 767 110 782 nw
rect 429 782 444 958
tri 444 951 457 964 nw
rect 530 883 545 1111
tri 67 761 73 767 se
rect 73 761 82 767
rect 67 745 82 761
tri 82 754 95 767 nw
rect 236 759 253 773
rect 285 759 302 773
tri 429 767 444 782 ne
tri 444 767 466 789 sw
rect 67 709 82 717
rect 148 745 208 759
rect 163 735 208 745
rect 163 717 191 735
tri 67 694 82 709 ne
tri 82 694 104 716 sw
rect 148 707 191 717
rect 206 731 208 735
rect 330 745 390 759
tri 444 754 457 767 ne
rect 457 761 466 767
tri 466 761 472 767 sw
rect 330 735 375 745
rect 206 707 280 731
rect 148 703 280 707
tri 280 703 308 731 sw
rect 330 721 332 735
tri 330 719 332 721 ne
rect 344 717 375 735
rect 344 707 390 717
rect 457 746 472 761
tri 82 682 94 694 ne
rect 94 689 104 694
tri 104 689 109 694 sw
rect -7 343 8 571
rect 94 581 109 689
rect 148 647 176 703
tri 268 685 286 703 ne
rect 286 683 308 703
tri 308 683 328 703 sw
tri 344 689 362 707 ne
rect 167 613 176 647
rect 210 674 252 675
rect 210 640 215 674
rect 245 640 252 674
rect 210 631 252 640
rect 286 674 328 683
rect 286 640 293 674
rect 323 640 328 674
rect 286 635 328 640
rect 362 647 390 707
tri 435 694 457 716 se
rect 457 709 472 717
tri 457 694 472 709 nw
tri 429 688 435 694 se
rect 435 688 444 694
rect 148 603 176 613
tri 176 603 200 627 sw
rect 94 533 110 581
rect 148 571 190 603
tri 207 595 208 596 sw
rect 207 571 208 595
tri 210 594 247 631 ne
rect 247 603 252 631
tri 252 603 278 629 sw
rect 362 613 371 647
rect 362 603 390 613
rect 247 594 331 603
tri 247 575 266 594 ne
rect 266 575 331 594
rect 148 549 208 571
rect 330 571 331 575
rect 348 571 390 603
rect 330 549 390 571
rect 236 533 253 547
rect 285 533 302 547
tri 73 497 95 519 se
rect 95 512 110 533
tri 95 497 110 512 nw
rect 429 512 444 688
tri 444 681 457 694 nw
rect 530 613 545 841
tri 67 491 73 497 se
rect 73 491 82 497
rect 67 475 82 491
tri 82 484 95 497 nw
rect 236 489 253 503
rect 285 489 302 503
tri 429 497 444 512 ne
tri 444 497 466 519 sw
rect 67 439 82 447
rect 148 475 208 489
rect 163 465 208 475
rect 163 447 191 465
tri 67 424 82 439 ne
tri 82 424 104 446 sw
rect 148 437 191 447
rect 206 461 208 465
rect 330 475 390 489
tri 444 484 457 497 ne
rect 457 491 466 497
tri 466 491 472 497 sw
rect 330 465 375 475
rect 206 437 280 461
rect 148 433 280 437
tri 280 433 308 461 sw
rect 330 451 332 465
tri 330 449 332 451 ne
rect 344 447 375 465
rect 344 437 390 447
rect 457 476 472 491
tri 82 412 94 424 ne
rect 94 419 104 424
tri 104 419 109 424 sw
rect -7 73 8 301
rect 94 263 109 419
rect 148 377 176 433
tri 268 415 286 433 ne
rect 286 413 308 433
tri 308 413 328 433 sw
tri 344 419 362 437 ne
rect 167 343 176 377
rect 210 404 252 405
rect 210 370 215 404
rect 245 370 252 404
rect 210 361 252 370
rect 286 404 328 413
rect 286 370 293 404
rect 323 370 328 404
rect 286 365 328 370
rect 362 377 390 437
tri 435 424 457 446 se
rect 457 439 472 447
tri 457 424 472 439 nw
tri 429 418 435 424 se
rect 435 418 444 424
rect 148 333 176 343
tri 176 333 200 357 sw
rect 148 301 190 333
tri 207 325 208 326 sw
rect 207 301 208 325
tri 210 324 247 361 ne
rect 247 333 252 361
tri 252 333 278 359 sw
rect 362 343 371 377
rect 362 333 390 343
rect 247 324 331 333
tri 247 305 266 324 ne
rect 266 305 331 324
rect 148 279 208 301
rect 330 301 331 305
rect 348 301 390 333
rect 330 279 390 301
rect 236 263 253 277
rect 285 263 302 277
tri 73 227 95 249 se
rect 95 242 110 263
tri 95 227 110 242 nw
rect 429 242 444 418
tri 444 411 457 424 nw
rect 530 343 545 571
tri 67 221 73 227 se
rect 73 221 82 227
rect 67 205 82 221
tri 82 214 95 227 nw
rect 236 219 253 233
rect 285 219 302 233
tri 429 227 444 242 ne
tri 444 227 466 249 sw
rect 67 169 82 177
rect 148 205 208 219
rect 163 195 208 205
rect 163 177 191 195
tri 67 154 82 169 ne
tri 82 154 104 176 sw
rect 148 167 191 177
rect 206 191 208 195
rect 330 205 390 219
tri 444 214 457 227 ne
rect 457 221 466 227
tri 466 221 472 227 sw
rect 330 195 375 205
rect 206 167 280 191
rect 148 163 280 167
tri 280 163 308 191 sw
rect 330 181 332 195
tri 330 179 332 181 ne
rect 344 177 375 195
rect 344 167 390 177
rect 457 206 472 221
tri 82 142 94 154 ne
rect 94 149 104 154
tri 104 149 109 154 sw
rect -7 -55 8 31
rect 94 -55 109 149
rect 148 107 176 163
tri 268 145 286 163 ne
rect 286 143 308 163
tri 308 143 328 163 sw
tri 344 149 362 167 ne
rect 167 73 176 107
rect 210 134 252 135
rect 210 100 215 134
rect 245 100 252 134
rect 210 91 252 100
rect 286 134 328 143
rect 286 100 293 134
rect 323 100 328 134
rect 286 95 328 100
rect 362 107 390 167
tri 435 154 457 176 se
rect 457 169 472 177
tri 457 154 472 169 nw
tri 429 148 435 154 se
rect 435 148 444 154
rect 148 63 176 73
tri 176 63 200 87 sw
rect 148 31 190 63
tri 207 55 208 56 sw
rect 207 31 208 55
tri 210 54 247 91 ne
rect 247 63 252 91
tri 252 63 278 89 sw
rect 362 73 371 107
rect 362 63 390 73
rect 247 54 331 63
tri 247 35 266 54 ne
rect 266 35 331 54
rect 148 9 208 31
rect 330 31 331 35
rect 348 31 390 63
rect 330 9 390 31
rect 236 -7 253 7
rect 285 -7 302 7
rect 429 -55 444 148
tri 444 141 457 154 nw
rect 530 73 545 301
rect 530 -55 545 31
rect 573 4123 588 4361
tri 653 4277 675 4299 se
rect 675 4292 690 4361
tri 675 4277 690 4292 nw
rect 1009 4292 1024 4361
tri 647 4271 653 4277 se
rect 653 4271 662 4277
rect 647 4255 662 4271
tri 662 4264 675 4277 nw
rect 816 4269 833 4283
rect 865 4269 882 4283
tri 1009 4277 1024 4292 ne
tri 1024 4277 1046 4299 sw
rect 647 4219 662 4227
rect 728 4255 788 4269
rect 743 4245 788 4255
rect 743 4227 771 4245
tri 647 4204 662 4219 ne
tri 662 4204 684 4226 sw
rect 728 4217 771 4227
rect 786 4241 788 4245
rect 910 4255 970 4269
tri 1024 4264 1037 4277 ne
rect 1037 4271 1046 4277
tri 1046 4271 1052 4277 sw
rect 910 4245 955 4255
rect 786 4217 860 4241
rect 728 4213 860 4217
tri 860 4213 888 4241 sw
rect 910 4231 912 4245
tri 910 4229 912 4231 ne
rect 924 4227 955 4245
rect 924 4217 970 4227
rect 1037 4256 1052 4271
tri 662 4192 674 4204 ne
rect 674 4199 684 4204
tri 684 4199 689 4204 sw
rect 573 3853 588 4081
rect 674 4043 689 4199
rect 728 4157 756 4213
tri 848 4195 866 4213 ne
rect 866 4193 888 4213
tri 888 4193 908 4213 sw
tri 924 4199 942 4217 ne
rect 747 4123 756 4157
rect 790 4184 832 4185
rect 790 4150 795 4184
rect 825 4150 832 4184
rect 790 4141 832 4150
rect 866 4184 908 4193
rect 866 4150 873 4184
rect 903 4150 908 4184
rect 866 4145 908 4150
rect 942 4157 970 4217
tri 1015 4204 1037 4226 se
rect 1037 4219 1052 4227
tri 1037 4204 1052 4219 nw
tri 1009 4198 1015 4204 se
rect 1015 4198 1024 4204
rect 728 4113 756 4123
tri 756 4113 780 4137 sw
rect 728 4081 770 4113
tri 787 4105 788 4106 sw
rect 787 4081 788 4105
tri 790 4104 827 4141 ne
rect 827 4113 832 4141
tri 832 4113 858 4139 sw
rect 942 4123 951 4157
rect 942 4113 970 4123
rect 827 4104 911 4113
tri 827 4085 846 4104 ne
rect 846 4085 911 4104
rect 728 4059 788 4081
rect 910 4081 911 4085
rect 928 4081 970 4113
rect 910 4059 970 4081
rect 816 4043 833 4057
rect 865 4043 882 4057
tri 653 4007 675 4029 se
rect 675 4022 690 4043
tri 675 4007 690 4022 nw
rect 1009 4022 1024 4198
tri 1024 4191 1037 4204 nw
rect 1110 4123 1125 4361
tri 647 4001 653 4007 se
rect 653 4001 662 4007
rect 647 3985 662 4001
tri 662 3994 675 4007 nw
rect 816 3999 833 4013
rect 865 3999 882 4013
tri 1009 4007 1024 4022 ne
tri 1024 4007 1046 4029 sw
rect 647 3949 662 3957
rect 728 3985 788 3999
rect 743 3975 788 3985
rect 743 3957 771 3975
tri 647 3934 662 3949 ne
tri 662 3934 684 3956 sw
rect 728 3947 771 3957
rect 786 3971 788 3975
rect 910 3985 970 3999
tri 1024 3994 1037 4007 ne
rect 1037 4001 1046 4007
tri 1046 4001 1052 4007 sw
rect 910 3975 955 3985
rect 786 3947 860 3971
rect 728 3943 860 3947
tri 860 3943 888 3971 sw
rect 910 3961 912 3975
tri 910 3959 912 3961 ne
rect 924 3957 955 3975
rect 924 3947 970 3957
rect 1037 3986 1052 4001
tri 662 3922 674 3934 ne
rect 674 3929 684 3934
tri 684 3929 689 3934 sw
rect 573 3583 588 3811
rect 674 3821 689 3929
rect 728 3887 756 3943
tri 848 3925 866 3943 ne
rect 866 3923 888 3943
tri 888 3923 908 3943 sw
tri 924 3929 942 3947 ne
rect 747 3853 756 3887
rect 790 3914 832 3915
rect 790 3880 795 3914
rect 825 3880 832 3914
rect 790 3871 832 3880
rect 866 3914 908 3923
rect 866 3880 873 3914
rect 903 3880 908 3914
rect 866 3875 908 3880
rect 942 3887 970 3947
tri 1015 3934 1037 3956 se
rect 1037 3949 1052 3957
tri 1037 3934 1052 3949 nw
tri 1009 3928 1015 3934 se
rect 1015 3928 1024 3934
rect 728 3843 756 3853
tri 756 3843 780 3867 sw
rect 674 3773 690 3821
rect 728 3811 770 3843
tri 787 3835 788 3836 sw
rect 787 3811 788 3835
tri 790 3834 827 3871 ne
rect 827 3843 832 3871
tri 832 3843 858 3869 sw
rect 942 3853 951 3887
rect 942 3843 970 3853
rect 827 3834 911 3843
tri 827 3815 846 3834 ne
rect 846 3815 911 3834
rect 728 3789 788 3811
rect 910 3811 911 3815
rect 928 3811 970 3843
rect 910 3789 970 3811
rect 816 3773 833 3787
rect 865 3773 882 3787
tri 653 3737 675 3759 se
rect 675 3752 690 3773
tri 675 3737 690 3752 nw
rect 1009 3752 1024 3928
tri 1024 3921 1037 3934 nw
rect 1110 3853 1125 4081
tri 647 3731 653 3737 se
rect 653 3731 662 3737
rect 647 3715 662 3731
tri 662 3724 675 3737 nw
rect 816 3729 833 3743
rect 865 3729 882 3743
tri 1009 3737 1024 3752 ne
tri 1024 3737 1046 3759 sw
rect 647 3679 662 3687
rect 728 3715 788 3729
rect 743 3705 788 3715
rect 743 3687 771 3705
tri 647 3664 662 3679 ne
tri 662 3664 684 3686 sw
rect 728 3677 771 3687
rect 786 3701 788 3705
rect 910 3715 970 3729
tri 1024 3724 1037 3737 ne
rect 1037 3731 1046 3737
tri 1046 3731 1052 3737 sw
rect 910 3705 955 3715
rect 786 3677 860 3701
rect 728 3673 860 3677
tri 860 3673 888 3701 sw
rect 910 3691 912 3705
tri 910 3689 912 3691 ne
rect 924 3687 955 3705
rect 924 3677 970 3687
rect 1037 3716 1052 3731
tri 662 3652 674 3664 ne
rect 674 3659 684 3664
tri 684 3659 689 3664 sw
rect 573 3313 588 3541
rect 674 3503 689 3659
rect 728 3617 756 3673
tri 848 3655 866 3673 ne
rect 866 3653 888 3673
tri 888 3653 908 3673 sw
tri 924 3659 942 3677 ne
rect 747 3583 756 3617
rect 790 3644 832 3645
rect 790 3610 795 3644
rect 825 3610 832 3644
rect 790 3601 832 3610
rect 866 3644 908 3653
rect 866 3610 873 3644
rect 903 3610 908 3644
rect 866 3605 908 3610
rect 942 3617 970 3677
tri 1015 3664 1037 3686 se
rect 1037 3679 1052 3687
tri 1037 3664 1052 3679 nw
tri 1009 3658 1015 3664 se
rect 1015 3658 1024 3664
rect 728 3573 756 3583
tri 756 3573 780 3597 sw
rect 728 3541 770 3573
tri 787 3565 788 3566 sw
rect 787 3541 788 3565
tri 790 3564 827 3601 ne
rect 827 3573 832 3601
tri 832 3573 858 3599 sw
rect 942 3583 951 3617
rect 942 3573 970 3583
rect 827 3564 911 3573
tri 827 3545 846 3564 ne
rect 846 3545 911 3564
rect 728 3519 788 3541
rect 910 3541 911 3545
rect 928 3541 970 3573
rect 910 3519 970 3541
rect 816 3503 833 3517
rect 865 3503 882 3517
tri 653 3467 675 3489 se
rect 675 3482 690 3503
tri 675 3467 690 3482 nw
rect 1009 3482 1024 3658
tri 1024 3651 1037 3664 nw
rect 1110 3583 1125 3811
tri 647 3461 653 3467 se
rect 653 3461 662 3467
rect 647 3445 662 3461
tri 662 3454 675 3467 nw
rect 816 3459 833 3473
rect 865 3459 882 3473
tri 1009 3467 1024 3482 ne
tri 1024 3467 1046 3489 sw
rect 647 3409 662 3417
rect 728 3445 788 3459
rect 743 3435 788 3445
rect 743 3417 771 3435
tri 647 3394 662 3409 ne
tri 662 3394 684 3416 sw
rect 728 3407 771 3417
rect 786 3431 788 3435
rect 910 3445 970 3459
tri 1024 3454 1037 3467 ne
rect 1037 3461 1046 3467
tri 1046 3461 1052 3467 sw
rect 910 3435 955 3445
rect 786 3407 860 3431
rect 728 3403 860 3407
tri 860 3403 888 3431 sw
rect 910 3421 912 3435
tri 910 3419 912 3421 ne
rect 924 3417 955 3435
rect 924 3407 970 3417
rect 1037 3446 1052 3461
tri 662 3382 674 3394 ne
rect 674 3389 684 3394
tri 684 3389 689 3394 sw
rect 573 3043 588 3271
rect 674 3281 689 3389
rect 728 3347 756 3403
tri 848 3385 866 3403 ne
rect 866 3383 888 3403
tri 888 3383 908 3403 sw
tri 924 3389 942 3407 ne
rect 747 3313 756 3347
rect 790 3374 832 3375
rect 790 3340 795 3374
rect 825 3340 832 3374
rect 790 3331 832 3340
rect 866 3374 908 3383
rect 866 3340 873 3374
rect 903 3340 908 3374
rect 866 3335 908 3340
rect 942 3347 970 3407
tri 1015 3394 1037 3416 se
rect 1037 3409 1052 3417
tri 1037 3394 1052 3409 nw
tri 1009 3388 1015 3394 se
rect 1015 3388 1024 3394
rect 728 3303 756 3313
tri 756 3303 780 3327 sw
rect 674 3233 690 3281
rect 728 3271 770 3303
tri 787 3295 788 3296 sw
rect 787 3271 788 3295
tri 790 3294 827 3331 ne
rect 827 3303 832 3331
tri 832 3303 858 3329 sw
rect 942 3313 951 3347
rect 942 3303 970 3313
rect 827 3294 911 3303
tri 827 3275 846 3294 ne
rect 846 3275 911 3294
rect 728 3249 788 3271
rect 910 3271 911 3275
rect 928 3271 970 3303
rect 910 3249 970 3271
rect 816 3233 833 3247
rect 865 3233 882 3247
tri 653 3197 675 3219 se
rect 675 3212 690 3233
tri 675 3197 690 3212 nw
rect 1009 3212 1024 3388
tri 1024 3381 1037 3394 nw
rect 1110 3313 1125 3541
tri 647 3191 653 3197 se
rect 653 3191 662 3197
rect 647 3175 662 3191
tri 662 3184 675 3197 nw
rect 816 3189 833 3203
rect 865 3189 882 3203
tri 1009 3197 1024 3212 ne
tri 1024 3197 1046 3219 sw
rect 647 3139 662 3147
rect 728 3175 788 3189
rect 743 3165 788 3175
rect 743 3147 771 3165
tri 647 3124 662 3139 ne
tri 662 3124 684 3146 sw
rect 728 3137 771 3147
rect 786 3161 788 3165
rect 910 3175 970 3189
tri 1024 3184 1037 3197 ne
rect 1037 3191 1046 3197
tri 1046 3191 1052 3197 sw
rect 910 3165 955 3175
rect 786 3137 860 3161
rect 728 3133 860 3137
tri 860 3133 888 3161 sw
rect 910 3151 912 3165
tri 910 3149 912 3151 ne
rect 924 3147 955 3165
rect 924 3137 970 3147
rect 1037 3176 1052 3191
tri 662 3112 674 3124 ne
rect 674 3119 684 3124
tri 684 3119 689 3124 sw
rect 573 2773 588 3001
rect 674 2963 689 3119
rect 728 3077 756 3133
tri 848 3115 866 3133 ne
rect 866 3113 888 3133
tri 888 3113 908 3133 sw
tri 924 3119 942 3137 ne
rect 747 3043 756 3077
rect 790 3104 832 3105
rect 790 3070 795 3104
rect 825 3070 832 3104
rect 790 3061 832 3070
rect 866 3104 908 3113
rect 866 3070 873 3104
rect 903 3070 908 3104
rect 866 3065 908 3070
rect 942 3077 970 3137
tri 1015 3124 1037 3146 se
rect 1037 3139 1052 3147
tri 1037 3124 1052 3139 nw
tri 1009 3118 1015 3124 se
rect 1015 3118 1024 3124
rect 728 3033 756 3043
tri 756 3033 780 3057 sw
rect 728 3001 770 3033
tri 787 3025 788 3026 sw
rect 787 3001 788 3025
tri 790 3024 827 3061 ne
rect 827 3033 832 3061
tri 832 3033 858 3059 sw
rect 942 3043 951 3077
rect 942 3033 970 3043
rect 827 3024 911 3033
tri 827 3005 846 3024 ne
rect 846 3005 911 3024
rect 728 2979 788 3001
rect 910 3001 911 3005
rect 928 3001 970 3033
rect 910 2979 970 3001
rect 816 2963 833 2977
rect 865 2963 882 2977
tri 653 2927 675 2949 se
rect 675 2942 690 2963
tri 675 2927 690 2942 nw
rect 1009 2942 1024 3118
tri 1024 3111 1037 3124 nw
rect 1110 3043 1125 3271
tri 647 2921 653 2927 se
rect 653 2921 662 2927
rect 647 2905 662 2921
tri 662 2914 675 2927 nw
rect 816 2919 833 2933
rect 865 2919 882 2933
tri 1009 2927 1024 2942 ne
tri 1024 2927 1046 2949 sw
rect 647 2869 662 2877
rect 728 2905 788 2919
rect 743 2895 788 2905
rect 743 2877 771 2895
tri 647 2854 662 2869 ne
tri 662 2854 684 2876 sw
rect 728 2867 771 2877
rect 786 2891 788 2895
rect 910 2905 970 2919
tri 1024 2914 1037 2927 ne
rect 1037 2921 1046 2927
tri 1046 2921 1052 2927 sw
rect 910 2895 955 2905
rect 786 2867 860 2891
rect 728 2863 860 2867
tri 860 2863 888 2891 sw
rect 910 2881 912 2895
tri 910 2879 912 2881 ne
rect 924 2877 955 2895
rect 924 2867 970 2877
rect 1037 2906 1052 2921
tri 662 2842 674 2854 ne
rect 674 2849 684 2854
tri 684 2849 689 2854 sw
rect 573 2503 588 2731
rect 674 2741 689 2849
rect 728 2807 756 2863
tri 848 2845 866 2863 ne
rect 866 2843 888 2863
tri 888 2843 908 2863 sw
tri 924 2849 942 2867 ne
rect 747 2773 756 2807
rect 790 2834 832 2835
rect 790 2800 795 2834
rect 825 2800 832 2834
rect 790 2791 832 2800
rect 866 2834 908 2843
rect 866 2800 873 2834
rect 903 2800 908 2834
rect 866 2795 908 2800
rect 942 2807 970 2867
tri 1015 2854 1037 2876 se
rect 1037 2869 1052 2877
tri 1037 2854 1052 2869 nw
tri 1009 2848 1015 2854 se
rect 1015 2848 1024 2854
rect 728 2763 756 2773
tri 756 2763 780 2787 sw
rect 674 2693 690 2741
rect 728 2731 770 2763
tri 787 2755 788 2756 sw
rect 787 2731 788 2755
tri 790 2754 827 2791 ne
rect 827 2763 832 2791
tri 832 2763 858 2789 sw
rect 942 2773 951 2807
rect 942 2763 970 2773
rect 827 2754 911 2763
tri 827 2735 846 2754 ne
rect 846 2735 911 2754
rect 728 2709 788 2731
rect 910 2731 911 2735
rect 928 2731 970 2763
rect 910 2709 970 2731
rect 816 2693 833 2707
rect 865 2693 882 2707
tri 653 2657 675 2679 se
rect 675 2672 690 2693
tri 675 2657 690 2672 nw
rect 1009 2672 1024 2848
tri 1024 2841 1037 2854 nw
rect 1110 2773 1125 3001
tri 647 2651 653 2657 se
rect 653 2651 662 2657
rect 647 2635 662 2651
tri 662 2644 675 2657 nw
rect 816 2649 833 2663
rect 865 2649 882 2663
tri 1009 2657 1024 2672 ne
tri 1024 2657 1046 2679 sw
rect 647 2599 662 2607
rect 728 2635 788 2649
rect 743 2625 788 2635
rect 743 2607 771 2625
tri 647 2584 662 2599 ne
tri 662 2584 684 2606 sw
rect 728 2597 771 2607
rect 786 2621 788 2625
rect 910 2635 970 2649
tri 1024 2644 1037 2657 ne
rect 1037 2651 1046 2657
tri 1046 2651 1052 2657 sw
rect 910 2625 955 2635
rect 786 2597 860 2621
rect 728 2593 860 2597
tri 860 2593 888 2621 sw
rect 910 2611 912 2625
tri 910 2609 912 2611 ne
rect 924 2607 955 2625
rect 924 2597 970 2607
rect 1037 2636 1052 2651
tri 662 2572 674 2584 ne
rect 674 2579 684 2584
tri 684 2579 689 2584 sw
rect 573 2233 588 2461
rect 674 2423 689 2579
rect 728 2537 756 2593
tri 848 2575 866 2593 ne
rect 866 2573 888 2593
tri 888 2573 908 2593 sw
tri 924 2579 942 2597 ne
rect 747 2503 756 2537
rect 790 2564 832 2565
rect 790 2530 795 2564
rect 825 2530 832 2564
rect 790 2521 832 2530
rect 866 2564 908 2573
rect 866 2530 873 2564
rect 903 2530 908 2564
rect 866 2525 908 2530
rect 942 2537 970 2597
tri 1015 2584 1037 2606 se
rect 1037 2599 1052 2607
tri 1037 2584 1052 2599 nw
tri 1009 2578 1015 2584 se
rect 1015 2578 1024 2584
rect 728 2493 756 2503
tri 756 2493 780 2517 sw
rect 728 2461 770 2493
tri 787 2485 788 2486 sw
rect 787 2461 788 2485
tri 790 2484 827 2521 ne
rect 827 2493 832 2521
tri 832 2493 858 2519 sw
rect 942 2503 951 2537
rect 942 2493 970 2503
rect 827 2484 911 2493
tri 827 2465 846 2484 ne
rect 846 2465 911 2484
rect 728 2439 788 2461
rect 910 2461 911 2465
rect 928 2461 970 2493
rect 910 2439 970 2461
rect 816 2423 833 2437
rect 865 2423 882 2437
tri 653 2387 675 2409 se
rect 675 2402 690 2423
tri 675 2387 690 2402 nw
rect 1009 2402 1024 2578
tri 1024 2571 1037 2584 nw
rect 1110 2503 1125 2731
tri 647 2381 653 2387 se
rect 653 2381 662 2387
rect 647 2365 662 2381
tri 662 2374 675 2387 nw
rect 816 2379 833 2393
rect 865 2379 882 2393
tri 1009 2387 1024 2402 ne
tri 1024 2387 1046 2409 sw
rect 647 2329 662 2337
rect 728 2365 788 2379
rect 743 2355 788 2365
rect 743 2337 771 2355
tri 647 2314 662 2329 ne
tri 662 2314 684 2336 sw
rect 728 2327 771 2337
rect 786 2351 788 2355
rect 910 2365 970 2379
tri 1024 2374 1037 2387 ne
rect 1037 2381 1046 2387
tri 1046 2381 1052 2387 sw
rect 910 2355 955 2365
rect 786 2327 860 2351
rect 728 2323 860 2327
tri 860 2323 888 2351 sw
rect 910 2341 912 2355
tri 910 2339 912 2341 ne
rect 924 2337 955 2355
rect 924 2327 970 2337
rect 1037 2366 1052 2381
tri 662 2302 674 2314 ne
rect 674 2309 684 2314
tri 684 2309 689 2314 sw
rect 573 1963 588 2191
rect 674 2201 689 2309
rect 728 2267 756 2323
tri 848 2305 866 2323 ne
rect 866 2303 888 2323
tri 888 2303 908 2323 sw
tri 924 2309 942 2327 ne
rect 747 2233 756 2267
rect 790 2294 832 2295
rect 790 2260 795 2294
rect 825 2260 832 2294
rect 790 2251 832 2260
rect 866 2294 908 2303
rect 866 2260 873 2294
rect 903 2260 908 2294
rect 866 2255 908 2260
rect 942 2267 970 2327
tri 1015 2314 1037 2336 se
rect 1037 2329 1052 2337
tri 1037 2314 1052 2329 nw
tri 1009 2308 1015 2314 se
rect 1015 2308 1024 2314
rect 728 2223 756 2233
tri 756 2223 780 2247 sw
rect 674 2153 690 2201
rect 728 2191 770 2223
tri 787 2215 788 2216 sw
rect 787 2191 788 2215
tri 790 2214 827 2251 ne
rect 827 2223 832 2251
tri 832 2223 858 2249 sw
rect 942 2233 951 2267
rect 942 2223 970 2233
rect 827 2214 911 2223
tri 827 2195 846 2214 ne
rect 846 2195 911 2214
rect 728 2169 788 2191
rect 910 2191 911 2195
rect 928 2191 970 2223
rect 910 2169 970 2191
rect 816 2153 833 2167
rect 865 2153 882 2167
tri 653 2117 675 2139 se
rect 675 2132 690 2153
tri 675 2117 690 2132 nw
rect 1009 2132 1024 2308
tri 1024 2301 1037 2314 nw
rect 1110 2233 1125 2461
tri 647 2111 653 2117 se
rect 653 2111 662 2117
rect 647 2095 662 2111
tri 662 2104 675 2117 nw
rect 816 2109 833 2123
rect 865 2109 882 2123
tri 1009 2117 1024 2132 ne
tri 1024 2117 1046 2139 sw
rect 647 2059 662 2067
rect 728 2095 788 2109
rect 743 2085 788 2095
rect 743 2067 771 2085
tri 647 2044 662 2059 ne
tri 662 2044 684 2066 sw
rect 728 2057 771 2067
rect 786 2081 788 2085
rect 910 2095 970 2109
tri 1024 2104 1037 2117 ne
rect 1037 2111 1046 2117
tri 1046 2111 1052 2117 sw
rect 910 2085 955 2095
rect 786 2057 860 2081
rect 728 2053 860 2057
tri 860 2053 888 2081 sw
rect 910 2071 912 2085
tri 910 2069 912 2071 ne
rect 924 2067 955 2085
rect 924 2057 970 2067
rect 1037 2096 1052 2111
tri 662 2032 674 2044 ne
rect 674 2039 684 2044
tri 684 2039 689 2044 sw
rect 573 1693 588 1921
rect 674 1883 689 2039
rect 728 1997 756 2053
tri 848 2035 866 2053 ne
rect 866 2033 888 2053
tri 888 2033 908 2053 sw
tri 924 2039 942 2057 ne
rect 747 1963 756 1997
rect 790 2024 832 2025
rect 790 1990 795 2024
rect 825 1990 832 2024
rect 790 1981 832 1990
rect 866 2024 908 2033
rect 866 1990 873 2024
rect 903 1990 908 2024
rect 866 1985 908 1990
rect 942 1997 970 2057
tri 1015 2044 1037 2066 se
rect 1037 2059 1052 2067
tri 1037 2044 1052 2059 nw
tri 1009 2038 1015 2044 se
rect 1015 2038 1024 2044
rect 728 1953 756 1963
tri 756 1953 780 1977 sw
rect 728 1921 770 1953
tri 787 1945 788 1946 sw
rect 787 1921 788 1945
tri 790 1944 827 1981 ne
rect 827 1953 832 1981
tri 832 1953 858 1979 sw
rect 942 1963 951 1997
rect 942 1953 970 1963
rect 827 1944 911 1953
tri 827 1925 846 1944 ne
rect 846 1925 911 1944
rect 728 1899 788 1921
rect 910 1921 911 1925
rect 928 1921 970 1953
rect 910 1899 970 1921
rect 816 1883 833 1897
rect 865 1883 882 1897
tri 653 1847 675 1869 se
rect 675 1862 690 1883
tri 675 1847 690 1862 nw
rect 1009 1862 1024 2038
tri 1024 2031 1037 2044 nw
rect 1110 1963 1125 2191
tri 647 1841 653 1847 se
rect 653 1841 662 1847
rect 647 1825 662 1841
tri 662 1834 675 1847 nw
rect 816 1839 833 1853
rect 865 1839 882 1853
tri 1009 1847 1024 1862 ne
tri 1024 1847 1046 1869 sw
rect 647 1789 662 1797
rect 728 1825 788 1839
rect 743 1815 788 1825
rect 743 1797 771 1815
tri 647 1774 662 1789 ne
tri 662 1774 684 1796 sw
rect 728 1787 771 1797
rect 786 1811 788 1815
rect 910 1825 970 1839
tri 1024 1834 1037 1847 ne
rect 1037 1841 1046 1847
tri 1046 1841 1052 1847 sw
rect 910 1815 955 1825
rect 786 1787 860 1811
rect 728 1783 860 1787
tri 860 1783 888 1811 sw
rect 910 1801 912 1815
tri 910 1799 912 1801 ne
rect 924 1797 955 1815
rect 924 1787 970 1797
rect 1037 1826 1052 1841
tri 662 1762 674 1774 ne
rect 674 1769 684 1774
tri 684 1769 689 1774 sw
rect 573 1423 588 1651
rect 674 1661 689 1769
rect 728 1727 756 1783
tri 848 1765 866 1783 ne
rect 866 1763 888 1783
tri 888 1763 908 1783 sw
tri 924 1769 942 1787 ne
rect 747 1693 756 1727
rect 790 1754 832 1755
rect 790 1720 795 1754
rect 825 1720 832 1754
rect 790 1711 832 1720
rect 866 1754 908 1763
rect 866 1720 873 1754
rect 903 1720 908 1754
rect 866 1715 908 1720
rect 942 1727 970 1787
tri 1015 1774 1037 1796 se
rect 1037 1789 1052 1797
tri 1037 1774 1052 1789 nw
tri 1009 1768 1015 1774 se
rect 1015 1768 1024 1774
rect 728 1683 756 1693
tri 756 1683 780 1707 sw
rect 674 1613 690 1661
rect 728 1651 770 1683
tri 787 1675 788 1676 sw
rect 787 1651 788 1675
tri 790 1674 827 1711 ne
rect 827 1683 832 1711
tri 832 1683 858 1709 sw
rect 942 1693 951 1727
rect 942 1683 970 1693
rect 827 1674 911 1683
tri 827 1655 846 1674 ne
rect 846 1655 911 1674
rect 728 1629 788 1651
rect 910 1651 911 1655
rect 928 1651 970 1683
rect 910 1629 970 1651
rect 816 1613 833 1627
rect 865 1613 882 1627
tri 653 1577 675 1599 se
rect 675 1592 690 1613
tri 675 1577 690 1592 nw
rect 1009 1592 1024 1768
tri 1024 1761 1037 1774 nw
rect 1110 1693 1125 1921
tri 647 1571 653 1577 se
rect 653 1571 662 1577
rect 647 1555 662 1571
tri 662 1564 675 1577 nw
rect 816 1569 833 1583
rect 865 1569 882 1583
tri 1009 1577 1024 1592 ne
tri 1024 1577 1046 1599 sw
rect 647 1519 662 1527
rect 728 1555 788 1569
rect 743 1545 788 1555
rect 743 1527 771 1545
tri 647 1504 662 1519 ne
tri 662 1504 684 1526 sw
rect 728 1517 771 1527
rect 786 1541 788 1545
rect 910 1555 970 1569
tri 1024 1564 1037 1577 ne
rect 1037 1571 1046 1577
tri 1046 1571 1052 1577 sw
rect 910 1545 955 1555
rect 786 1517 860 1541
rect 728 1513 860 1517
tri 860 1513 888 1541 sw
rect 910 1531 912 1545
tri 910 1529 912 1531 ne
rect 924 1527 955 1545
rect 924 1517 970 1527
rect 1037 1556 1052 1571
tri 662 1492 674 1504 ne
rect 674 1499 684 1504
tri 684 1499 689 1504 sw
rect 573 1153 588 1381
rect 674 1343 689 1499
rect 728 1457 756 1513
tri 848 1495 866 1513 ne
rect 866 1493 888 1513
tri 888 1493 908 1513 sw
tri 924 1499 942 1517 ne
rect 747 1423 756 1457
rect 790 1484 832 1485
rect 790 1450 795 1484
rect 825 1450 832 1484
rect 790 1441 832 1450
rect 866 1484 908 1493
rect 866 1450 873 1484
rect 903 1450 908 1484
rect 866 1445 908 1450
rect 942 1457 970 1517
tri 1015 1504 1037 1526 se
rect 1037 1519 1052 1527
tri 1037 1504 1052 1519 nw
tri 1009 1498 1015 1504 se
rect 1015 1498 1024 1504
rect 728 1413 756 1423
tri 756 1413 780 1437 sw
rect 728 1381 770 1413
tri 787 1405 788 1406 sw
rect 787 1381 788 1405
tri 790 1404 827 1441 ne
rect 827 1413 832 1441
tri 832 1413 858 1439 sw
rect 942 1423 951 1457
rect 942 1413 970 1423
rect 827 1404 911 1413
tri 827 1385 846 1404 ne
rect 846 1385 911 1404
rect 728 1359 788 1381
rect 910 1381 911 1385
rect 928 1381 970 1413
rect 910 1359 970 1381
rect 816 1343 833 1357
rect 865 1343 882 1357
tri 653 1307 675 1329 se
rect 675 1322 690 1343
tri 675 1307 690 1322 nw
rect 1009 1322 1024 1498
tri 1024 1491 1037 1504 nw
rect 1110 1423 1125 1651
tri 647 1301 653 1307 se
rect 653 1301 662 1307
rect 647 1285 662 1301
tri 662 1294 675 1307 nw
rect 816 1299 833 1313
rect 865 1299 882 1313
tri 1009 1307 1024 1322 ne
tri 1024 1307 1046 1329 sw
rect 647 1249 662 1257
rect 728 1285 788 1299
rect 743 1275 788 1285
rect 743 1257 771 1275
tri 647 1234 662 1249 ne
tri 662 1234 684 1256 sw
rect 728 1247 771 1257
rect 786 1271 788 1275
rect 910 1285 970 1299
tri 1024 1294 1037 1307 ne
rect 1037 1301 1046 1307
tri 1046 1301 1052 1307 sw
rect 910 1275 955 1285
rect 786 1247 860 1271
rect 728 1243 860 1247
tri 860 1243 888 1271 sw
rect 910 1261 912 1275
tri 910 1259 912 1261 ne
rect 924 1257 955 1275
rect 924 1247 970 1257
rect 1037 1286 1052 1301
tri 662 1222 674 1234 ne
rect 674 1229 684 1234
tri 684 1229 689 1234 sw
rect 573 883 588 1111
rect 674 1121 689 1229
rect 728 1187 756 1243
tri 848 1225 866 1243 ne
rect 866 1223 888 1243
tri 888 1223 908 1243 sw
tri 924 1229 942 1247 ne
rect 747 1153 756 1187
rect 790 1214 832 1215
rect 790 1180 795 1214
rect 825 1180 832 1214
rect 790 1171 832 1180
rect 866 1214 908 1223
rect 866 1180 873 1214
rect 903 1180 908 1214
rect 866 1175 908 1180
rect 942 1187 970 1247
tri 1015 1234 1037 1256 se
rect 1037 1249 1052 1257
tri 1037 1234 1052 1249 nw
tri 1009 1228 1015 1234 se
rect 1015 1228 1024 1234
rect 728 1143 756 1153
tri 756 1143 780 1167 sw
rect 674 1073 690 1121
rect 728 1111 770 1143
tri 787 1135 788 1136 sw
rect 787 1111 788 1135
tri 790 1134 827 1171 ne
rect 827 1143 832 1171
tri 832 1143 858 1169 sw
rect 942 1153 951 1187
rect 942 1143 970 1153
rect 827 1134 911 1143
tri 827 1115 846 1134 ne
rect 846 1115 911 1134
rect 728 1089 788 1111
rect 910 1111 911 1115
rect 928 1111 970 1143
rect 910 1089 970 1111
rect 816 1073 833 1087
rect 865 1073 882 1087
tri 653 1037 675 1059 se
rect 675 1052 690 1073
tri 675 1037 690 1052 nw
rect 1009 1052 1024 1228
tri 1024 1221 1037 1234 nw
rect 1110 1153 1125 1381
tri 647 1031 653 1037 se
rect 653 1031 662 1037
rect 647 1015 662 1031
tri 662 1024 675 1037 nw
rect 816 1029 833 1043
rect 865 1029 882 1043
tri 1009 1037 1024 1052 ne
tri 1024 1037 1046 1059 sw
rect 647 979 662 987
rect 728 1015 788 1029
rect 743 1005 788 1015
rect 743 987 771 1005
tri 647 964 662 979 ne
tri 662 964 684 986 sw
rect 728 977 771 987
rect 786 1001 788 1005
rect 910 1015 970 1029
tri 1024 1024 1037 1037 ne
rect 1037 1031 1046 1037
tri 1046 1031 1052 1037 sw
rect 910 1005 955 1015
rect 786 977 860 1001
rect 728 973 860 977
tri 860 973 888 1001 sw
rect 910 991 912 1005
tri 910 989 912 991 ne
rect 924 987 955 1005
rect 924 977 970 987
rect 1037 1016 1052 1031
tri 662 952 674 964 ne
rect 674 959 684 964
tri 684 959 689 964 sw
rect 573 613 588 841
rect 674 803 689 959
rect 728 917 756 973
tri 848 955 866 973 ne
rect 866 953 888 973
tri 888 953 908 973 sw
tri 924 959 942 977 ne
rect 747 883 756 917
rect 790 944 832 945
rect 790 910 795 944
rect 825 910 832 944
rect 790 901 832 910
rect 866 944 908 953
rect 866 910 873 944
rect 903 910 908 944
rect 866 905 908 910
rect 942 917 970 977
tri 1015 964 1037 986 se
rect 1037 979 1052 987
tri 1037 964 1052 979 nw
tri 1009 958 1015 964 se
rect 1015 958 1024 964
rect 728 873 756 883
tri 756 873 780 897 sw
rect 728 841 770 873
tri 787 865 788 866 sw
rect 787 841 788 865
tri 790 864 827 901 ne
rect 827 873 832 901
tri 832 873 858 899 sw
rect 942 883 951 917
rect 942 873 970 883
rect 827 864 911 873
tri 827 845 846 864 ne
rect 846 845 911 864
rect 728 819 788 841
rect 910 841 911 845
rect 928 841 970 873
rect 910 819 970 841
rect 816 803 833 817
rect 865 803 882 817
tri 653 767 675 789 se
rect 675 782 690 803
tri 675 767 690 782 nw
rect 1009 782 1024 958
tri 1024 951 1037 964 nw
rect 1110 883 1125 1111
tri 647 761 653 767 se
rect 653 761 662 767
rect 647 745 662 761
tri 662 754 675 767 nw
rect 816 759 833 773
rect 865 759 882 773
tri 1009 767 1024 782 ne
tri 1024 767 1046 789 sw
rect 647 709 662 717
rect 728 745 788 759
rect 743 735 788 745
rect 743 717 771 735
tri 647 694 662 709 ne
tri 662 694 684 716 sw
rect 728 707 771 717
rect 786 731 788 735
rect 910 745 970 759
tri 1024 754 1037 767 ne
rect 1037 761 1046 767
tri 1046 761 1052 767 sw
rect 910 735 955 745
rect 786 707 860 731
rect 728 703 860 707
tri 860 703 888 731 sw
rect 910 721 912 735
tri 910 719 912 721 ne
rect 924 717 955 735
rect 924 707 970 717
rect 1037 746 1052 761
tri 662 682 674 694 ne
rect 674 689 684 694
tri 684 689 689 694 sw
rect 573 343 588 571
rect 674 581 689 689
rect 728 647 756 703
tri 848 685 866 703 ne
rect 866 683 888 703
tri 888 683 908 703 sw
tri 924 689 942 707 ne
rect 747 613 756 647
rect 790 674 832 675
rect 790 640 795 674
rect 825 640 832 674
rect 790 631 832 640
rect 866 674 908 683
rect 866 640 873 674
rect 903 640 908 674
rect 866 635 908 640
rect 942 647 970 707
tri 1015 694 1037 716 se
rect 1037 709 1052 717
tri 1037 694 1052 709 nw
tri 1009 688 1015 694 se
rect 1015 688 1024 694
rect 728 603 756 613
tri 756 603 780 627 sw
rect 674 533 690 581
rect 728 571 770 603
tri 787 595 788 596 sw
rect 787 571 788 595
tri 790 594 827 631 ne
rect 827 603 832 631
tri 832 603 858 629 sw
rect 942 613 951 647
rect 942 603 970 613
rect 827 594 911 603
tri 827 575 846 594 ne
rect 846 575 911 594
rect 728 549 788 571
rect 910 571 911 575
rect 928 571 970 603
rect 910 549 970 571
rect 816 533 833 547
rect 865 533 882 547
tri 653 497 675 519 se
rect 675 512 690 533
tri 675 497 690 512 nw
rect 1009 512 1024 688
tri 1024 681 1037 694 nw
rect 1110 613 1125 841
tri 647 491 653 497 se
rect 653 491 662 497
rect 647 475 662 491
tri 662 484 675 497 nw
rect 816 489 833 503
rect 865 489 882 503
tri 1009 497 1024 512 ne
tri 1024 497 1046 519 sw
rect 647 439 662 447
rect 728 475 788 489
rect 743 465 788 475
rect 743 447 771 465
tri 647 424 662 439 ne
tri 662 424 684 446 sw
rect 728 437 771 447
rect 786 461 788 465
rect 910 475 970 489
tri 1024 484 1037 497 ne
rect 1037 491 1046 497
tri 1046 491 1052 497 sw
rect 910 465 955 475
rect 786 437 860 461
rect 728 433 860 437
tri 860 433 888 461 sw
rect 910 451 912 465
tri 910 449 912 451 ne
rect 924 447 955 465
rect 924 437 970 447
rect 1037 476 1052 491
tri 662 412 674 424 ne
rect 674 419 684 424
tri 684 419 689 424 sw
rect 573 73 588 301
rect 674 263 689 419
rect 728 377 756 433
tri 848 415 866 433 ne
rect 866 413 888 433
tri 888 413 908 433 sw
tri 924 419 942 437 ne
rect 747 343 756 377
rect 790 404 832 405
rect 790 370 795 404
rect 825 370 832 404
rect 790 361 832 370
rect 866 404 908 413
rect 866 370 873 404
rect 903 370 908 404
rect 866 365 908 370
rect 942 377 970 437
tri 1015 424 1037 446 se
rect 1037 439 1052 447
tri 1037 424 1052 439 nw
tri 1009 418 1015 424 se
rect 1015 418 1024 424
rect 728 333 756 343
tri 756 333 780 357 sw
rect 728 301 770 333
tri 787 325 788 326 sw
rect 787 301 788 325
tri 790 324 827 361 ne
rect 827 333 832 361
tri 832 333 858 359 sw
rect 942 343 951 377
rect 942 333 970 343
rect 827 324 911 333
tri 827 305 846 324 ne
rect 846 305 911 324
rect 728 279 788 301
rect 910 301 911 305
rect 928 301 970 333
rect 910 279 970 301
rect 816 263 833 277
rect 865 263 882 277
tri 653 227 675 249 se
rect 675 242 690 263
tri 675 227 690 242 nw
rect 1009 242 1024 418
tri 1024 411 1037 424 nw
rect 1110 343 1125 571
tri 647 221 653 227 se
rect 653 221 662 227
rect 647 205 662 221
tri 662 214 675 227 nw
rect 816 219 833 233
rect 865 219 882 233
tri 1009 227 1024 242 ne
tri 1024 227 1046 249 sw
rect 647 169 662 177
rect 728 205 788 219
rect 743 195 788 205
rect 743 177 771 195
tri 647 154 662 169 ne
tri 662 154 684 176 sw
rect 728 167 771 177
rect 786 191 788 195
rect 910 205 970 219
tri 1024 214 1037 227 ne
rect 1037 221 1046 227
tri 1046 221 1052 227 sw
rect 910 195 955 205
rect 786 167 860 191
rect 728 163 860 167
tri 860 163 888 191 sw
rect 910 181 912 195
tri 910 179 912 181 ne
rect 924 177 955 195
rect 924 167 970 177
rect 1037 206 1052 221
tri 662 142 674 154 ne
rect 674 149 684 154
tri 684 149 689 154 sw
rect 573 -55 588 31
rect 674 -55 689 149
rect 728 107 756 163
tri 848 145 866 163 ne
rect 866 143 888 163
tri 888 143 908 163 sw
tri 924 149 942 167 ne
rect 747 73 756 107
rect 790 134 832 135
rect 790 100 795 134
rect 825 100 832 134
rect 790 91 832 100
rect 866 134 908 143
rect 866 100 873 134
rect 903 100 908 134
rect 866 95 908 100
rect 942 107 970 167
tri 1015 154 1037 176 se
rect 1037 169 1052 177
tri 1037 154 1052 169 nw
tri 1009 148 1015 154 se
rect 1015 148 1024 154
rect 728 63 756 73
tri 756 63 780 87 sw
rect 728 31 770 63
tri 787 55 788 56 sw
rect 787 31 788 55
tri 790 54 827 91 ne
rect 827 63 832 91
tri 832 63 858 89 sw
rect 942 73 951 107
rect 942 63 970 73
rect 827 54 911 63
tri 827 35 846 54 ne
rect 846 35 911 54
rect 728 9 788 31
rect 910 31 911 35
rect 928 31 970 63
rect 910 9 970 31
rect 816 -7 833 7
rect 865 -7 882 7
rect 1009 -55 1024 148
tri 1024 141 1037 154 nw
rect 1110 73 1125 301
rect 1110 -55 1125 31
rect 1153 4123 1168 4361
tri 1233 4277 1255 4299 se
rect 1255 4292 1270 4361
tri 1255 4277 1270 4292 nw
rect 1589 4292 1604 4361
tri 1227 4271 1233 4277 se
rect 1233 4271 1242 4277
rect 1227 4255 1242 4271
tri 1242 4264 1255 4277 nw
rect 1396 4269 1413 4283
rect 1445 4269 1462 4283
tri 1589 4277 1604 4292 ne
tri 1604 4277 1626 4299 sw
rect 1227 4219 1242 4227
rect 1308 4255 1368 4269
rect 1323 4245 1368 4255
rect 1323 4227 1351 4245
tri 1227 4204 1242 4219 ne
tri 1242 4204 1264 4226 sw
rect 1308 4217 1351 4227
rect 1366 4241 1368 4245
rect 1490 4255 1550 4269
tri 1604 4264 1617 4277 ne
rect 1617 4271 1626 4277
tri 1626 4271 1632 4277 sw
rect 1490 4245 1535 4255
rect 1366 4217 1440 4241
rect 1308 4213 1440 4217
tri 1440 4213 1468 4241 sw
rect 1490 4231 1492 4245
tri 1490 4229 1492 4231 ne
rect 1504 4227 1535 4245
rect 1504 4217 1550 4227
rect 1617 4256 1632 4271
tri 1242 4192 1254 4204 ne
rect 1254 4199 1264 4204
tri 1264 4199 1269 4204 sw
rect 1153 3853 1168 4081
rect 1254 4043 1269 4199
rect 1308 4157 1336 4213
tri 1428 4195 1446 4213 ne
rect 1446 4193 1468 4213
tri 1468 4193 1488 4213 sw
tri 1504 4199 1522 4217 ne
rect 1327 4123 1336 4157
rect 1370 4184 1412 4185
rect 1370 4150 1375 4184
rect 1405 4150 1412 4184
rect 1370 4141 1412 4150
rect 1446 4184 1488 4193
rect 1446 4150 1453 4184
rect 1483 4150 1488 4184
rect 1446 4145 1488 4150
rect 1522 4157 1550 4217
tri 1595 4204 1617 4226 se
rect 1617 4219 1632 4227
tri 1617 4204 1632 4219 nw
tri 1589 4198 1595 4204 se
rect 1595 4198 1604 4204
rect 1308 4113 1336 4123
tri 1336 4113 1360 4137 sw
rect 1308 4081 1350 4113
tri 1367 4105 1368 4106 sw
rect 1367 4081 1368 4105
tri 1370 4104 1407 4141 ne
rect 1407 4113 1412 4141
tri 1412 4113 1438 4139 sw
rect 1522 4123 1531 4157
rect 1522 4113 1550 4123
rect 1407 4104 1491 4113
tri 1407 4085 1426 4104 ne
rect 1426 4085 1491 4104
rect 1308 4059 1368 4081
rect 1490 4081 1491 4085
rect 1508 4081 1550 4113
rect 1490 4059 1550 4081
rect 1396 4043 1413 4057
rect 1445 4043 1462 4057
tri 1233 4007 1255 4029 se
rect 1255 4022 1270 4043
tri 1255 4007 1270 4022 nw
rect 1589 4022 1604 4198
tri 1604 4191 1617 4204 nw
rect 1690 4123 1705 4361
tri 1227 4001 1233 4007 se
rect 1233 4001 1242 4007
rect 1227 3985 1242 4001
tri 1242 3994 1255 4007 nw
rect 1396 3999 1413 4013
rect 1445 3999 1462 4013
tri 1589 4007 1604 4022 ne
tri 1604 4007 1626 4029 sw
rect 1227 3949 1242 3957
rect 1308 3985 1368 3999
rect 1323 3975 1368 3985
rect 1323 3957 1351 3975
tri 1227 3934 1242 3949 ne
tri 1242 3934 1264 3956 sw
rect 1308 3947 1351 3957
rect 1366 3971 1368 3975
rect 1490 3985 1550 3999
tri 1604 3994 1617 4007 ne
rect 1617 4001 1626 4007
tri 1626 4001 1632 4007 sw
rect 1490 3975 1535 3985
rect 1366 3947 1440 3971
rect 1308 3943 1440 3947
tri 1440 3943 1468 3971 sw
rect 1490 3961 1492 3975
tri 1490 3959 1492 3961 ne
rect 1504 3957 1535 3975
rect 1504 3947 1550 3957
rect 1617 3986 1632 4001
tri 1242 3922 1254 3934 ne
rect 1254 3929 1264 3934
tri 1264 3929 1269 3934 sw
rect 1153 3583 1168 3811
rect 1254 3821 1269 3929
rect 1308 3887 1336 3943
tri 1428 3925 1446 3943 ne
rect 1446 3923 1468 3943
tri 1468 3923 1488 3943 sw
tri 1504 3929 1522 3947 ne
rect 1327 3853 1336 3887
rect 1370 3914 1412 3915
rect 1370 3880 1375 3914
rect 1405 3880 1412 3914
rect 1370 3871 1412 3880
rect 1446 3914 1488 3923
rect 1446 3880 1453 3914
rect 1483 3880 1488 3914
rect 1446 3875 1488 3880
rect 1522 3887 1550 3947
tri 1595 3934 1617 3956 se
rect 1617 3949 1632 3957
tri 1617 3934 1632 3949 nw
tri 1589 3928 1595 3934 se
rect 1595 3928 1604 3934
rect 1308 3843 1336 3853
tri 1336 3843 1360 3867 sw
rect 1254 3773 1270 3821
rect 1308 3811 1350 3843
tri 1367 3835 1368 3836 sw
rect 1367 3811 1368 3835
tri 1370 3834 1407 3871 ne
rect 1407 3843 1412 3871
tri 1412 3843 1438 3869 sw
rect 1522 3853 1531 3887
rect 1522 3843 1550 3853
rect 1407 3834 1491 3843
tri 1407 3815 1426 3834 ne
rect 1426 3815 1491 3834
rect 1308 3789 1368 3811
rect 1490 3811 1491 3815
rect 1508 3811 1550 3843
rect 1490 3789 1550 3811
rect 1396 3773 1413 3787
rect 1445 3773 1462 3787
tri 1233 3737 1255 3759 se
rect 1255 3752 1270 3773
tri 1255 3737 1270 3752 nw
rect 1589 3752 1604 3928
tri 1604 3921 1617 3934 nw
rect 1690 3853 1705 4081
tri 1227 3731 1233 3737 se
rect 1233 3731 1242 3737
rect 1227 3715 1242 3731
tri 1242 3724 1255 3737 nw
rect 1396 3729 1413 3743
rect 1445 3729 1462 3743
tri 1589 3737 1604 3752 ne
tri 1604 3737 1626 3759 sw
rect 1227 3679 1242 3687
rect 1308 3715 1368 3729
rect 1323 3705 1368 3715
rect 1323 3687 1351 3705
tri 1227 3664 1242 3679 ne
tri 1242 3664 1264 3686 sw
rect 1308 3677 1351 3687
rect 1366 3701 1368 3705
rect 1490 3715 1550 3729
tri 1604 3724 1617 3737 ne
rect 1617 3731 1626 3737
tri 1626 3731 1632 3737 sw
rect 1490 3705 1535 3715
rect 1366 3677 1440 3701
rect 1308 3673 1440 3677
tri 1440 3673 1468 3701 sw
rect 1490 3691 1492 3705
tri 1490 3689 1492 3691 ne
rect 1504 3687 1535 3705
rect 1504 3677 1550 3687
rect 1617 3716 1632 3731
tri 1242 3652 1254 3664 ne
rect 1254 3659 1264 3664
tri 1264 3659 1269 3664 sw
rect 1153 3313 1168 3541
rect 1254 3503 1269 3659
rect 1308 3617 1336 3673
tri 1428 3655 1446 3673 ne
rect 1446 3653 1468 3673
tri 1468 3653 1488 3673 sw
tri 1504 3659 1522 3677 ne
rect 1327 3583 1336 3617
rect 1370 3644 1412 3645
rect 1370 3610 1375 3644
rect 1405 3610 1412 3644
rect 1370 3601 1412 3610
rect 1446 3644 1488 3653
rect 1446 3610 1453 3644
rect 1483 3610 1488 3644
rect 1446 3605 1488 3610
rect 1522 3617 1550 3677
tri 1595 3664 1617 3686 se
rect 1617 3679 1632 3687
tri 1617 3664 1632 3679 nw
tri 1589 3658 1595 3664 se
rect 1595 3658 1604 3664
rect 1308 3573 1336 3583
tri 1336 3573 1360 3597 sw
rect 1308 3541 1350 3573
tri 1367 3565 1368 3566 sw
rect 1367 3541 1368 3565
tri 1370 3564 1407 3601 ne
rect 1407 3573 1412 3601
tri 1412 3573 1438 3599 sw
rect 1522 3583 1531 3617
rect 1522 3573 1550 3583
rect 1407 3564 1491 3573
tri 1407 3545 1426 3564 ne
rect 1426 3545 1491 3564
rect 1308 3519 1368 3541
rect 1490 3541 1491 3545
rect 1508 3541 1550 3573
rect 1490 3519 1550 3541
rect 1396 3503 1413 3517
rect 1445 3503 1462 3517
tri 1233 3467 1255 3489 se
rect 1255 3482 1270 3503
tri 1255 3467 1270 3482 nw
rect 1589 3482 1604 3658
tri 1604 3651 1617 3664 nw
rect 1690 3583 1705 3811
tri 1227 3461 1233 3467 se
rect 1233 3461 1242 3467
rect 1227 3445 1242 3461
tri 1242 3454 1255 3467 nw
rect 1396 3459 1413 3473
rect 1445 3459 1462 3473
tri 1589 3467 1604 3482 ne
tri 1604 3467 1626 3489 sw
rect 1227 3409 1242 3417
rect 1308 3445 1368 3459
rect 1323 3435 1368 3445
rect 1323 3417 1351 3435
tri 1227 3394 1242 3409 ne
tri 1242 3394 1264 3416 sw
rect 1308 3407 1351 3417
rect 1366 3431 1368 3435
rect 1490 3445 1550 3459
tri 1604 3454 1617 3467 ne
rect 1617 3461 1626 3467
tri 1626 3461 1632 3467 sw
rect 1490 3435 1535 3445
rect 1366 3407 1440 3431
rect 1308 3403 1440 3407
tri 1440 3403 1468 3431 sw
rect 1490 3421 1492 3435
tri 1490 3419 1492 3421 ne
rect 1504 3417 1535 3435
rect 1504 3407 1550 3417
rect 1617 3446 1632 3461
tri 1242 3382 1254 3394 ne
rect 1254 3389 1264 3394
tri 1264 3389 1269 3394 sw
rect 1153 3043 1168 3271
rect 1254 3281 1269 3389
rect 1308 3347 1336 3403
tri 1428 3385 1446 3403 ne
rect 1446 3383 1468 3403
tri 1468 3383 1488 3403 sw
tri 1504 3389 1522 3407 ne
rect 1327 3313 1336 3347
rect 1370 3374 1412 3375
rect 1370 3340 1375 3374
rect 1405 3340 1412 3374
rect 1370 3331 1412 3340
rect 1446 3374 1488 3383
rect 1446 3340 1453 3374
rect 1483 3340 1488 3374
rect 1446 3335 1488 3340
rect 1522 3347 1550 3407
tri 1595 3394 1617 3416 se
rect 1617 3409 1632 3417
tri 1617 3394 1632 3409 nw
tri 1589 3388 1595 3394 se
rect 1595 3388 1604 3394
rect 1308 3303 1336 3313
tri 1336 3303 1360 3327 sw
rect 1254 3233 1270 3281
rect 1308 3271 1350 3303
tri 1367 3295 1368 3296 sw
rect 1367 3271 1368 3295
tri 1370 3294 1407 3331 ne
rect 1407 3303 1412 3331
tri 1412 3303 1438 3329 sw
rect 1522 3313 1531 3347
rect 1522 3303 1550 3313
rect 1407 3294 1491 3303
tri 1407 3275 1426 3294 ne
rect 1426 3275 1491 3294
rect 1308 3249 1368 3271
rect 1490 3271 1491 3275
rect 1508 3271 1550 3303
rect 1490 3249 1550 3271
rect 1396 3233 1413 3247
rect 1445 3233 1462 3247
tri 1233 3197 1255 3219 se
rect 1255 3212 1270 3233
tri 1255 3197 1270 3212 nw
rect 1589 3212 1604 3388
tri 1604 3381 1617 3394 nw
rect 1690 3313 1705 3541
tri 1227 3191 1233 3197 se
rect 1233 3191 1242 3197
rect 1227 3175 1242 3191
tri 1242 3184 1255 3197 nw
rect 1396 3189 1413 3203
rect 1445 3189 1462 3203
tri 1589 3197 1604 3212 ne
tri 1604 3197 1626 3219 sw
rect 1227 3139 1242 3147
rect 1308 3175 1368 3189
rect 1323 3165 1368 3175
rect 1323 3147 1351 3165
tri 1227 3124 1242 3139 ne
tri 1242 3124 1264 3146 sw
rect 1308 3137 1351 3147
rect 1366 3161 1368 3165
rect 1490 3175 1550 3189
tri 1604 3184 1617 3197 ne
rect 1617 3191 1626 3197
tri 1626 3191 1632 3197 sw
rect 1490 3165 1535 3175
rect 1366 3137 1440 3161
rect 1308 3133 1440 3137
tri 1440 3133 1468 3161 sw
rect 1490 3151 1492 3165
tri 1490 3149 1492 3151 ne
rect 1504 3147 1535 3165
rect 1504 3137 1550 3147
rect 1617 3176 1632 3191
tri 1242 3112 1254 3124 ne
rect 1254 3119 1264 3124
tri 1264 3119 1269 3124 sw
rect 1153 2773 1168 3001
rect 1254 2963 1269 3119
rect 1308 3077 1336 3133
tri 1428 3115 1446 3133 ne
rect 1446 3113 1468 3133
tri 1468 3113 1488 3133 sw
tri 1504 3119 1522 3137 ne
rect 1327 3043 1336 3077
rect 1370 3104 1412 3105
rect 1370 3070 1375 3104
rect 1405 3070 1412 3104
rect 1370 3061 1412 3070
rect 1446 3104 1488 3113
rect 1446 3070 1453 3104
rect 1483 3070 1488 3104
rect 1446 3065 1488 3070
rect 1522 3077 1550 3137
tri 1595 3124 1617 3146 se
rect 1617 3139 1632 3147
tri 1617 3124 1632 3139 nw
tri 1589 3118 1595 3124 se
rect 1595 3118 1604 3124
rect 1308 3033 1336 3043
tri 1336 3033 1360 3057 sw
rect 1308 3001 1350 3033
tri 1367 3025 1368 3026 sw
rect 1367 3001 1368 3025
tri 1370 3024 1407 3061 ne
rect 1407 3033 1412 3061
tri 1412 3033 1438 3059 sw
rect 1522 3043 1531 3077
rect 1522 3033 1550 3043
rect 1407 3024 1491 3033
tri 1407 3005 1426 3024 ne
rect 1426 3005 1491 3024
rect 1308 2979 1368 3001
rect 1490 3001 1491 3005
rect 1508 3001 1550 3033
rect 1490 2979 1550 3001
rect 1396 2963 1413 2977
rect 1445 2963 1462 2977
tri 1233 2927 1255 2949 se
rect 1255 2942 1270 2963
tri 1255 2927 1270 2942 nw
rect 1589 2942 1604 3118
tri 1604 3111 1617 3124 nw
rect 1690 3043 1705 3271
tri 1227 2921 1233 2927 se
rect 1233 2921 1242 2927
rect 1227 2905 1242 2921
tri 1242 2914 1255 2927 nw
rect 1396 2919 1413 2933
rect 1445 2919 1462 2933
tri 1589 2927 1604 2942 ne
tri 1604 2927 1626 2949 sw
rect 1227 2869 1242 2877
rect 1308 2905 1368 2919
rect 1323 2895 1368 2905
rect 1323 2877 1351 2895
tri 1227 2854 1242 2869 ne
tri 1242 2854 1264 2876 sw
rect 1308 2867 1351 2877
rect 1366 2891 1368 2895
rect 1490 2905 1550 2919
tri 1604 2914 1617 2927 ne
rect 1617 2921 1626 2927
tri 1626 2921 1632 2927 sw
rect 1490 2895 1535 2905
rect 1366 2867 1440 2891
rect 1308 2863 1440 2867
tri 1440 2863 1468 2891 sw
rect 1490 2881 1492 2895
tri 1490 2879 1492 2881 ne
rect 1504 2877 1535 2895
rect 1504 2867 1550 2877
rect 1617 2906 1632 2921
tri 1242 2842 1254 2854 ne
rect 1254 2849 1264 2854
tri 1264 2849 1269 2854 sw
rect 1153 2503 1168 2731
rect 1254 2741 1269 2849
rect 1308 2807 1336 2863
tri 1428 2845 1446 2863 ne
rect 1446 2843 1468 2863
tri 1468 2843 1488 2863 sw
tri 1504 2849 1522 2867 ne
rect 1327 2773 1336 2807
rect 1370 2834 1412 2835
rect 1370 2800 1375 2834
rect 1405 2800 1412 2834
rect 1370 2791 1412 2800
rect 1446 2834 1488 2843
rect 1446 2800 1453 2834
rect 1483 2800 1488 2834
rect 1446 2795 1488 2800
rect 1522 2807 1550 2867
tri 1595 2854 1617 2876 se
rect 1617 2869 1632 2877
tri 1617 2854 1632 2869 nw
tri 1589 2848 1595 2854 se
rect 1595 2848 1604 2854
rect 1308 2763 1336 2773
tri 1336 2763 1360 2787 sw
rect 1254 2693 1270 2741
rect 1308 2731 1350 2763
tri 1367 2755 1368 2756 sw
rect 1367 2731 1368 2755
tri 1370 2754 1407 2791 ne
rect 1407 2763 1412 2791
tri 1412 2763 1438 2789 sw
rect 1522 2773 1531 2807
rect 1522 2763 1550 2773
rect 1407 2754 1491 2763
tri 1407 2735 1426 2754 ne
rect 1426 2735 1491 2754
rect 1308 2709 1368 2731
rect 1490 2731 1491 2735
rect 1508 2731 1550 2763
rect 1490 2709 1550 2731
rect 1396 2693 1413 2707
rect 1445 2693 1462 2707
tri 1233 2657 1255 2679 se
rect 1255 2672 1270 2693
tri 1255 2657 1270 2672 nw
rect 1589 2672 1604 2848
tri 1604 2841 1617 2854 nw
rect 1690 2773 1705 3001
tri 1227 2651 1233 2657 se
rect 1233 2651 1242 2657
rect 1227 2635 1242 2651
tri 1242 2644 1255 2657 nw
rect 1396 2649 1413 2663
rect 1445 2649 1462 2663
tri 1589 2657 1604 2672 ne
tri 1604 2657 1626 2679 sw
rect 1227 2599 1242 2607
rect 1308 2635 1368 2649
rect 1323 2625 1368 2635
rect 1323 2607 1351 2625
tri 1227 2584 1242 2599 ne
tri 1242 2584 1264 2606 sw
rect 1308 2597 1351 2607
rect 1366 2621 1368 2625
rect 1490 2635 1550 2649
tri 1604 2644 1617 2657 ne
rect 1617 2651 1626 2657
tri 1626 2651 1632 2657 sw
rect 1490 2625 1535 2635
rect 1366 2597 1440 2621
rect 1308 2593 1440 2597
tri 1440 2593 1468 2621 sw
rect 1490 2611 1492 2625
tri 1490 2609 1492 2611 ne
rect 1504 2607 1535 2625
rect 1504 2597 1550 2607
rect 1617 2636 1632 2651
tri 1242 2572 1254 2584 ne
rect 1254 2579 1264 2584
tri 1264 2579 1269 2584 sw
rect 1153 2233 1168 2461
rect 1254 2423 1269 2579
rect 1308 2537 1336 2593
tri 1428 2575 1446 2593 ne
rect 1446 2573 1468 2593
tri 1468 2573 1488 2593 sw
tri 1504 2579 1522 2597 ne
rect 1327 2503 1336 2537
rect 1370 2564 1412 2565
rect 1370 2530 1375 2564
rect 1405 2530 1412 2564
rect 1370 2521 1412 2530
rect 1446 2564 1488 2573
rect 1446 2530 1453 2564
rect 1483 2530 1488 2564
rect 1446 2525 1488 2530
rect 1522 2537 1550 2597
tri 1595 2584 1617 2606 se
rect 1617 2599 1632 2607
tri 1617 2584 1632 2599 nw
tri 1589 2578 1595 2584 se
rect 1595 2578 1604 2584
rect 1308 2493 1336 2503
tri 1336 2493 1360 2517 sw
rect 1308 2461 1350 2493
tri 1367 2485 1368 2486 sw
rect 1367 2461 1368 2485
tri 1370 2484 1407 2521 ne
rect 1407 2493 1412 2521
tri 1412 2493 1438 2519 sw
rect 1522 2503 1531 2537
rect 1522 2493 1550 2503
rect 1407 2484 1491 2493
tri 1407 2465 1426 2484 ne
rect 1426 2465 1491 2484
rect 1308 2439 1368 2461
rect 1490 2461 1491 2465
rect 1508 2461 1550 2493
rect 1490 2439 1550 2461
rect 1396 2423 1413 2437
rect 1445 2423 1462 2437
tri 1233 2387 1255 2409 se
rect 1255 2402 1270 2423
tri 1255 2387 1270 2402 nw
rect 1589 2402 1604 2578
tri 1604 2571 1617 2584 nw
rect 1690 2503 1705 2731
tri 1227 2381 1233 2387 se
rect 1233 2381 1242 2387
rect 1227 2365 1242 2381
tri 1242 2374 1255 2387 nw
rect 1396 2379 1413 2393
rect 1445 2379 1462 2393
tri 1589 2387 1604 2402 ne
tri 1604 2387 1626 2409 sw
rect 1227 2329 1242 2337
rect 1308 2365 1368 2379
rect 1323 2355 1368 2365
rect 1323 2337 1351 2355
tri 1227 2314 1242 2329 ne
tri 1242 2314 1264 2336 sw
rect 1308 2327 1351 2337
rect 1366 2351 1368 2355
rect 1490 2365 1550 2379
tri 1604 2374 1617 2387 ne
rect 1617 2381 1626 2387
tri 1626 2381 1632 2387 sw
rect 1490 2355 1535 2365
rect 1366 2327 1440 2351
rect 1308 2323 1440 2327
tri 1440 2323 1468 2351 sw
rect 1490 2341 1492 2355
tri 1490 2339 1492 2341 ne
rect 1504 2337 1535 2355
rect 1504 2327 1550 2337
rect 1617 2366 1632 2381
tri 1242 2302 1254 2314 ne
rect 1254 2309 1264 2314
tri 1264 2309 1269 2314 sw
rect 1153 1963 1168 2191
rect 1254 2201 1269 2309
rect 1308 2267 1336 2323
tri 1428 2305 1446 2323 ne
rect 1446 2303 1468 2323
tri 1468 2303 1488 2323 sw
tri 1504 2309 1522 2327 ne
rect 1327 2233 1336 2267
rect 1370 2294 1412 2295
rect 1370 2260 1375 2294
rect 1405 2260 1412 2294
rect 1370 2251 1412 2260
rect 1446 2294 1488 2303
rect 1446 2260 1453 2294
rect 1483 2260 1488 2294
rect 1446 2255 1488 2260
rect 1522 2267 1550 2327
tri 1595 2314 1617 2336 se
rect 1617 2329 1632 2337
tri 1617 2314 1632 2329 nw
tri 1589 2308 1595 2314 se
rect 1595 2308 1604 2314
rect 1308 2223 1336 2233
tri 1336 2223 1360 2247 sw
rect 1254 2153 1270 2201
rect 1308 2191 1350 2223
tri 1367 2215 1368 2216 sw
rect 1367 2191 1368 2215
tri 1370 2214 1407 2251 ne
rect 1407 2223 1412 2251
tri 1412 2223 1438 2249 sw
rect 1522 2233 1531 2267
rect 1522 2223 1550 2233
rect 1407 2214 1491 2223
tri 1407 2195 1426 2214 ne
rect 1426 2195 1491 2214
rect 1308 2169 1368 2191
rect 1490 2191 1491 2195
rect 1508 2191 1550 2223
rect 1490 2169 1550 2191
rect 1396 2153 1413 2167
rect 1445 2153 1462 2167
tri 1233 2117 1255 2139 se
rect 1255 2132 1270 2153
tri 1255 2117 1270 2132 nw
rect 1589 2132 1604 2308
tri 1604 2301 1617 2314 nw
rect 1690 2233 1705 2461
tri 1227 2111 1233 2117 se
rect 1233 2111 1242 2117
rect 1227 2095 1242 2111
tri 1242 2104 1255 2117 nw
rect 1396 2109 1413 2123
rect 1445 2109 1462 2123
tri 1589 2117 1604 2132 ne
tri 1604 2117 1626 2139 sw
rect 1227 2059 1242 2067
rect 1308 2095 1368 2109
rect 1323 2085 1368 2095
rect 1323 2067 1351 2085
tri 1227 2044 1242 2059 ne
tri 1242 2044 1264 2066 sw
rect 1308 2057 1351 2067
rect 1366 2081 1368 2085
rect 1490 2095 1550 2109
tri 1604 2104 1617 2117 ne
rect 1617 2111 1626 2117
tri 1626 2111 1632 2117 sw
rect 1490 2085 1535 2095
rect 1366 2057 1440 2081
rect 1308 2053 1440 2057
tri 1440 2053 1468 2081 sw
rect 1490 2071 1492 2085
tri 1490 2069 1492 2071 ne
rect 1504 2067 1535 2085
rect 1504 2057 1550 2067
rect 1617 2096 1632 2111
tri 1242 2032 1254 2044 ne
rect 1254 2039 1264 2044
tri 1264 2039 1269 2044 sw
rect 1153 1693 1168 1921
rect 1254 1883 1269 2039
rect 1308 1997 1336 2053
tri 1428 2035 1446 2053 ne
rect 1446 2033 1468 2053
tri 1468 2033 1488 2053 sw
tri 1504 2039 1522 2057 ne
rect 1327 1963 1336 1997
rect 1370 2024 1412 2025
rect 1370 1990 1375 2024
rect 1405 1990 1412 2024
rect 1370 1981 1412 1990
rect 1446 2024 1488 2033
rect 1446 1990 1453 2024
rect 1483 1990 1488 2024
rect 1446 1985 1488 1990
rect 1522 1997 1550 2057
tri 1595 2044 1617 2066 se
rect 1617 2059 1632 2067
tri 1617 2044 1632 2059 nw
tri 1589 2038 1595 2044 se
rect 1595 2038 1604 2044
rect 1308 1953 1336 1963
tri 1336 1953 1360 1977 sw
rect 1308 1921 1350 1953
tri 1367 1945 1368 1946 sw
rect 1367 1921 1368 1945
tri 1370 1944 1407 1981 ne
rect 1407 1953 1412 1981
tri 1412 1953 1438 1979 sw
rect 1522 1963 1531 1997
rect 1522 1953 1550 1963
rect 1407 1944 1491 1953
tri 1407 1925 1426 1944 ne
rect 1426 1925 1491 1944
rect 1308 1899 1368 1921
rect 1490 1921 1491 1925
rect 1508 1921 1550 1953
rect 1490 1899 1550 1921
rect 1396 1883 1413 1897
rect 1445 1883 1462 1897
tri 1233 1847 1255 1869 se
rect 1255 1862 1270 1883
tri 1255 1847 1270 1862 nw
rect 1589 1862 1604 2038
tri 1604 2031 1617 2044 nw
rect 1690 1963 1705 2191
tri 1227 1841 1233 1847 se
rect 1233 1841 1242 1847
rect 1227 1825 1242 1841
tri 1242 1834 1255 1847 nw
rect 1396 1839 1413 1853
rect 1445 1839 1462 1853
tri 1589 1847 1604 1862 ne
tri 1604 1847 1626 1869 sw
rect 1227 1789 1242 1797
rect 1308 1825 1368 1839
rect 1323 1815 1368 1825
rect 1323 1797 1351 1815
tri 1227 1774 1242 1789 ne
tri 1242 1774 1264 1796 sw
rect 1308 1787 1351 1797
rect 1366 1811 1368 1815
rect 1490 1825 1550 1839
tri 1604 1834 1617 1847 ne
rect 1617 1841 1626 1847
tri 1626 1841 1632 1847 sw
rect 1490 1815 1535 1825
rect 1366 1787 1440 1811
rect 1308 1783 1440 1787
tri 1440 1783 1468 1811 sw
rect 1490 1801 1492 1815
tri 1490 1799 1492 1801 ne
rect 1504 1797 1535 1815
rect 1504 1787 1550 1797
rect 1617 1826 1632 1841
tri 1242 1762 1254 1774 ne
rect 1254 1769 1264 1774
tri 1264 1769 1269 1774 sw
rect 1153 1423 1168 1651
rect 1254 1661 1269 1769
rect 1308 1727 1336 1783
tri 1428 1765 1446 1783 ne
rect 1446 1763 1468 1783
tri 1468 1763 1488 1783 sw
tri 1504 1769 1522 1787 ne
rect 1327 1693 1336 1727
rect 1370 1754 1412 1755
rect 1370 1720 1375 1754
rect 1405 1720 1412 1754
rect 1370 1711 1412 1720
rect 1446 1754 1488 1763
rect 1446 1720 1453 1754
rect 1483 1720 1488 1754
rect 1446 1715 1488 1720
rect 1522 1727 1550 1787
tri 1595 1774 1617 1796 se
rect 1617 1789 1632 1797
tri 1617 1774 1632 1789 nw
tri 1589 1768 1595 1774 se
rect 1595 1768 1604 1774
rect 1308 1683 1336 1693
tri 1336 1683 1360 1707 sw
rect 1254 1613 1270 1661
rect 1308 1651 1350 1683
tri 1367 1675 1368 1676 sw
rect 1367 1651 1368 1675
tri 1370 1674 1407 1711 ne
rect 1407 1683 1412 1711
tri 1412 1683 1438 1709 sw
rect 1522 1693 1531 1727
rect 1522 1683 1550 1693
rect 1407 1674 1491 1683
tri 1407 1655 1426 1674 ne
rect 1426 1655 1491 1674
rect 1308 1629 1368 1651
rect 1490 1651 1491 1655
rect 1508 1651 1550 1683
rect 1490 1629 1550 1651
rect 1396 1613 1413 1627
rect 1445 1613 1462 1627
tri 1233 1577 1255 1599 se
rect 1255 1592 1270 1613
tri 1255 1577 1270 1592 nw
rect 1589 1592 1604 1768
tri 1604 1761 1617 1774 nw
rect 1690 1693 1705 1921
tri 1227 1571 1233 1577 se
rect 1233 1571 1242 1577
rect 1227 1555 1242 1571
tri 1242 1564 1255 1577 nw
rect 1396 1569 1413 1583
rect 1445 1569 1462 1583
tri 1589 1577 1604 1592 ne
tri 1604 1577 1626 1599 sw
rect 1227 1519 1242 1527
rect 1308 1555 1368 1569
rect 1323 1545 1368 1555
rect 1323 1527 1351 1545
tri 1227 1504 1242 1519 ne
tri 1242 1504 1264 1526 sw
rect 1308 1517 1351 1527
rect 1366 1541 1368 1545
rect 1490 1555 1550 1569
tri 1604 1564 1617 1577 ne
rect 1617 1571 1626 1577
tri 1626 1571 1632 1577 sw
rect 1490 1545 1535 1555
rect 1366 1517 1440 1541
rect 1308 1513 1440 1517
tri 1440 1513 1468 1541 sw
rect 1490 1531 1492 1545
tri 1490 1529 1492 1531 ne
rect 1504 1527 1535 1545
rect 1504 1517 1550 1527
rect 1617 1556 1632 1571
tri 1242 1492 1254 1504 ne
rect 1254 1499 1264 1504
tri 1264 1499 1269 1504 sw
rect 1153 1153 1168 1381
rect 1254 1343 1269 1499
rect 1308 1457 1336 1513
tri 1428 1495 1446 1513 ne
rect 1446 1493 1468 1513
tri 1468 1493 1488 1513 sw
tri 1504 1499 1522 1517 ne
rect 1327 1423 1336 1457
rect 1370 1484 1412 1485
rect 1370 1450 1375 1484
rect 1405 1450 1412 1484
rect 1370 1441 1412 1450
rect 1446 1484 1488 1493
rect 1446 1450 1453 1484
rect 1483 1450 1488 1484
rect 1446 1445 1488 1450
rect 1522 1457 1550 1517
tri 1595 1504 1617 1526 se
rect 1617 1519 1632 1527
tri 1617 1504 1632 1519 nw
tri 1589 1498 1595 1504 se
rect 1595 1498 1604 1504
rect 1308 1413 1336 1423
tri 1336 1413 1360 1437 sw
rect 1308 1381 1350 1413
tri 1367 1405 1368 1406 sw
rect 1367 1381 1368 1405
tri 1370 1404 1407 1441 ne
rect 1407 1413 1412 1441
tri 1412 1413 1438 1439 sw
rect 1522 1423 1531 1457
rect 1522 1413 1550 1423
rect 1407 1404 1491 1413
tri 1407 1385 1426 1404 ne
rect 1426 1385 1491 1404
rect 1308 1359 1368 1381
rect 1490 1381 1491 1385
rect 1508 1381 1550 1413
rect 1490 1359 1550 1381
rect 1396 1343 1413 1357
rect 1445 1343 1462 1357
tri 1233 1307 1255 1329 se
rect 1255 1322 1270 1343
tri 1255 1307 1270 1322 nw
rect 1589 1322 1604 1498
tri 1604 1491 1617 1504 nw
rect 1690 1423 1705 1651
tri 1227 1301 1233 1307 se
rect 1233 1301 1242 1307
rect 1227 1285 1242 1301
tri 1242 1294 1255 1307 nw
rect 1396 1299 1413 1313
rect 1445 1299 1462 1313
tri 1589 1307 1604 1322 ne
tri 1604 1307 1626 1329 sw
rect 1227 1249 1242 1257
rect 1308 1285 1368 1299
rect 1323 1275 1368 1285
rect 1323 1257 1351 1275
tri 1227 1234 1242 1249 ne
tri 1242 1234 1264 1256 sw
rect 1308 1247 1351 1257
rect 1366 1271 1368 1275
rect 1490 1285 1550 1299
tri 1604 1294 1617 1307 ne
rect 1617 1301 1626 1307
tri 1626 1301 1632 1307 sw
rect 1490 1275 1535 1285
rect 1366 1247 1440 1271
rect 1308 1243 1440 1247
tri 1440 1243 1468 1271 sw
rect 1490 1261 1492 1275
tri 1490 1259 1492 1261 ne
rect 1504 1257 1535 1275
rect 1504 1247 1550 1257
rect 1617 1286 1632 1301
tri 1242 1222 1254 1234 ne
rect 1254 1229 1264 1234
tri 1264 1229 1269 1234 sw
rect 1153 883 1168 1111
rect 1254 1121 1269 1229
rect 1308 1187 1336 1243
tri 1428 1225 1446 1243 ne
rect 1446 1223 1468 1243
tri 1468 1223 1488 1243 sw
tri 1504 1229 1522 1247 ne
rect 1327 1153 1336 1187
rect 1370 1214 1412 1215
rect 1370 1180 1375 1214
rect 1405 1180 1412 1214
rect 1370 1171 1412 1180
rect 1446 1214 1488 1223
rect 1446 1180 1453 1214
rect 1483 1180 1488 1214
rect 1446 1175 1488 1180
rect 1522 1187 1550 1247
tri 1595 1234 1617 1256 se
rect 1617 1249 1632 1257
tri 1617 1234 1632 1249 nw
tri 1589 1228 1595 1234 se
rect 1595 1228 1604 1234
rect 1308 1143 1336 1153
tri 1336 1143 1360 1167 sw
rect 1254 1073 1270 1121
rect 1308 1111 1350 1143
tri 1367 1135 1368 1136 sw
rect 1367 1111 1368 1135
tri 1370 1134 1407 1171 ne
rect 1407 1143 1412 1171
tri 1412 1143 1438 1169 sw
rect 1522 1153 1531 1187
rect 1522 1143 1550 1153
rect 1407 1134 1491 1143
tri 1407 1115 1426 1134 ne
rect 1426 1115 1491 1134
rect 1308 1089 1368 1111
rect 1490 1111 1491 1115
rect 1508 1111 1550 1143
rect 1490 1089 1550 1111
rect 1396 1073 1413 1087
rect 1445 1073 1462 1087
tri 1233 1037 1255 1059 se
rect 1255 1052 1270 1073
tri 1255 1037 1270 1052 nw
rect 1589 1052 1604 1228
tri 1604 1221 1617 1234 nw
rect 1690 1153 1705 1381
tri 1227 1031 1233 1037 se
rect 1233 1031 1242 1037
rect 1227 1015 1242 1031
tri 1242 1024 1255 1037 nw
rect 1396 1029 1413 1043
rect 1445 1029 1462 1043
tri 1589 1037 1604 1052 ne
tri 1604 1037 1626 1059 sw
rect 1227 979 1242 987
rect 1308 1015 1368 1029
rect 1323 1005 1368 1015
rect 1323 987 1351 1005
tri 1227 964 1242 979 ne
tri 1242 964 1264 986 sw
rect 1308 977 1351 987
rect 1366 1001 1368 1005
rect 1490 1015 1550 1029
tri 1604 1024 1617 1037 ne
rect 1617 1031 1626 1037
tri 1626 1031 1632 1037 sw
rect 1490 1005 1535 1015
rect 1366 977 1440 1001
rect 1308 973 1440 977
tri 1440 973 1468 1001 sw
rect 1490 991 1492 1005
tri 1490 989 1492 991 ne
rect 1504 987 1535 1005
rect 1504 977 1550 987
rect 1617 1016 1632 1031
tri 1242 952 1254 964 ne
rect 1254 959 1264 964
tri 1264 959 1269 964 sw
rect 1153 613 1168 841
rect 1254 803 1269 959
rect 1308 917 1336 973
tri 1428 955 1446 973 ne
rect 1446 953 1468 973
tri 1468 953 1488 973 sw
tri 1504 959 1522 977 ne
rect 1327 883 1336 917
rect 1370 944 1412 945
rect 1370 910 1375 944
rect 1405 910 1412 944
rect 1370 901 1412 910
rect 1446 944 1488 953
rect 1446 910 1453 944
rect 1483 910 1488 944
rect 1446 905 1488 910
rect 1522 917 1550 977
tri 1595 964 1617 986 se
rect 1617 979 1632 987
tri 1617 964 1632 979 nw
tri 1589 958 1595 964 se
rect 1595 958 1604 964
rect 1308 873 1336 883
tri 1336 873 1360 897 sw
rect 1308 841 1350 873
tri 1367 865 1368 866 sw
rect 1367 841 1368 865
tri 1370 864 1407 901 ne
rect 1407 873 1412 901
tri 1412 873 1438 899 sw
rect 1522 883 1531 917
rect 1522 873 1550 883
rect 1407 864 1491 873
tri 1407 845 1426 864 ne
rect 1426 845 1491 864
rect 1308 819 1368 841
rect 1490 841 1491 845
rect 1508 841 1550 873
rect 1490 819 1550 841
rect 1396 803 1413 817
rect 1445 803 1462 817
tri 1233 767 1255 789 se
rect 1255 782 1270 803
tri 1255 767 1270 782 nw
rect 1589 782 1604 958
tri 1604 951 1617 964 nw
rect 1690 883 1705 1111
tri 1227 761 1233 767 se
rect 1233 761 1242 767
rect 1227 745 1242 761
tri 1242 754 1255 767 nw
rect 1396 759 1413 773
rect 1445 759 1462 773
tri 1589 767 1604 782 ne
tri 1604 767 1626 789 sw
rect 1227 709 1242 717
rect 1308 745 1368 759
rect 1323 735 1368 745
rect 1323 717 1351 735
tri 1227 694 1242 709 ne
tri 1242 694 1264 716 sw
rect 1308 707 1351 717
rect 1366 731 1368 735
rect 1490 745 1550 759
tri 1604 754 1617 767 ne
rect 1617 761 1626 767
tri 1626 761 1632 767 sw
rect 1490 735 1535 745
rect 1366 707 1440 731
rect 1308 703 1440 707
tri 1440 703 1468 731 sw
rect 1490 721 1492 735
tri 1490 719 1492 721 ne
rect 1504 717 1535 735
rect 1504 707 1550 717
rect 1617 746 1632 761
tri 1242 682 1254 694 ne
rect 1254 689 1264 694
tri 1264 689 1269 694 sw
rect 1153 343 1168 571
rect 1254 581 1269 689
rect 1308 647 1336 703
tri 1428 685 1446 703 ne
rect 1446 683 1468 703
tri 1468 683 1488 703 sw
tri 1504 689 1522 707 ne
rect 1327 613 1336 647
rect 1370 674 1412 675
rect 1370 640 1375 674
rect 1405 640 1412 674
rect 1370 631 1412 640
rect 1446 674 1488 683
rect 1446 640 1453 674
rect 1483 640 1488 674
rect 1446 635 1488 640
rect 1522 647 1550 707
tri 1595 694 1617 716 se
rect 1617 709 1632 717
tri 1617 694 1632 709 nw
tri 1589 688 1595 694 se
rect 1595 688 1604 694
rect 1308 603 1336 613
tri 1336 603 1360 627 sw
rect 1254 533 1270 581
rect 1308 571 1350 603
tri 1367 595 1368 596 sw
rect 1367 571 1368 595
tri 1370 594 1407 631 ne
rect 1407 603 1412 631
tri 1412 603 1438 629 sw
rect 1522 613 1531 647
rect 1522 603 1550 613
rect 1407 594 1491 603
tri 1407 575 1426 594 ne
rect 1426 575 1491 594
rect 1308 549 1368 571
rect 1490 571 1491 575
rect 1508 571 1550 603
rect 1490 549 1550 571
rect 1396 533 1413 547
rect 1445 533 1462 547
tri 1233 497 1255 519 se
rect 1255 512 1270 533
tri 1255 497 1270 512 nw
rect 1589 512 1604 688
tri 1604 681 1617 694 nw
rect 1690 613 1705 841
tri 1227 491 1233 497 se
rect 1233 491 1242 497
rect 1227 475 1242 491
tri 1242 484 1255 497 nw
rect 1396 489 1413 503
rect 1445 489 1462 503
tri 1589 497 1604 512 ne
tri 1604 497 1626 519 sw
rect 1227 439 1242 447
rect 1308 475 1368 489
rect 1323 465 1368 475
rect 1323 447 1351 465
tri 1227 424 1242 439 ne
tri 1242 424 1264 446 sw
rect 1308 437 1351 447
rect 1366 461 1368 465
rect 1490 475 1550 489
tri 1604 484 1617 497 ne
rect 1617 491 1626 497
tri 1626 491 1632 497 sw
rect 1490 465 1535 475
rect 1366 437 1440 461
rect 1308 433 1440 437
tri 1440 433 1468 461 sw
rect 1490 451 1492 465
tri 1490 449 1492 451 ne
rect 1504 447 1535 465
rect 1504 437 1550 447
rect 1617 476 1632 491
tri 1242 412 1254 424 ne
rect 1254 419 1264 424
tri 1264 419 1269 424 sw
rect 1153 73 1168 301
rect 1254 263 1269 419
rect 1308 377 1336 433
tri 1428 415 1446 433 ne
rect 1446 413 1468 433
tri 1468 413 1488 433 sw
tri 1504 419 1522 437 ne
rect 1327 343 1336 377
rect 1370 404 1412 405
rect 1370 370 1375 404
rect 1405 370 1412 404
rect 1370 361 1412 370
rect 1446 404 1488 413
rect 1446 370 1453 404
rect 1483 370 1488 404
rect 1446 365 1488 370
rect 1522 377 1550 437
tri 1595 424 1617 446 se
rect 1617 439 1632 447
tri 1617 424 1632 439 nw
tri 1589 418 1595 424 se
rect 1595 418 1604 424
rect 1308 333 1336 343
tri 1336 333 1360 357 sw
rect 1308 301 1350 333
tri 1367 325 1368 326 sw
rect 1367 301 1368 325
tri 1370 324 1407 361 ne
rect 1407 333 1412 361
tri 1412 333 1438 359 sw
rect 1522 343 1531 377
rect 1522 333 1550 343
rect 1407 324 1491 333
tri 1407 305 1426 324 ne
rect 1426 305 1491 324
rect 1308 279 1368 301
rect 1490 301 1491 305
rect 1508 301 1550 333
rect 1490 279 1550 301
rect 1396 263 1413 277
rect 1445 263 1462 277
tri 1233 227 1255 249 se
rect 1255 242 1270 263
tri 1255 227 1270 242 nw
rect 1589 242 1604 418
tri 1604 411 1617 424 nw
rect 1690 343 1705 571
tri 1227 221 1233 227 se
rect 1233 221 1242 227
rect 1227 205 1242 221
tri 1242 214 1255 227 nw
rect 1396 219 1413 233
rect 1445 219 1462 233
tri 1589 227 1604 242 ne
tri 1604 227 1626 249 sw
rect 1227 169 1242 177
rect 1308 205 1368 219
rect 1323 195 1368 205
rect 1323 177 1351 195
tri 1227 154 1242 169 ne
tri 1242 154 1264 176 sw
rect 1308 167 1351 177
rect 1366 191 1368 195
rect 1490 205 1550 219
tri 1604 214 1617 227 ne
rect 1617 221 1626 227
tri 1626 221 1632 227 sw
rect 1490 195 1535 205
rect 1366 167 1440 191
rect 1308 163 1440 167
tri 1440 163 1468 191 sw
rect 1490 181 1492 195
tri 1490 179 1492 181 ne
rect 1504 177 1535 195
rect 1504 167 1550 177
rect 1617 206 1632 221
tri 1242 142 1254 154 ne
rect 1254 149 1264 154
tri 1264 149 1269 154 sw
rect 1153 -55 1168 31
rect 1254 -55 1269 149
rect 1308 107 1336 163
tri 1428 145 1446 163 ne
rect 1446 143 1468 163
tri 1468 143 1488 163 sw
tri 1504 149 1522 167 ne
rect 1327 73 1336 107
rect 1370 134 1412 135
rect 1370 100 1375 134
rect 1405 100 1412 134
rect 1370 91 1412 100
rect 1446 134 1488 143
rect 1446 100 1453 134
rect 1483 100 1488 134
rect 1446 95 1488 100
rect 1522 107 1550 167
tri 1595 154 1617 176 se
rect 1617 169 1632 177
tri 1617 154 1632 169 nw
tri 1589 148 1595 154 se
rect 1595 148 1604 154
rect 1308 63 1336 73
tri 1336 63 1360 87 sw
rect 1308 31 1350 63
tri 1367 55 1368 56 sw
rect 1367 31 1368 55
tri 1370 54 1407 91 ne
rect 1407 63 1412 91
tri 1412 63 1438 89 sw
rect 1522 73 1531 107
rect 1522 63 1550 73
rect 1407 54 1491 63
tri 1407 35 1426 54 ne
rect 1426 35 1491 54
rect 1308 9 1368 31
rect 1490 31 1491 35
rect 1508 31 1550 63
rect 1490 9 1550 31
rect 1396 -7 1413 7
rect 1445 -7 1462 7
rect 1589 -55 1604 148
tri 1604 141 1617 154 nw
rect 1690 73 1705 301
rect 1690 -55 1705 31
rect 1733 4123 1748 4361
tri 1813 4277 1835 4299 se
rect 1835 4292 1850 4361
tri 1835 4277 1850 4292 nw
rect 2169 4292 2184 4361
tri 1807 4271 1813 4277 se
rect 1813 4271 1822 4277
rect 1807 4255 1822 4271
tri 1822 4264 1835 4277 nw
rect 1976 4269 1993 4283
rect 2025 4269 2042 4283
tri 2169 4277 2184 4292 ne
tri 2184 4277 2206 4299 sw
rect 1807 4219 1822 4227
rect 1888 4255 1948 4269
rect 1903 4245 1948 4255
rect 1903 4227 1931 4245
tri 1807 4204 1822 4219 ne
tri 1822 4204 1844 4226 sw
rect 1888 4217 1931 4227
rect 1946 4241 1948 4245
rect 2070 4255 2130 4269
tri 2184 4264 2197 4277 ne
rect 2197 4271 2206 4277
tri 2206 4271 2212 4277 sw
rect 2070 4245 2115 4255
rect 1946 4217 2020 4241
rect 1888 4213 2020 4217
tri 2020 4213 2048 4241 sw
rect 2070 4231 2072 4245
tri 2070 4229 2072 4231 ne
rect 2084 4227 2115 4245
rect 2084 4217 2130 4227
rect 2197 4256 2212 4271
tri 1822 4192 1834 4204 ne
rect 1834 4199 1844 4204
tri 1844 4199 1849 4204 sw
rect 1733 3853 1748 4081
rect 1834 4043 1849 4199
rect 1888 4157 1916 4213
tri 2008 4195 2026 4213 ne
rect 2026 4193 2048 4213
tri 2048 4193 2068 4213 sw
tri 2084 4199 2102 4217 ne
rect 1907 4123 1916 4157
rect 1950 4184 1992 4185
rect 1950 4150 1955 4184
rect 1985 4150 1992 4184
rect 1950 4141 1992 4150
rect 2026 4184 2068 4193
rect 2026 4150 2033 4184
rect 2063 4150 2068 4184
rect 2026 4145 2068 4150
rect 2102 4157 2130 4217
tri 2175 4204 2197 4226 se
rect 2197 4219 2212 4227
tri 2197 4204 2212 4219 nw
tri 2169 4198 2175 4204 se
rect 2175 4198 2184 4204
rect 1888 4113 1916 4123
tri 1916 4113 1940 4137 sw
rect 1888 4081 1930 4113
tri 1947 4105 1948 4106 sw
rect 1947 4081 1948 4105
tri 1950 4104 1987 4141 ne
rect 1987 4113 1992 4141
tri 1992 4113 2018 4139 sw
rect 2102 4123 2111 4157
rect 2102 4113 2130 4123
rect 1987 4104 2071 4113
tri 1987 4085 2006 4104 ne
rect 2006 4085 2071 4104
rect 1888 4059 1948 4081
rect 2070 4081 2071 4085
rect 2088 4081 2130 4113
rect 2070 4059 2130 4081
rect 1976 4043 1993 4057
rect 2025 4043 2042 4057
tri 1813 4007 1835 4029 se
rect 1835 4022 1850 4043
tri 1835 4007 1850 4022 nw
rect 2169 4022 2184 4198
tri 2184 4191 2197 4204 nw
rect 2270 4123 2285 4361
tri 1807 4001 1813 4007 se
rect 1813 4001 1822 4007
rect 1807 3985 1822 4001
tri 1822 3994 1835 4007 nw
rect 1976 3999 1993 4013
rect 2025 3999 2042 4013
tri 2169 4007 2184 4022 ne
tri 2184 4007 2206 4029 sw
rect 1807 3949 1822 3957
rect 1888 3985 1948 3999
rect 1903 3975 1948 3985
rect 1903 3957 1931 3975
tri 1807 3934 1822 3949 ne
tri 1822 3934 1844 3956 sw
rect 1888 3947 1931 3957
rect 1946 3971 1948 3975
rect 2070 3985 2130 3999
tri 2184 3994 2197 4007 ne
rect 2197 4001 2206 4007
tri 2206 4001 2212 4007 sw
rect 2070 3975 2115 3985
rect 1946 3947 2020 3971
rect 1888 3943 2020 3947
tri 2020 3943 2048 3971 sw
rect 2070 3961 2072 3975
tri 2070 3959 2072 3961 ne
rect 2084 3957 2115 3975
rect 2084 3947 2130 3957
rect 2197 3986 2212 4001
tri 1822 3922 1834 3934 ne
rect 1834 3929 1844 3934
tri 1844 3929 1849 3934 sw
rect 1733 3583 1748 3811
rect 1834 3821 1849 3929
rect 1888 3887 1916 3943
tri 2008 3925 2026 3943 ne
rect 2026 3923 2048 3943
tri 2048 3923 2068 3943 sw
tri 2084 3929 2102 3947 ne
rect 1907 3853 1916 3887
rect 1950 3914 1992 3915
rect 1950 3880 1955 3914
rect 1985 3880 1992 3914
rect 1950 3871 1992 3880
rect 2026 3914 2068 3923
rect 2026 3880 2033 3914
rect 2063 3880 2068 3914
rect 2026 3875 2068 3880
rect 2102 3887 2130 3947
tri 2175 3934 2197 3956 se
rect 2197 3949 2212 3957
tri 2197 3934 2212 3949 nw
tri 2169 3928 2175 3934 se
rect 2175 3928 2184 3934
rect 1888 3843 1916 3853
tri 1916 3843 1940 3867 sw
rect 1834 3773 1850 3821
rect 1888 3811 1930 3843
tri 1947 3835 1948 3836 sw
rect 1947 3811 1948 3835
tri 1950 3834 1987 3871 ne
rect 1987 3843 1992 3871
tri 1992 3843 2018 3869 sw
rect 2102 3853 2111 3887
rect 2102 3843 2130 3853
rect 1987 3834 2071 3843
tri 1987 3815 2006 3834 ne
rect 2006 3815 2071 3834
rect 1888 3789 1948 3811
rect 2070 3811 2071 3815
rect 2088 3811 2130 3843
rect 2070 3789 2130 3811
rect 1976 3773 1993 3787
rect 2025 3773 2042 3787
tri 1813 3737 1835 3759 se
rect 1835 3752 1850 3773
tri 1835 3737 1850 3752 nw
rect 2169 3752 2184 3928
tri 2184 3921 2197 3934 nw
rect 2270 3853 2285 4081
tri 1807 3731 1813 3737 se
rect 1813 3731 1822 3737
rect 1807 3715 1822 3731
tri 1822 3724 1835 3737 nw
rect 1976 3729 1993 3743
rect 2025 3729 2042 3743
tri 2169 3737 2184 3752 ne
tri 2184 3737 2206 3759 sw
rect 1807 3679 1822 3687
rect 1888 3715 1948 3729
rect 1903 3705 1948 3715
rect 1903 3687 1931 3705
tri 1807 3664 1822 3679 ne
tri 1822 3664 1844 3686 sw
rect 1888 3677 1931 3687
rect 1946 3701 1948 3705
rect 2070 3715 2130 3729
tri 2184 3724 2197 3737 ne
rect 2197 3731 2206 3737
tri 2206 3731 2212 3737 sw
rect 2070 3705 2115 3715
rect 1946 3677 2020 3701
rect 1888 3673 2020 3677
tri 2020 3673 2048 3701 sw
rect 2070 3691 2072 3705
tri 2070 3689 2072 3691 ne
rect 2084 3687 2115 3705
rect 2084 3677 2130 3687
rect 2197 3716 2212 3731
tri 1822 3652 1834 3664 ne
rect 1834 3659 1844 3664
tri 1844 3659 1849 3664 sw
rect 1733 3313 1748 3541
rect 1834 3503 1849 3659
rect 1888 3617 1916 3673
tri 2008 3655 2026 3673 ne
rect 2026 3653 2048 3673
tri 2048 3653 2068 3673 sw
tri 2084 3659 2102 3677 ne
rect 1907 3583 1916 3617
rect 1950 3644 1992 3645
rect 1950 3610 1955 3644
rect 1985 3610 1992 3644
rect 1950 3601 1992 3610
rect 2026 3644 2068 3653
rect 2026 3610 2033 3644
rect 2063 3610 2068 3644
rect 2026 3605 2068 3610
rect 2102 3617 2130 3677
tri 2175 3664 2197 3686 se
rect 2197 3679 2212 3687
tri 2197 3664 2212 3679 nw
tri 2169 3658 2175 3664 se
rect 2175 3658 2184 3664
rect 1888 3573 1916 3583
tri 1916 3573 1940 3597 sw
rect 1888 3541 1930 3573
tri 1947 3565 1948 3566 sw
rect 1947 3541 1948 3565
tri 1950 3564 1987 3601 ne
rect 1987 3573 1992 3601
tri 1992 3573 2018 3599 sw
rect 2102 3583 2111 3617
rect 2102 3573 2130 3583
rect 1987 3564 2071 3573
tri 1987 3545 2006 3564 ne
rect 2006 3545 2071 3564
rect 1888 3519 1948 3541
rect 2070 3541 2071 3545
rect 2088 3541 2130 3573
rect 2070 3519 2130 3541
rect 1976 3503 1993 3517
rect 2025 3503 2042 3517
tri 1813 3467 1835 3489 se
rect 1835 3482 1850 3503
tri 1835 3467 1850 3482 nw
rect 2169 3482 2184 3658
tri 2184 3651 2197 3664 nw
rect 2270 3583 2285 3811
tri 1807 3461 1813 3467 se
rect 1813 3461 1822 3467
rect 1807 3445 1822 3461
tri 1822 3454 1835 3467 nw
rect 1976 3459 1993 3473
rect 2025 3459 2042 3473
tri 2169 3467 2184 3482 ne
tri 2184 3467 2206 3489 sw
rect 1807 3409 1822 3417
rect 1888 3445 1948 3459
rect 1903 3435 1948 3445
rect 1903 3417 1931 3435
tri 1807 3394 1822 3409 ne
tri 1822 3394 1844 3416 sw
rect 1888 3407 1931 3417
rect 1946 3431 1948 3435
rect 2070 3445 2130 3459
tri 2184 3454 2197 3467 ne
rect 2197 3461 2206 3467
tri 2206 3461 2212 3467 sw
rect 2070 3435 2115 3445
rect 1946 3407 2020 3431
rect 1888 3403 2020 3407
tri 2020 3403 2048 3431 sw
rect 2070 3421 2072 3435
tri 2070 3419 2072 3421 ne
rect 2084 3417 2115 3435
rect 2084 3407 2130 3417
rect 2197 3446 2212 3461
tri 1822 3382 1834 3394 ne
rect 1834 3389 1844 3394
tri 1844 3389 1849 3394 sw
rect 1733 3043 1748 3271
rect 1834 3281 1849 3389
rect 1888 3347 1916 3403
tri 2008 3385 2026 3403 ne
rect 2026 3383 2048 3403
tri 2048 3383 2068 3403 sw
tri 2084 3389 2102 3407 ne
rect 1907 3313 1916 3347
rect 1950 3374 1992 3375
rect 1950 3340 1955 3374
rect 1985 3340 1992 3374
rect 1950 3331 1992 3340
rect 2026 3374 2068 3383
rect 2026 3340 2033 3374
rect 2063 3340 2068 3374
rect 2026 3335 2068 3340
rect 2102 3347 2130 3407
tri 2175 3394 2197 3416 se
rect 2197 3409 2212 3417
tri 2197 3394 2212 3409 nw
tri 2169 3388 2175 3394 se
rect 2175 3388 2184 3394
rect 1888 3303 1916 3313
tri 1916 3303 1940 3327 sw
rect 1834 3233 1850 3281
rect 1888 3271 1930 3303
tri 1947 3295 1948 3296 sw
rect 1947 3271 1948 3295
tri 1950 3294 1987 3331 ne
rect 1987 3303 1992 3331
tri 1992 3303 2018 3329 sw
rect 2102 3313 2111 3347
rect 2102 3303 2130 3313
rect 1987 3294 2071 3303
tri 1987 3275 2006 3294 ne
rect 2006 3275 2071 3294
rect 1888 3249 1948 3271
rect 2070 3271 2071 3275
rect 2088 3271 2130 3303
rect 2070 3249 2130 3271
rect 1976 3233 1993 3247
rect 2025 3233 2042 3247
tri 1813 3197 1835 3219 se
rect 1835 3212 1850 3233
tri 1835 3197 1850 3212 nw
rect 2169 3212 2184 3388
tri 2184 3381 2197 3394 nw
rect 2270 3313 2285 3541
tri 1807 3191 1813 3197 se
rect 1813 3191 1822 3197
rect 1807 3175 1822 3191
tri 1822 3184 1835 3197 nw
rect 1976 3189 1993 3203
rect 2025 3189 2042 3203
tri 2169 3197 2184 3212 ne
tri 2184 3197 2206 3219 sw
rect 1807 3139 1822 3147
rect 1888 3175 1948 3189
rect 1903 3165 1948 3175
rect 1903 3147 1931 3165
tri 1807 3124 1822 3139 ne
tri 1822 3124 1844 3146 sw
rect 1888 3137 1931 3147
rect 1946 3161 1948 3165
rect 2070 3175 2130 3189
tri 2184 3184 2197 3197 ne
rect 2197 3191 2206 3197
tri 2206 3191 2212 3197 sw
rect 2070 3165 2115 3175
rect 1946 3137 2020 3161
rect 1888 3133 2020 3137
tri 2020 3133 2048 3161 sw
rect 2070 3151 2072 3165
tri 2070 3149 2072 3151 ne
rect 2084 3147 2115 3165
rect 2084 3137 2130 3147
rect 2197 3176 2212 3191
tri 1822 3112 1834 3124 ne
rect 1834 3119 1844 3124
tri 1844 3119 1849 3124 sw
rect 1733 2773 1748 3001
rect 1834 2963 1849 3119
rect 1888 3077 1916 3133
tri 2008 3115 2026 3133 ne
rect 2026 3113 2048 3133
tri 2048 3113 2068 3133 sw
tri 2084 3119 2102 3137 ne
rect 1907 3043 1916 3077
rect 1950 3104 1992 3105
rect 1950 3070 1955 3104
rect 1985 3070 1992 3104
rect 1950 3061 1992 3070
rect 2026 3104 2068 3113
rect 2026 3070 2033 3104
rect 2063 3070 2068 3104
rect 2026 3065 2068 3070
rect 2102 3077 2130 3137
tri 2175 3124 2197 3146 se
rect 2197 3139 2212 3147
tri 2197 3124 2212 3139 nw
tri 2169 3118 2175 3124 se
rect 2175 3118 2184 3124
rect 1888 3033 1916 3043
tri 1916 3033 1940 3057 sw
rect 1888 3001 1930 3033
tri 1947 3025 1948 3026 sw
rect 1947 3001 1948 3025
tri 1950 3024 1987 3061 ne
rect 1987 3033 1992 3061
tri 1992 3033 2018 3059 sw
rect 2102 3043 2111 3077
rect 2102 3033 2130 3043
rect 1987 3024 2071 3033
tri 1987 3005 2006 3024 ne
rect 2006 3005 2071 3024
rect 1888 2979 1948 3001
rect 2070 3001 2071 3005
rect 2088 3001 2130 3033
rect 2070 2979 2130 3001
rect 1976 2963 1993 2977
rect 2025 2963 2042 2977
tri 1813 2927 1835 2949 se
rect 1835 2942 1850 2963
tri 1835 2927 1850 2942 nw
rect 2169 2942 2184 3118
tri 2184 3111 2197 3124 nw
rect 2270 3043 2285 3271
tri 1807 2921 1813 2927 se
rect 1813 2921 1822 2927
rect 1807 2905 1822 2921
tri 1822 2914 1835 2927 nw
rect 1976 2919 1993 2933
rect 2025 2919 2042 2933
tri 2169 2927 2184 2942 ne
tri 2184 2927 2206 2949 sw
rect 1807 2869 1822 2877
rect 1888 2905 1948 2919
rect 1903 2895 1948 2905
rect 1903 2877 1931 2895
tri 1807 2854 1822 2869 ne
tri 1822 2854 1844 2876 sw
rect 1888 2867 1931 2877
rect 1946 2891 1948 2895
rect 2070 2905 2130 2919
tri 2184 2914 2197 2927 ne
rect 2197 2921 2206 2927
tri 2206 2921 2212 2927 sw
rect 2070 2895 2115 2905
rect 1946 2867 2020 2891
rect 1888 2863 2020 2867
tri 2020 2863 2048 2891 sw
rect 2070 2881 2072 2895
tri 2070 2879 2072 2881 ne
rect 2084 2877 2115 2895
rect 2084 2867 2130 2877
rect 2197 2906 2212 2921
tri 1822 2842 1834 2854 ne
rect 1834 2849 1844 2854
tri 1844 2849 1849 2854 sw
rect 1733 2503 1748 2731
rect 1834 2741 1849 2849
rect 1888 2807 1916 2863
tri 2008 2845 2026 2863 ne
rect 2026 2843 2048 2863
tri 2048 2843 2068 2863 sw
tri 2084 2849 2102 2867 ne
rect 1907 2773 1916 2807
rect 1950 2834 1992 2835
rect 1950 2800 1955 2834
rect 1985 2800 1992 2834
rect 1950 2791 1992 2800
rect 2026 2834 2068 2843
rect 2026 2800 2033 2834
rect 2063 2800 2068 2834
rect 2026 2795 2068 2800
rect 2102 2807 2130 2867
tri 2175 2854 2197 2876 se
rect 2197 2869 2212 2877
tri 2197 2854 2212 2869 nw
tri 2169 2848 2175 2854 se
rect 2175 2848 2184 2854
rect 1888 2763 1916 2773
tri 1916 2763 1940 2787 sw
rect 1834 2693 1850 2741
rect 1888 2731 1930 2763
tri 1947 2755 1948 2756 sw
rect 1947 2731 1948 2755
tri 1950 2754 1987 2791 ne
rect 1987 2763 1992 2791
tri 1992 2763 2018 2789 sw
rect 2102 2773 2111 2807
rect 2102 2763 2130 2773
rect 1987 2754 2071 2763
tri 1987 2735 2006 2754 ne
rect 2006 2735 2071 2754
rect 1888 2709 1948 2731
rect 2070 2731 2071 2735
rect 2088 2731 2130 2763
rect 2070 2709 2130 2731
rect 1976 2693 1993 2707
rect 2025 2693 2042 2707
tri 1813 2657 1835 2679 se
rect 1835 2672 1850 2693
tri 1835 2657 1850 2672 nw
rect 2169 2672 2184 2848
tri 2184 2841 2197 2854 nw
rect 2270 2773 2285 3001
tri 1807 2651 1813 2657 se
rect 1813 2651 1822 2657
rect 1807 2635 1822 2651
tri 1822 2644 1835 2657 nw
rect 1976 2649 1993 2663
rect 2025 2649 2042 2663
tri 2169 2657 2184 2672 ne
tri 2184 2657 2206 2679 sw
rect 1807 2599 1822 2607
rect 1888 2635 1948 2649
rect 1903 2625 1948 2635
rect 1903 2607 1931 2625
tri 1807 2584 1822 2599 ne
tri 1822 2584 1844 2606 sw
rect 1888 2597 1931 2607
rect 1946 2621 1948 2625
rect 2070 2635 2130 2649
tri 2184 2644 2197 2657 ne
rect 2197 2651 2206 2657
tri 2206 2651 2212 2657 sw
rect 2070 2625 2115 2635
rect 1946 2597 2020 2621
rect 1888 2593 2020 2597
tri 2020 2593 2048 2621 sw
rect 2070 2611 2072 2625
tri 2070 2609 2072 2611 ne
rect 2084 2607 2115 2625
rect 2084 2597 2130 2607
rect 2197 2636 2212 2651
tri 1822 2572 1834 2584 ne
rect 1834 2579 1844 2584
tri 1844 2579 1849 2584 sw
rect 1733 2233 1748 2461
rect 1834 2423 1849 2579
rect 1888 2537 1916 2593
tri 2008 2575 2026 2593 ne
rect 2026 2573 2048 2593
tri 2048 2573 2068 2593 sw
tri 2084 2579 2102 2597 ne
rect 1907 2503 1916 2537
rect 1950 2564 1992 2565
rect 1950 2530 1955 2564
rect 1985 2530 1992 2564
rect 1950 2521 1992 2530
rect 2026 2564 2068 2573
rect 2026 2530 2033 2564
rect 2063 2530 2068 2564
rect 2026 2525 2068 2530
rect 2102 2537 2130 2597
tri 2175 2584 2197 2606 se
rect 2197 2599 2212 2607
tri 2197 2584 2212 2599 nw
tri 2169 2578 2175 2584 se
rect 2175 2578 2184 2584
rect 1888 2493 1916 2503
tri 1916 2493 1940 2517 sw
rect 1888 2461 1930 2493
tri 1947 2485 1948 2486 sw
rect 1947 2461 1948 2485
tri 1950 2484 1987 2521 ne
rect 1987 2493 1992 2521
tri 1992 2493 2018 2519 sw
rect 2102 2503 2111 2537
rect 2102 2493 2130 2503
rect 1987 2484 2071 2493
tri 1987 2465 2006 2484 ne
rect 2006 2465 2071 2484
rect 1888 2439 1948 2461
rect 2070 2461 2071 2465
rect 2088 2461 2130 2493
rect 2070 2439 2130 2461
rect 1976 2423 1993 2437
rect 2025 2423 2042 2437
tri 1813 2387 1835 2409 se
rect 1835 2402 1850 2423
tri 1835 2387 1850 2402 nw
rect 2169 2402 2184 2578
tri 2184 2571 2197 2584 nw
rect 2270 2503 2285 2731
tri 1807 2381 1813 2387 se
rect 1813 2381 1822 2387
rect 1807 2365 1822 2381
tri 1822 2374 1835 2387 nw
rect 1976 2379 1993 2393
rect 2025 2379 2042 2393
tri 2169 2387 2184 2402 ne
tri 2184 2387 2206 2409 sw
rect 1807 2329 1822 2337
rect 1888 2365 1948 2379
rect 1903 2355 1948 2365
rect 1903 2337 1931 2355
tri 1807 2314 1822 2329 ne
tri 1822 2314 1844 2336 sw
rect 1888 2327 1931 2337
rect 1946 2351 1948 2355
rect 2070 2365 2130 2379
tri 2184 2374 2197 2387 ne
rect 2197 2381 2206 2387
tri 2206 2381 2212 2387 sw
rect 2070 2355 2115 2365
rect 1946 2327 2020 2351
rect 1888 2323 2020 2327
tri 2020 2323 2048 2351 sw
rect 2070 2341 2072 2355
tri 2070 2339 2072 2341 ne
rect 2084 2337 2115 2355
rect 2084 2327 2130 2337
rect 2197 2366 2212 2381
tri 1822 2302 1834 2314 ne
rect 1834 2309 1844 2314
tri 1844 2309 1849 2314 sw
rect 1733 1963 1748 2191
rect 1834 2201 1849 2309
rect 1888 2267 1916 2323
tri 2008 2305 2026 2323 ne
rect 2026 2303 2048 2323
tri 2048 2303 2068 2323 sw
tri 2084 2309 2102 2327 ne
rect 1907 2233 1916 2267
rect 1950 2294 1992 2295
rect 1950 2260 1955 2294
rect 1985 2260 1992 2294
rect 1950 2251 1992 2260
rect 2026 2294 2068 2303
rect 2026 2260 2033 2294
rect 2063 2260 2068 2294
rect 2026 2255 2068 2260
rect 2102 2267 2130 2327
tri 2175 2314 2197 2336 se
rect 2197 2329 2212 2337
tri 2197 2314 2212 2329 nw
tri 2169 2308 2175 2314 se
rect 2175 2308 2184 2314
rect 1888 2223 1916 2233
tri 1916 2223 1940 2247 sw
rect 1834 2153 1850 2201
rect 1888 2191 1930 2223
tri 1947 2215 1948 2216 sw
rect 1947 2191 1948 2215
tri 1950 2214 1987 2251 ne
rect 1987 2223 1992 2251
tri 1992 2223 2018 2249 sw
rect 2102 2233 2111 2267
rect 2102 2223 2130 2233
rect 1987 2214 2071 2223
tri 1987 2195 2006 2214 ne
rect 2006 2195 2071 2214
rect 1888 2169 1948 2191
rect 2070 2191 2071 2195
rect 2088 2191 2130 2223
rect 2070 2169 2130 2191
rect 1976 2153 1993 2167
rect 2025 2153 2042 2167
tri 1813 2117 1835 2139 se
rect 1835 2132 1850 2153
tri 1835 2117 1850 2132 nw
rect 2169 2132 2184 2308
tri 2184 2301 2197 2314 nw
rect 2270 2233 2285 2461
tri 1807 2111 1813 2117 se
rect 1813 2111 1822 2117
rect 1807 2095 1822 2111
tri 1822 2104 1835 2117 nw
rect 1976 2109 1993 2123
rect 2025 2109 2042 2123
tri 2169 2117 2184 2132 ne
tri 2184 2117 2206 2139 sw
rect 1807 2059 1822 2067
rect 1888 2095 1948 2109
rect 1903 2085 1948 2095
rect 1903 2067 1931 2085
tri 1807 2044 1822 2059 ne
tri 1822 2044 1844 2066 sw
rect 1888 2057 1931 2067
rect 1946 2081 1948 2085
rect 2070 2095 2130 2109
tri 2184 2104 2197 2117 ne
rect 2197 2111 2206 2117
tri 2206 2111 2212 2117 sw
rect 2070 2085 2115 2095
rect 1946 2057 2020 2081
rect 1888 2053 2020 2057
tri 2020 2053 2048 2081 sw
rect 2070 2071 2072 2085
tri 2070 2069 2072 2071 ne
rect 2084 2067 2115 2085
rect 2084 2057 2130 2067
rect 2197 2096 2212 2111
tri 1822 2032 1834 2044 ne
rect 1834 2039 1844 2044
tri 1844 2039 1849 2044 sw
rect 1733 1693 1748 1921
rect 1834 1883 1849 2039
rect 1888 1997 1916 2053
tri 2008 2035 2026 2053 ne
rect 2026 2033 2048 2053
tri 2048 2033 2068 2053 sw
tri 2084 2039 2102 2057 ne
rect 1907 1963 1916 1997
rect 1950 2024 1992 2025
rect 1950 1990 1955 2024
rect 1985 1990 1992 2024
rect 1950 1981 1992 1990
rect 2026 2024 2068 2033
rect 2026 1990 2033 2024
rect 2063 1990 2068 2024
rect 2026 1985 2068 1990
rect 2102 1997 2130 2057
tri 2175 2044 2197 2066 se
rect 2197 2059 2212 2067
tri 2197 2044 2212 2059 nw
tri 2169 2038 2175 2044 se
rect 2175 2038 2184 2044
rect 1888 1953 1916 1963
tri 1916 1953 1940 1977 sw
rect 1888 1921 1930 1953
tri 1947 1945 1948 1946 sw
rect 1947 1921 1948 1945
tri 1950 1944 1987 1981 ne
rect 1987 1953 1992 1981
tri 1992 1953 2018 1979 sw
rect 2102 1963 2111 1997
rect 2102 1953 2130 1963
rect 1987 1944 2071 1953
tri 1987 1925 2006 1944 ne
rect 2006 1925 2071 1944
rect 1888 1899 1948 1921
rect 2070 1921 2071 1925
rect 2088 1921 2130 1953
rect 2070 1899 2130 1921
rect 1976 1883 1993 1897
rect 2025 1883 2042 1897
tri 1813 1847 1835 1869 se
rect 1835 1862 1850 1883
tri 1835 1847 1850 1862 nw
rect 2169 1862 2184 2038
tri 2184 2031 2197 2044 nw
rect 2270 1963 2285 2191
tri 1807 1841 1813 1847 se
rect 1813 1841 1822 1847
rect 1807 1825 1822 1841
tri 1822 1834 1835 1847 nw
rect 1976 1839 1993 1853
rect 2025 1839 2042 1853
tri 2169 1847 2184 1862 ne
tri 2184 1847 2206 1869 sw
rect 1807 1789 1822 1797
rect 1888 1825 1948 1839
rect 1903 1815 1948 1825
rect 1903 1797 1931 1815
tri 1807 1774 1822 1789 ne
tri 1822 1774 1844 1796 sw
rect 1888 1787 1931 1797
rect 1946 1811 1948 1815
rect 2070 1825 2130 1839
tri 2184 1834 2197 1847 ne
rect 2197 1841 2206 1847
tri 2206 1841 2212 1847 sw
rect 2070 1815 2115 1825
rect 1946 1787 2020 1811
rect 1888 1783 2020 1787
tri 2020 1783 2048 1811 sw
rect 2070 1801 2072 1815
tri 2070 1799 2072 1801 ne
rect 2084 1797 2115 1815
rect 2084 1787 2130 1797
rect 2197 1826 2212 1841
tri 1822 1762 1834 1774 ne
rect 1834 1769 1844 1774
tri 1844 1769 1849 1774 sw
rect 1733 1423 1748 1651
rect 1834 1661 1849 1769
rect 1888 1727 1916 1783
tri 2008 1765 2026 1783 ne
rect 2026 1763 2048 1783
tri 2048 1763 2068 1783 sw
tri 2084 1769 2102 1787 ne
rect 1907 1693 1916 1727
rect 1950 1754 1992 1755
rect 1950 1720 1955 1754
rect 1985 1720 1992 1754
rect 1950 1711 1992 1720
rect 2026 1754 2068 1763
rect 2026 1720 2033 1754
rect 2063 1720 2068 1754
rect 2026 1715 2068 1720
rect 2102 1727 2130 1787
tri 2175 1774 2197 1796 se
rect 2197 1789 2212 1797
tri 2197 1774 2212 1789 nw
tri 2169 1768 2175 1774 se
rect 2175 1768 2184 1774
rect 1888 1683 1916 1693
tri 1916 1683 1940 1707 sw
rect 1834 1613 1850 1661
rect 1888 1651 1930 1683
tri 1947 1675 1948 1676 sw
rect 1947 1651 1948 1675
tri 1950 1674 1987 1711 ne
rect 1987 1683 1992 1711
tri 1992 1683 2018 1709 sw
rect 2102 1693 2111 1727
rect 2102 1683 2130 1693
rect 1987 1674 2071 1683
tri 1987 1655 2006 1674 ne
rect 2006 1655 2071 1674
rect 1888 1629 1948 1651
rect 2070 1651 2071 1655
rect 2088 1651 2130 1683
rect 2070 1629 2130 1651
rect 1976 1613 1993 1627
rect 2025 1613 2042 1627
tri 1813 1577 1835 1599 se
rect 1835 1592 1850 1613
tri 1835 1577 1850 1592 nw
rect 2169 1592 2184 1768
tri 2184 1761 2197 1774 nw
rect 2270 1693 2285 1921
tri 1807 1571 1813 1577 se
rect 1813 1571 1822 1577
rect 1807 1555 1822 1571
tri 1822 1564 1835 1577 nw
rect 1976 1569 1993 1583
rect 2025 1569 2042 1583
tri 2169 1577 2184 1592 ne
tri 2184 1577 2206 1599 sw
rect 1807 1519 1822 1527
rect 1888 1555 1948 1569
rect 1903 1545 1948 1555
rect 1903 1527 1931 1545
tri 1807 1504 1822 1519 ne
tri 1822 1504 1844 1526 sw
rect 1888 1517 1931 1527
rect 1946 1541 1948 1545
rect 2070 1555 2130 1569
tri 2184 1564 2197 1577 ne
rect 2197 1571 2206 1577
tri 2206 1571 2212 1577 sw
rect 2070 1545 2115 1555
rect 1946 1517 2020 1541
rect 1888 1513 2020 1517
tri 2020 1513 2048 1541 sw
rect 2070 1531 2072 1545
tri 2070 1529 2072 1531 ne
rect 2084 1527 2115 1545
rect 2084 1517 2130 1527
rect 2197 1556 2212 1571
tri 1822 1492 1834 1504 ne
rect 1834 1499 1844 1504
tri 1844 1499 1849 1504 sw
rect 1733 1153 1748 1381
rect 1834 1343 1849 1499
rect 1888 1457 1916 1513
tri 2008 1495 2026 1513 ne
rect 2026 1493 2048 1513
tri 2048 1493 2068 1513 sw
tri 2084 1499 2102 1517 ne
rect 1907 1423 1916 1457
rect 1950 1484 1992 1485
rect 1950 1450 1955 1484
rect 1985 1450 1992 1484
rect 1950 1441 1992 1450
rect 2026 1484 2068 1493
rect 2026 1450 2033 1484
rect 2063 1450 2068 1484
rect 2026 1445 2068 1450
rect 2102 1457 2130 1517
tri 2175 1504 2197 1526 se
rect 2197 1519 2212 1527
tri 2197 1504 2212 1519 nw
tri 2169 1498 2175 1504 se
rect 2175 1498 2184 1504
rect 1888 1413 1916 1423
tri 1916 1413 1940 1437 sw
rect 1888 1381 1930 1413
tri 1947 1405 1948 1406 sw
rect 1947 1381 1948 1405
tri 1950 1404 1987 1441 ne
rect 1987 1413 1992 1441
tri 1992 1413 2018 1439 sw
rect 2102 1423 2111 1457
rect 2102 1413 2130 1423
rect 1987 1404 2071 1413
tri 1987 1385 2006 1404 ne
rect 2006 1385 2071 1404
rect 1888 1359 1948 1381
rect 2070 1381 2071 1385
rect 2088 1381 2130 1413
rect 2070 1359 2130 1381
rect 1976 1343 1993 1357
rect 2025 1343 2042 1357
tri 1813 1307 1835 1329 se
rect 1835 1322 1850 1343
tri 1835 1307 1850 1322 nw
rect 2169 1322 2184 1498
tri 2184 1491 2197 1504 nw
rect 2270 1423 2285 1651
tri 1807 1301 1813 1307 se
rect 1813 1301 1822 1307
rect 1807 1285 1822 1301
tri 1822 1294 1835 1307 nw
rect 1976 1299 1993 1313
rect 2025 1299 2042 1313
tri 2169 1307 2184 1322 ne
tri 2184 1307 2206 1329 sw
rect 1807 1249 1822 1257
rect 1888 1285 1948 1299
rect 1903 1275 1948 1285
rect 1903 1257 1931 1275
tri 1807 1234 1822 1249 ne
tri 1822 1234 1844 1256 sw
rect 1888 1247 1931 1257
rect 1946 1271 1948 1275
rect 2070 1285 2130 1299
tri 2184 1294 2197 1307 ne
rect 2197 1301 2206 1307
tri 2206 1301 2212 1307 sw
rect 2070 1275 2115 1285
rect 1946 1247 2020 1271
rect 1888 1243 2020 1247
tri 2020 1243 2048 1271 sw
rect 2070 1261 2072 1275
tri 2070 1259 2072 1261 ne
rect 2084 1257 2115 1275
rect 2084 1247 2130 1257
rect 2197 1286 2212 1301
tri 1822 1222 1834 1234 ne
rect 1834 1229 1844 1234
tri 1844 1229 1849 1234 sw
rect 1733 883 1748 1111
rect 1834 1121 1849 1229
rect 1888 1187 1916 1243
tri 2008 1225 2026 1243 ne
rect 2026 1223 2048 1243
tri 2048 1223 2068 1243 sw
tri 2084 1229 2102 1247 ne
rect 1907 1153 1916 1187
rect 1950 1214 1992 1215
rect 1950 1180 1955 1214
rect 1985 1180 1992 1214
rect 1950 1171 1992 1180
rect 2026 1214 2068 1223
rect 2026 1180 2033 1214
rect 2063 1180 2068 1214
rect 2026 1175 2068 1180
rect 2102 1187 2130 1247
tri 2175 1234 2197 1256 se
rect 2197 1249 2212 1257
tri 2197 1234 2212 1249 nw
tri 2169 1228 2175 1234 se
rect 2175 1228 2184 1234
rect 1888 1143 1916 1153
tri 1916 1143 1940 1167 sw
rect 1834 1073 1850 1121
rect 1888 1111 1930 1143
tri 1947 1135 1948 1136 sw
rect 1947 1111 1948 1135
tri 1950 1134 1987 1171 ne
rect 1987 1143 1992 1171
tri 1992 1143 2018 1169 sw
rect 2102 1153 2111 1187
rect 2102 1143 2130 1153
rect 1987 1134 2071 1143
tri 1987 1115 2006 1134 ne
rect 2006 1115 2071 1134
rect 1888 1089 1948 1111
rect 2070 1111 2071 1115
rect 2088 1111 2130 1143
rect 2070 1089 2130 1111
rect 1976 1073 1993 1087
rect 2025 1073 2042 1087
tri 1813 1037 1835 1059 se
rect 1835 1052 1850 1073
tri 1835 1037 1850 1052 nw
rect 2169 1052 2184 1228
tri 2184 1221 2197 1234 nw
rect 2270 1153 2285 1381
tri 1807 1031 1813 1037 se
rect 1813 1031 1822 1037
rect 1807 1015 1822 1031
tri 1822 1024 1835 1037 nw
rect 1976 1029 1993 1043
rect 2025 1029 2042 1043
tri 2169 1037 2184 1052 ne
tri 2184 1037 2206 1059 sw
rect 1807 979 1822 987
rect 1888 1015 1948 1029
rect 1903 1005 1948 1015
rect 1903 987 1931 1005
tri 1807 964 1822 979 ne
tri 1822 964 1844 986 sw
rect 1888 977 1931 987
rect 1946 1001 1948 1005
rect 2070 1015 2130 1029
tri 2184 1024 2197 1037 ne
rect 2197 1031 2206 1037
tri 2206 1031 2212 1037 sw
rect 2070 1005 2115 1015
rect 1946 977 2020 1001
rect 1888 973 2020 977
tri 2020 973 2048 1001 sw
rect 2070 991 2072 1005
tri 2070 989 2072 991 ne
rect 2084 987 2115 1005
rect 2084 977 2130 987
rect 2197 1016 2212 1031
tri 1822 952 1834 964 ne
rect 1834 959 1844 964
tri 1844 959 1849 964 sw
rect 1733 613 1748 841
rect 1834 803 1849 959
rect 1888 917 1916 973
tri 2008 955 2026 973 ne
rect 2026 953 2048 973
tri 2048 953 2068 973 sw
tri 2084 959 2102 977 ne
rect 1907 883 1916 917
rect 1950 944 1992 945
rect 1950 910 1955 944
rect 1985 910 1992 944
rect 1950 901 1992 910
rect 2026 944 2068 953
rect 2026 910 2033 944
rect 2063 910 2068 944
rect 2026 905 2068 910
rect 2102 917 2130 977
tri 2175 964 2197 986 se
rect 2197 979 2212 987
tri 2197 964 2212 979 nw
tri 2169 958 2175 964 se
rect 2175 958 2184 964
rect 1888 873 1916 883
tri 1916 873 1940 897 sw
rect 1888 841 1930 873
tri 1947 865 1948 866 sw
rect 1947 841 1948 865
tri 1950 864 1987 901 ne
rect 1987 873 1992 901
tri 1992 873 2018 899 sw
rect 2102 883 2111 917
rect 2102 873 2130 883
rect 1987 864 2071 873
tri 1987 845 2006 864 ne
rect 2006 845 2071 864
rect 1888 819 1948 841
rect 2070 841 2071 845
rect 2088 841 2130 873
rect 2070 819 2130 841
rect 1976 803 1993 817
rect 2025 803 2042 817
tri 1813 767 1835 789 se
rect 1835 782 1850 803
tri 1835 767 1850 782 nw
rect 2169 782 2184 958
tri 2184 951 2197 964 nw
rect 2270 883 2285 1111
tri 1807 761 1813 767 se
rect 1813 761 1822 767
rect 1807 745 1822 761
tri 1822 754 1835 767 nw
rect 1976 759 1993 773
rect 2025 759 2042 773
tri 2169 767 2184 782 ne
tri 2184 767 2206 789 sw
rect 1807 709 1822 717
rect 1888 745 1948 759
rect 1903 735 1948 745
rect 1903 717 1931 735
tri 1807 694 1822 709 ne
tri 1822 694 1844 716 sw
rect 1888 707 1931 717
rect 1946 731 1948 735
rect 2070 745 2130 759
tri 2184 754 2197 767 ne
rect 2197 761 2206 767
tri 2206 761 2212 767 sw
rect 2070 735 2115 745
rect 1946 707 2020 731
rect 1888 703 2020 707
tri 2020 703 2048 731 sw
rect 2070 721 2072 735
tri 2070 719 2072 721 ne
rect 2084 717 2115 735
rect 2084 707 2130 717
rect 2197 746 2212 761
tri 1822 682 1834 694 ne
rect 1834 689 1844 694
tri 1844 689 1849 694 sw
rect 1733 343 1748 571
rect 1834 581 1849 689
rect 1888 647 1916 703
tri 2008 685 2026 703 ne
rect 2026 683 2048 703
tri 2048 683 2068 703 sw
tri 2084 689 2102 707 ne
rect 1907 613 1916 647
rect 1950 674 1992 675
rect 1950 640 1955 674
rect 1985 640 1992 674
rect 1950 631 1992 640
rect 2026 674 2068 683
rect 2026 640 2033 674
rect 2063 640 2068 674
rect 2026 635 2068 640
rect 2102 647 2130 707
tri 2175 694 2197 716 se
rect 2197 709 2212 717
tri 2197 694 2212 709 nw
tri 2169 688 2175 694 se
rect 2175 688 2184 694
rect 1888 603 1916 613
tri 1916 603 1940 627 sw
rect 1834 533 1850 581
rect 1888 571 1930 603
tri 1947 595 1948 596 sw
rect 1947 571 1948 595
tri 1950 594 1987 631 ne
rect 1987 603 1992 631
tri 1992 603 2018 629 sw
rect 2102 613 2111 647
rect 2102 603 2130 613
rect 1987 594 2071 603
tri 1987 575 2006 594 ne
rect 2006 575 2071 594
rect 1888 549 1948 571
rect 2070 571 2071 575
rect 2088 571 2130 603
rect 2070 549 2130 571
rect 1976 533 1993 547
rect 2025 533 2042 547
tri 1813 497 1835 519 se
rect 1835 512 1850 533
tri 1835 497 1850 512 nw
rect 2169 512 2184 688
tri 2184 681 2197 694 nw
rect 2270 613 2285 841
tri 1807 491 1813 497 se
rect 1813 491 1822 497
rect 1807 475 1822 491
tri 1822 484 1835 497 nw
rect 1976 489 1993 503
rect 2025 489 2042 503
tri 2169 497 2184 512 ne
tri 2184 497 2206 519 sw
rect 1807 439 1822 447
rect 1888 475 1948 489
rect 1903 465 1948 475
rect 1903 447 1931 465
tri 1807 424 1822 439 ne
tri 1822 424 1844 446 sw
rect 1888 437 1931 447
rect 1946 461 1948 465
rect 2070 475 2130 489
tri 2184 484 2197 497 ne
rect 2197 491 2206 497
tri 2206 491 2212 497 sw
rect 2070 465 2115 475
rect 1946 437 2020 461
rect 1888 433 2020 437
tri 2020 433 2048 461 sw
rect 2070 451 2072 465
tri 2070 449 2072 451 ne
rect 2084 447 2115 465
rect 2084 437 2130 447
rect 2197 476 2212 491
tri 1822 412 1834 424 ne
rect 1834 419 1844 424
tri 1844 419 1849 424 sw
rect 1733 73 1748 301
rect 1834 263 1849 419
rect 1888 377 1916 433
tri 2008 415 2026 433 ne
rect 2026 413 2048 433
tri 2048 413 2068 433 sw
tri 2084 419 2102 437 ne
rect 1907 343 1916 377
rect 1950 404 1992 405
rect 1950 370 1955 404
rect 1985 370 1992 404
rect 1950 361 1992 370
rect 2026 404 2068 413
rect 2026 370 2033 404
rect 2063 370 2068 404
rect 2026 365 2068 370
rect 2102 377 2130 437
tri 2175 424 2197 446 se
rect 2197 439 2212 447
tri 2197 424 2212 439 nw
tri 2169 418 2175 424 se
rect 2175 418 2184 424
rect 1888 333 1916 343
tri 1916 333 1940 357 sw
rect 1888 301 1930 333
tri 1947 325 1948 326 sw
rect 1947 301 1948 325
tri 1950 324 1987 361 ne
rect 1987 333 1992 361
tri 1992 333 2018 359 sw
rect 2102 343 2111 377
rect 2102 333 2130 343
rect 1987 324 2071 333
tri 1987 305 2006 324 ne
rect 2006 305 2071 324
rect 1888 279 1948 301
rect 2070 301 2071 305
rect 2088 301 2130 333
rect 2070 279 2130 301
rect 1976 263 1993 277
rect 2025 263 2042 277
tri 1813 227 1835 249 se
rect 1835 242 1850 263
tri 1835 227 1850 242 nw
rect 2169 242 2184 418
tri 2184 411 2197 424 nw
rect 2270 343 2285 571
tri 1807 221 1813 227 se
rect 1813 221 1822 227
rect 1807 205 1822 221
tri 1822 214 1835 227 nw
rect 1976 219 1993 233
rect 2025 219 2042 233
tri 2169 227 2184 242 ne
tri 2184 227 2206 249 sw
rect 1807 169 1822 177
rect 1888 205 1948 219
rect 1903 195 1948 205
rect 1903 177 1931 195
tri 1807 154 1822 169 ne
tri 1822 154 1844 176 sw
rect 1888 167 1931 177
rect 1946 191 1948 195
rect 2070 205 2130 219
tri 2184 214 2197 227 ne
rect 2197 221 2206 227
tri 2206 221 2212 227 sw
rect 2070 195 2115 205
rect 1946 167 2020 191
rect 1888 163 2020 167
tri 2020 163 2048 191 sw
rect 2070 181 2072 195
tri 2070 179 2072 181 ne
rect 2084 177 2115 195
rect 2084 167 2130 177
rect 2197 206 2212 221
tri 1822 142 1834 154 ne
rect 1834 149 1844 154
tri 1844 149 1849 154 sw
rect 1733 -55 1748 31
rect 1834 -55 1849 149
rect 1888 107 1916 163
tri 2008 145 2026 163 ne
rect 2026 143 2048 163
tri 2048 143 2068 163 sw
tri 2084 149 2102 167 ne
rect 1907 73 1916 107
rect 1950 134 1992 135
rect 1950 100 1955 134
rect 1985 100 1992 134
rect 1950 91 1992 100
rect 2026 134 2068 143
rect 2026 100 2033 134
rect 2063 100 2068 134
rect 2026 95 2068 100
rect 2102 107 2130 167
tri 2175 154 2197 176 se
rect 2197 169 2212 177
tri 2197 154 2212 169 nw
tri 2169 148 2175 154 se
rect 2175 148 2184 154
rect 1888 63 1916 73
tri 1916 63 1940 87 sw
rect 1888 31 1930 63
tri 1947 55 1948 56 sw
rect 1947 31 1948 55
tri 1950 54 1987 91 ne
rect 1987 63 1992 91
tri 1992 63 2018 89 sw
rect 2102 73 2111 107
rect 2102 63 2130 73
rect 1987 54 2071 63
tri 1987 35 2006 54 ne
rect 2006 35 2071 54
rect 1888 9 1948 31
rect 2070 31 2071 35
rect 2088 31 2130 63
rect 2070 9 2130 31
rect 1976 -7 1993 7
rect 2025 -7 2042 7
rect 2169 -55 2184 148
tri 2184 141 2197 154 nw
rect 2270 73 2285 301
rect 2270 -55 2285 31
rect 2313 4123 2328 4361
tri 2393 4277 2415 4299 se
rect 2415 4292 2430 4361
tri 2415 4277 2430 4292 nw
rect 2749 4292 2764 4361
tri 2387 4271 2393 4277 se
rect 2393 4271 2402 4277
rect 2387 4255 2402 4271
tri 2402 4264 2415 4277 nw
rect 2556 4269 2573 4283
rect 2605 4269 2622 4283
tri 2749 4277 2764 4292 ne
tri 2764 4277 2786 4299 sw
rect 2387 4219 2402 4227
rect 2468 4255 2528 4269
rect 2483 4245 2528 4255
rect 2483 4227 2511 4245
tri 2387 4204 2402 4219 ne
tri 2402 4204 2424 4226 sw
rect 2468 4217 2511 4227
rect 2526 4241 2528 4245
rect 2650 4255 2710 4269
tri 2764 4264 2777 4277 ne
rect 2777 4271 2786 4277
tri 2786 4271 2792 4277 sw
rect 2650 4245 2695 4255
rect 2526 4217 2600 4241
rect 2468 4213 2600 4217
tri 2600 4213 2628 4241 sw
rect 2650 4231 2652 4245
tri 2650 4229 2652 4231 ne
rect 2664 4227 2695 4245
rect 2664 4217 2710 4227
rect 2777 4256 2792 4271
tri 2402 4192 2414 4204 ne
rect 2414 4199 2424 4204
tri 2424 4199 2429 4204 sw
rect 2313 3853 2328 4081
rect 2414 4043 2429 4199
rect 2468 4157 2496 4213
tri 2588 4195 2606 4213 ne
rect 2606 4193 2628 4213
tri 2628 4193 2648 4213 sw
tri 2664 4199 2682 4217 ne
rect 2487 4123 2496 4157
rect 2530 4184 2572 4185
rect 2530 4150 2535 4184
rect 2565 4150 2572 4184
rect 2530 4141 2572 4150
rect 2606 4184 2648 4193
rect 2606 4150 2613 4184
rect 2643 4150 2648 4184
rect 2606 4145 2648 4150
rect 2682 4157 2710 4217
tri 2755 4204 2777 4226 se
rect 2777 4219 2792 4227
tri 2777 4204 2792 4219 nw
tri 2749 4198 2755 4204 se
rect 2755 4198 2764 4204
rect 2468 4113 2496 4123
tri 2496 4113 2520 4137 sw
rect 2468 4081 2510 4113
tri 2527 4105 2528 4106 sw
rect 2527 4081 2528 4105
tri 2530 4104 2567 4141 ne
rect 2567 4113 2572 4141
tri 2572 4113 2598 4139 sw
rect 2682 4123 2691 4157
rect 2682 4113 2710 4123
rect 2567 4104 2651 4113
tri 2567 4085 2586 4104 ne
rect 2586 4085 2651 4104
rect 2468 4059 2528 4081
rect 2650 4081 2651 4085
rect 2668 4081 2710 4113
rect 2650 4059 2710 4081
rect 2556 4043 2573 4057
rect 2605 4043 2622 4057
tri 2393 4007 2415 4029 se
rect 2415 4022 2430 4043
tri 2415 4007 2430 4022 nw
rect 2749 4022 2764 4198
tri 2764 4191 2777 4204 nw
rect 2850 4123 2865 4361
tri 2387 4001 2393 4007 se
rect 2393 4001 2402 4007
rect 2387 3985 2402 4001
tri 2402 3994 2415 4007 nw
rect 2556 3999 2573 4013
rect 2605 3999 2622 4013
tri 2749 4007 2764 4022 ne
tri 2764 4007 2786 4029 sw
rect 2387 3949 2402 3957
rect 2468 3985 2528 3999
rect 2483 3975 2528 3985
rect 2483 3957 2511 3975
tri 2387 3934 2402 3949 ne
tri 2402 3934 2424 3956 sw
rect 2468 3947 2511 3957
rect 2526 3971 2528 3975
rect 2650 3985 2710 3999
tri 2764 3994 2777 4007 ne
rect 2777 4001 2786 4007
tri 2786 4001 2792 4007 sw
rect 2650 3975 2695 3985
rect 2526 3947 2600 3971
rect 2468 3943 2600 3947
tri 2600 3943 2628 3971 sw
rect 2650 3961 2652 3975
tri 2650 3959 2652 3961 ne
rect 2664 3957 2695 3975
rect 2664 3947 2710 3957
rect 2777 3986 2792 4001
tri 2402 3922 2414 3934 ne
rect 2414 3929 2424 3934
tri 2424 3929 2429 3934 sw
rect 2313 3583 2328 3811
rect 2414 3821 2429 3929
rect 2468 3887 2496 3943
tri 2588 3925 2606 3943 ne
rect 2606 3923 2628 3943
tri 2628 3923 2648 3943 sw
tri 2664 3929 2682 3947 ne
rect 2487 3853 2496 3887
rect 2530 3914 2572 3915
rect 2530 3880 2535 3914
rect 2565 3880 2572 3914
rect 2530 3871 2572 3880
rect 2606 3914 2648 3923
rect 2606 3880 2613 3914
rect 2643 3880 2648 3914
rect 2606 3875 2648 3880
rect 2682 3887 2710 3947
tri 2755 3934 2777 3956 se
rect 2777 3949 2792 3957
tri 2777 3934 2792 3949 nw
tri 2749 3928 2755 3934 se
rect 2755 3928 2764 3934
rect 2468 3843 2496 3853
tri 2496 3843 2520 3867 sw
rect 2414 3773 2430 3821
rect 2468 3811 2510 3843
tri 2527 3835 2528 3836 sw
rect 2527 3811 2528 3835
tri 2530 3834 2567 3871 ne
rect 2567 3843 2572 3871
tri 2572 3843 2598 3869 sw
rect 2682 3853 2691 3887
rect 2682 3843 2710 3853
rect 2567 3834 2651 3843
tri 2567 3815 2586 3834 ne
rect 2586 3815 2651 3834
rect 2468 3789 2528 3811
rect 2650 3811 2651 3815
rect 2668 3811 2710 3843
rect 2650 3789 2710 3811
rect 2556 3773 2573 3787
rect 2605 3773 2622 3787
tri 2393 3737 2415 3759 se
rect 2415 3752 2430 3773
tri 2415 3737 2430 3752 nw
rect 2749 3752 2764 3928
tri 2764 3921 2777 3934 nw
rect 2850 3853 2865 4081
tri 2387 3731 2393 3737 se
rect 2393 3731 2402 3737
rect 2387 3715 2402 3731
tri 2402 3724 2415 3737 nw
rect 2556 3729 2573 3743
rect 2605 3729 2622 3743
tri 2749 3737 2764 3752 ne
tri 2764 3737 2786 3759 sw
rect 2387 3679 2402 3687
rect 2468 3715 2528 3729
rect 2483 3705 2528 3715
rect 2483 3687 2511 3705
tri 2387 3664 2402 3679 ne
tri 2402 3664 2424 3686 sw
rect 2468 3677 2511 3687
rect 2526 3701 2528 3705
rect 2650 3715 2710 3729
tri 2764 3724 2777 3737 ne
rect 2777 3731 2786 3737
tri 2786 3731 2792 3737 sw
rect 2650 3705 2695 3715
rect 2526 3677 2600 3701
rect 2468 3673 2600 3677
tri 2600 3673 2628 3701 sw
rect 2650 3691 2652 3705
tri 2650 3689 2652 3691 ne
rect 2664 3687 2695 3705
rect 2664 3677 2710 3687
rect 2777 3716 2792 3731
tri 2402 3652 2414 3664 ne
rect 2414 3659 2424 3664
tri 2424 3659 2429 3664 sw
rect 2313 3313 2328 3541
rect 2414 3503 2429 3659
rect 2468 3617 2496 3673
tri 2588 3655 2606 3673 ne
rect 2606 3653 2628 3673
tri 2628 3653 2648 3673 sw
tri 2664 3659 2682 3677 ne
rect 2487 3583 2496 3617
rect 2530 3644 2572 3645
rect 2530 3610 2535 3644
rect 2565 3610 2572 3644
rect 2530 3601 2572 3610
rect 2606 3644 2648 3653
rect 2606 3610 2613 3644
rect 2643 3610 2648 3644
rect 2606 3605 2648 3610
rect 2682 3617 2710 3677
tri 2755 3664 2777 3686 se
rect 2777 3679 2792 3687
tri 2777 3664 2792 3679 nw
tri 2749 3658 2755 3664 se
rect 2755 3658 2764 3664
rect 2468 3573 2496 3583
tri 2496 3573 2520 3597 sw
rect 2468 3541 2510 3573
tri 2527 3565 2528 3566 sw
rect 2527 3541 2528 3565
tri 2530 3564 2567 3601 ne
rect 2567 3573 2572 3601
tri 2572 3573 2598 3599 sw
rect 2682 3583 2691 3617
rect 2682 3573 2710 3583
rect 2567 3564 2651 3573
tri 2567 3545 2586 3564 ne
rect 2586 3545 2651 3564
rect 2468 3519 2528 3541
rect 2650 3541 2651 3545
rect 2668 3541 2710 3573
rect 2650 3519 2710 3541
rect 2556 3503 2573 3517
rect 2605 3503 2622 3517
tri 2393 3467 2415 3489 se
rect 2415 3482 2430 3503
tri 2415 3467 2430 3482 nw
rect 2749 3482 2764 3658
tri 2764 3651 2777 3664 nw
rect 2850 3583 2865 3811
tri 2387 3461 2393 3467 se
rect 2393 3461 2402 3467
rect 2387 3445 2402 3461
tri 2402 3454 2415 3467 nw
rect 2556 3459 2573 3473
rect 2605 3459 2622 3473
tri 2749 3467 2764 3482 ne
tri 2764 3467 2786 3489 sw
rect 2387 3409 2402 3417
rect 2468 3445 2528 3459
rect 2483 3435 2528 3445
rect 2483 3417 2511 3435
tri 2387 3394 2402 3409 ne
tri 2402 3394 2424 3416 sw
rect 2468 3407 2511 3417
rect 2526 3431 2528 3435
rect 2650 3445 2710 3459
tri 2764 3454 2777 3467 ne
rect 2777 3461 2786 3467
tri 2786 3461 2792 3467 sw
rect 2650 3435 2695 3445
rect 2526 3407 2600 3431
rect 2468 3403 2600 3407
tri 2600 3403 2628 3431 sw
rect 2650 3421 2652 3435
tri 2650 3419 2652 3421 ne
rect 2664 3417 2695 3435
rect 2664 3407 2710 3417
rect 2777 3446 2792 3461
tri 2402 3382 2414 3394 ne
rect 2414 3389 2424 3394
tri 2424 3389 2429 3394 sw
rect 2313 3043 2328 3271
rect 2414 3281 2429 3389
rect 2468 3347 2496 3403
tri 2588 3385 2606 3403 ne
rect 2606 3383 2628 3403
tri 2628 3383 2648 3403 sw
tri 2664 3389 2682 3407 ne
rect 2487 3313 2496 3347
rect 2530 3374 2572 3375
rect 2530 3340 2535 3374
rect 2565 3340 2572 3374
rect 2530 3331 2572 3340
rect 2606 3374 2648 3383
rect 2606 3340 2613 3374
rect 2643 3340 2648 3374
rect 2606 3335 2648 3340
rect 2682 3347 2710 3407
tri 2755 3394 2777 3416 se
rect 2777 3409 2792 3417
tri 2777 3394 2792 3409 nw
tri 2749 3388 2755 3394 se
rect 2755 3388 2764 3394
rect 2468 3303 2496 3313
tri 2496 3303 2520 3327 sw
rect 2414 3233 2430 3281
rect 2468 3271 2510 3303
tri 2527 3295 2528 3296 sw
rect 2527 3271 2528 3295
tri 2530 3294 2567 3331 ne
rect 2567 3303 2572 3331
tri 2572 3303 2598 3329 sw
rect 2682 3313 2691 3347
rect 2682 3303 2710 3313
rect 2567 3294 2651 3303
tri 2567 3275 2586 3294 ne
rect 2586 3275 2651 3294
rect 2468 3249 2528 3271
rect 2650 3271 2651 3275
rect 2668 3271 2710 3303
rect 2650 3249 2710 3271
rect 2556 3233 2573 3247
rect 2605 3233 2622 3247
tri 2393 3197 2415 3219 se
rect 2415 3212 2430 3233
tri 2415 3197 2430 3212 nw
rect 2749 3212 2764 3388
tri 2764 3381 2777 3394 nw
rect 2850 3313 2865 3541
tri 2387 3191 2393 3197 se
rect 2393 3191 2402 3197
rect 2387 3175 2402 3191
tri 2402 3184 2415 3197 nw
rect 2556 3189 2573 3203
rect 2605 3189 2622 3203
tri 2749 3197 2764 3212 ne
tri 2764 3197 2786 3219 sw
rect 2387 3139 2402 3147
rect 2468 3175 2528 3189
rect 2483 3165 2528 3175
rect 2483 3147 2511 3165
tri 2387 3124 2402 3139 ne
tri 2402 3124 2424 3146 sw
rect 2468 3137 2511 3147
rect 2526 3161 2528 3165
rect 2650 3175 2710 3189
tri 2764 3184 2777 3197 ne
rect 2777 3191 2786 3197
tri 2786 3191 2792 3197 sw
rect 2650 3165 2695 3175
rect 2526 3137 2600 3161
rect 2468 3133 2600 3137
tri 2600 3133 2628 3161 sw
rect 2650 3151 2652 3165
tri 2650 3149 2652 3151 ne
rect 2664 3147 2695 3165
rect 2664 3137 2710 3147
rect 2777 3176 2792 3191
tri 2402 3112 2414 3124 ne
rect 2414 3119 2424 3124
tri 2424 3119 2429 3124 sw
rect 2313 2773 2328 3001
rect 2414 2963 2429 3119
rect 2468 3077 2496 3133
tri 2588 3115 2606 3133 ne
rect 2606 3113 2628 3133
tri 2628 3113 2648 3133 sw
tri 2664 3119 2682 3137 ne
rect 2487 3043 2496 3077
rect 2530 3104 2572 3105
rect 2530 3070 2535 3104
rect 2565 3070 2572 3104
rect 2530 3061 2572 3070
rect 2606 3104 2648 3113
rect 2606 3070 2613 3104
rect 2643 3070 2648 3104
rect 2606 3065 2648 3070
rect 2682 3077 2710 3137
tri 2755 3124 2777 3146 se
rect 2777 3139 2792 3147
tri 2777 3124 2792 3139 nw
tri 2749 3118 2755 3124 se
rect 2755 3118 2764 3124
rect 2468 3033 2496 3043
tri 2496 3033 2520 3057 sw
rect 2468 3001 2510 3033
tri 2527 3025 2528 3026 sw
rect 2527 3001 2528 3025
tri 2530 3024 2567 3061 ne
rect 2567 3033 2572 3061
tri 2572 3033 2598 3059 sw
rect 2682 3043 2691 3077
rect 2682 3033 2710 3043
rect 2567 3024 2651 3033
tri 2567 3005 2586 3024 ne
rect 2586 3005 2651 3024
rect 2468 2979 2528 3001
rect 2650 3001 2651 3005
rect 2668 3001 2710 3033
rect 2650 2979 2710 3001
rect 2556 2963 2573 2977
rect 2605 2963 2622 2977
tri 2393 2927 2415 2949 se
rect 2415 2942 2430 2963
tri 2415 2927 2430 2942 nw
rect 2749 2942 2764 3118
tri 2764 3111 2777 3124 nw
rect 2850 3043 2865 3271
tri 2387 2921 2393 2927 se
rect 2393 2921 2402 2927
rect 2387 2905 2402 2921
tri 2402 2914 2415 2927 nw
rect 2556 2919 2573 2933
rect 2605 2919 2622 2933
tri 2749 2927 2764 2942 ne
tri 2764 2927 2786 2949 sw
rect 2387 2869 2402 2877
rect 2468 2905 2528 2919
rect 2483 2895 2528 2905
rect 2483 2877 2511 2895
tri 2387 2854 2402 2869 ne
tri 2402 2854 2424 2876 sw
rect 2468 2867 2511 2877
rect 2526 2891 2528 2895
rect 2650 2905 2710 2919
tri 2764 2914 2777 2927 ne
rect 2777 2921 2786 2927
tri 2786 2921 2792 2927 sw
rect 2650 2895 2695 2905
rect 2526 2867 2600 2891
rect 2468 2863 2600 2867
tri 2600 2863 2628 2891 sw
rect 2650 2881 2652 2895
tri 2650 2879 2652 2881 ne
rect 2664 2877 2695 2895
rect 2664 2867 2710 2877
rect 2777 2906 2792 2921
tri 2402 2842 2414 2854 ne
rect 2414 2849 2424 2854
tri 2424 2849 2429 2854 sw
rect 2313 2503 2328 2731
rect 2414 2741 2429 2849
rect 2468 2807 2496 2863
tri 2588 2845 2606 2863 ne
rect 2606 2843 2628 2863
tri 2628 2843 2648 2863 sw
tri 2664 2849 2682 2867 ne
rect 2487 2773 2496 2807
rect 2530 2834 2572 2835
rect 2530 2800 2535 2834
rect 2565 2800 2572 2834
rect 2530 2791 2572 2800
rect 2606 2834 2648 2843
rect 2606 2800 2613 2834
rect 2643 2800 2648 2834
rect 2606 2795 2648 2800
rect 2682 2807 2710 2867
tri 2755 2854 2777 2876 se
rect 2777 2869 2792 2877
tri 2777 2854 2792 2869 nw
tri 2749 2848 2755 2854 se
rect 2755 2848 2764 2854
rect 2468 2763 2496 2773
tri 2496 2763 2520 2787 sw
rect 2414 2693 2430 2741
rect 2468 2731 2510 2763
tri 2527 2755 2528 2756 sw
rect 2527 2731 2528 2755
tri 2530 2754 2567 2791 ne
rect 2567 2763 2572 2791
tri 2572 2763 2598 2789 sw
rect 2682 2773 2691 2807
rect 2682 2763 2710 2773
rect 2567 2754 2651 2763
tri 2567 2735 2586 2754 ne
rect 2586 2735 2651 2754
rect 2468 2709 2528 2731
rect 2650 2731 2651 2735
rect 2668 2731 2710 2763
rect 2650 2709 2710 2731
rect 2556 2693 2573 2707
rect 2605 2693 2622 2707
tri 2393 2657 2415 2679 se
rect 2415 2672 2430 2693
tri 2415 2657 2430 2672 nw
rect 2749 2672 2764 2848
tri 2764 2841 2777 2854 nw
rect 2850 2773 2865 3001
tri 2387 2651 2393 2657 se
rect 2393 2651 2402 2657
rect 2387 2635 2402 2651
tri 2402 2644 2415 2657 nw
rect 2556 2649 2573 2663
rect 2605 2649 2622 2663
tri 2749 2657 2764 2672 ne
tri 2764 2657 2786 2679 sw
rect 2387 2599 2402 2607
rect 2468 2635 2528 2649
rect 2483 2625 2528 2635
rect 2483 2607 2511 2625
tri 2387 2584 2402 2599 ne
tri 2402 2584 2424 2606 sw
rect 2468 2597 2511 2607
rect 2526 2621 2528 2625
rect 2650 2635 2710 2649
tri 2764 2644 2777 2657 ne
rect 2777 2651 2786 2657
tri 2786 2651 2792 2657 sw
rect 2650 2625 2695 2635
rect 2526 2597 2600 2621
rect 2468 2593 2600 2597
tri 2600 2593 2628 2621 sw
rect 2650 2611 2652 2625
tri 2650 2609 2652 2611 ne
rect 2664 2607 2695 2625
rect 2664 2597 2710 2607
rect 2777 2636 2792 2651
tri 2402 2572 2414 2584 ne
rect 2414 2579 2424 2584
tri 2424 2579 2429 2584 sw
rect 2313 2233 2328 2461
rect 2414 2423 2429 2579
rect 2468 2537 2496 2593
tri 2588 2575 2606 2593 ne
rect 2606 2573 2628 2593
tri 2628 2573 2648 2593 sw
tri 2664 2579 2682 2597 ne
rect 2487 2503 2496 2537
rect 2530 2564 2572 2565
rect 2530 2530 2535 2564
rect 2565 2530 2572 2564
rect 2530 2521 2572 2530
rect 2606 2564 2648 2573
rect 2606 2530 2613 2564
rect 2643 2530 2648 2564
rect 2606 2525 2648 2530
rect 2682 2537 2710 2597
tri 2755 2584 2777 2606 se
rect 2777 2599 2792 2607
tri 2777 2584 2792 2599 nw
tri 2749 2578 2755 2584 se
rect 2755 2578 2764 2584
rect 2468 2493 2496 2503
tri 2496 2493 2520 2517 sw
rect 2468 2461 2510 2493
tri 2527 2485 2528 2486 sw
rect 2527 2461 2528 2485
tri 2530 2484 2567 2521 ne
rect 2567 2493 2572 2521
tri 2572 2493 2598 2519 sw
rect 2682 2503 2691 2537
rect 2682 2493 2710 2503
rect 2567 2484 2651 2493
tri 2567 2465 2586 2484 ne
rect 2586 2465 2651 2484
rect 2468 2439 2528 2461
rect 2650 2461 2651 2465
rect 2668 2461 2710 2493
rect 2650 2439 2710 2461
rect 2556 2423 2573 2437
rect 2605 2423 2622 2437
tri 2393 2387 2415 2409 se
rect 2415 2402 2430 2423
tri 2415 2387 2430 2402 nw
rect 2749 2402 2764 2578
tri 2764 2571 2777 2584 nw
rect 2850 2503 2865 2731
tri 2387 2381 2393 2387 se
rect 2393 2381 2402 2387
rect 2387 2365 2402 2381
tri 2402 2374 2415 2387 nw
rect 2556 2379 2573 2393
rect 2605 2379 2622 2393
tri 2749 2387 2764 2402 ne
tri 2764 2387 2786 2409 sw
rect 2387 2329 2402 2337
rect 2468 2365 2528 2379
rect 2483 2355 2528 2365
rect 2483 2337 2511 2355
tri 2387 2314 2402 2329 ne
tri 2402 2314 2424 2336 sw
rect 2468 2327 2511 2337
rect 2526 2351 2528 2355
rect 2650 2365 2710 2379
tri 2764 2374 2777 2387 ne
rect 2777 2381 2786 2387
tri 2786 2381 2792 2387 sw
rect 2650 2355 2695 2365
rect 2526 2327 2600 2351
rect 2468 2323 2600 2327
tri 2600 2323 2628 2351 sw
rect 2650 2341 2652 2355
tri 2650 2339 2652 2341 ne
rect 2664 2337 2695 2355
rect 2664 2327 2710 2337
rect 2777 2366 2792 2381
tri 2402 2302 2414 2314 ne
rect 2414 2309 2424 2314
tri 2424 2309 2429 2314 sw
rect 2313 1963 2328 2191
rect 2414 2201 2429 2309
rect 2468 2267 2496 2323
tri 2588 2305 2606 2323 ne
rect 2606 2303 2628 2323
tri 2628 2303 2648 2323 sw
tri 2664 2309 2682 2327 ne
rect 2487 2233 2496 2267
rect 2530 2294 2572 2295
rect 2530 2260 2535 2294
rect 2565 2260 2572 2294
rect 2530 2251 2572 2260
rect 2606 2294 2648 2303
rect 2606 2260 2613 2294
rect 2643 2260 2648 2294
rect 2606 2255 2648 2260
rect 2682 2267 2710 2327
tri 2755 2314 2777 2336 se
rect 2777 2329 2792 2337
tri 2777 2314 2792 2329 nw
tri 2749 2308 2755 2314 se
rect 2755 2308 2764 2314
rect 2468 2223 2496 2233
tri 2496 2223 2520 2247 sw
rect 2414 2153 2430 2201
rect 2468 2191 2510 2223
tri 2527 2215 2528 2216 sw
rect 2527 2191 2528 2215
tri 2530 2214 2567 2251 ne
rect 2567 2223 2572 2251
tri 2572 2223 2598 2249 sw
rect 2682 2233 2691 2267
rect 2682 2223 2710 2233
rect 2567 2214 2651 2223
tri 2567 2195 2586 2214 ne
rect 2586 2195 2651 2214
rect 2468 2169 2528 2191
rect 2650 2191 2651 2195
rect 2668 2191 2710 2223
rect 2650 2169 2710 2191
rect 2556 2153 2573 2167
rect 2605 2153 2622 2167
tri 2393 2117 2415 2139 se
rect 2415 2132 2430 2153
tri 2415 2117 2430 2132 nw
rect 2749 2132 2764 2308
tri 2764 2301 2777 2314 nw
rect 2850 2233 2865 2461
tri 2387 2111 2393 2117 se
rect 2393 2111 2402 2117
rect 2387 2095 2402 2111
tri 2402 2104 2415 2117 nw
rect 2556 2109 2573 2123
rect 2605 2109 2622 2123
tri 2749 2117 2764 2132 ne
tri 2764 2117 2786 2139 sw
rect 2387 2059 2402 2067
rect 2468 2095 2528 2109
rect 2483 2085 2528 2095
rect 2483 2067 2511 2085
tri 2387 2044 2402 2059 ne
tri 2402 2044 2424 2066 sw
rect 2468 2057 2511 2067
rect 2526 2081 2528 2085
rect 2650 2095 2710 2109
tri 2764 2104 2777 2117 ne
rect 2777 2111 2786 2117
tri 2786 2111 2792 2117 sw
rect 2650 2085 2695 2095
rect 2526 2057 2600 2081
rect 2468 2053 2600 2057
tri 2600 2053 2628 2081 sw
rect 2650 2071 2652 2085
tri 2650 2069 2652 2071 ne
rect 2664 2067 2695 2085
rect 2664 2057 2710 2067
rect 2777 2096 2792 2111
tri 2402 2032 2414 2044 ne
rect 2414 2039 2424 2044
tri 2424 2039 2429 2044 sw
rect 2313 1693 2328 1921
rect 2414 1883 2429 2039
rect 2468 1997 2496 2053
tri 2588 2035 2606 2053 ne
rect 2606 2033 2628 2053
tri 2628 2033 2648 2053 sw
tri 2664 2039 2682 2057 ne
rect 2487 1963 2496 1997
rect 2530 2024 2572 2025
rect 2530 1990 2535 2024
rect 2565 1990 2572 2024
rect 2530 1981 2572 1990
rect 2606 2024 2648 2033
rect 2606 1990 2613 2024
rect 2643 1990 2648 2024
rect 2606 1985 2648 1990
rect 2682 1997 2710 2057
tri 2755 2044 2777 2066 se
rect 2777 2059 2792 2067
tri 2777 2044 2792 2059 nw
tri 2749 2038 2755 2044 se
rect 2755 2038 2764 2044
rect 2468 1953 2496 1963
tri 2496 1953 2520 1977 sw
rect 2468 1921 2510 1953
tri 2527 1945 2528 1946 sw
rect 2527 1921 2528 1945
tri 2530 1944 2567 1981 ne
rect 2567 1953 2572 1981
tri 2572 1953 2598 1979 sw
rect 2682 1963 2691 1997
rect 2682 1953 2710 1963
rect 2567 1944 2651 1953
tri 2567 1925 2586 1944 ne
rect 2586 1925 2651 1944
rect 2468 1899 2528 1921
rect 2650 1921 2651 1925
rect 2668 1921 2710 1953
rect 2650 1899 2710 1921
rect 2556 1883 2573 1897
rect 2605 1883 2622 1897
tri 2393 1847 2415 1869 se
rect 2415 1862 2430 1883
tri 2415 1847 2430 1862 nw
rect 2749 1862 2764 2038
tri 2764 2031 2777 2044 nw
rect 2850 1963 2865 2191
tri 2387 1841 2393 1847 se
rect 2393 1841 2402 1847
rect 2387 1825 2402 1841
tri 2402 1834 2415 1847 nw
rect 2556 1839 2573 1853
rect 2605 1839 2622 1853
tri 2749 1847 2764 1862 ne
tri 2764 1847 2786 1869 sw
rect 2387 1789 2402 1797
rect 2468 1825 2528 1839
rect 2483 1815 2528 1825
rect 2483 1797 2511 1815
tri 2387 1774 2402 1789 ne
tri 2402 1774 2424 1796 sw
rect 2468 1787 2511 1797
rect 2526 1811 2528 1815
rect 2650 1825 2710 1839
tri 2764 1834 2777 1847 ne
rect 2777 1841 2786 1847
tri 2786 1841 2792 1847 sw
rect 2650 1815 2695 1825
rect 2526 1787 2600 1811
rect 2468 1783 2600 1787
tri 2600 1783 2628 1811 sw
rect 2650 1801 2652 1815
tri 2650 1799 2652 1801 ne
rect 2664 1797 2695 1815
rect 2664 1787 2710 1797
rect 2777 1826 2792 1841
tri 2402 1762 2414 1774 ne
rect 2414 1769 2424 1774
tri 2424 1769 2429 1774 sw
rect 2313 1423 2328 1651
rect 2414 1661 2429 1769
rect 2468 1727 2496 1783
tri 2588 1765 2606 1783 ne
rect 2606 1763 2628 1783
tri 2628 1763 2648 1783 sw
tri 2664 1769 2682 1787 ne
rect 2487 1693 2496 1727
rect 2530 1754 2572 1755
rect 2530 1720 2535 1754
rect 2565 1720 2572 1754
rect 2530 1711 2572 1720
rect 2606 1754 2648 1763
rect 2606 1720 2613 1754
rect 2643 1720 2648 1754
rect 2606 1715 2648 1720
rect 2682 1727 2710 1787
tri 2755 1774 2777 1796 se
rect 2777 1789 2792 1797
tri 2777 1774 2792 1789 nw
tri 2749 1768 2755 1774 se
rect 2755 1768 2764 1774
rect 2468 1683 2496 1693
tri 2496 1683 2520 1707 sw
rect 2414 1613 2430 1661
rect 2468 1651 2510 1683
tri 2527 1675 2528 1676 sw
rect 2527 1651 2528 1675
tri 2530 1674 2567 1711 ne
rect 2567 1683 2572 1711
tri 2572 1683 2598 1709 sw
rect 2682 1693 2691 1727
rect 2682 1683 2710 1693
rect 2567 1674 2651 1683
tri 2567 1655 2586 1674 ne
rect 2586 1655 2651 1674
rect 2468 1629 2528 1651
rect 2650 1651 2651 1655
rect 2668 1651 2710 1683
rect 2650 1629 2710 1651
rect 2556 1613 2573 1627
rect 2605 1613 2622 1627
tri 2393 1577 2415 1599 se
rect 2415 1592 2430 1613
tri 2415 1577 2430 1592 nw
rect 2749 1592 2764 1768
tri 2764 1761 2777 1774 nw
rect 2850 1693 2865 1921
tri 2387 1571 2393 1577 se
rect 2393 1571 2402 1577
rect 2387 1555 2402 1571
tri 2402 1564 2415 1577 nw
rect 2556 1569 2573 1583
rect 2605 1569 2622 1583
tri 2749 1577 2764 1592 ne
tri 2764 1577 2786 1599 sw
rect 2387 1519 2402 1527
rect 2468 1555 2528 1569
rect 2483 1545 2528 1555
rect 2483 1527 2511 1545
tri 2387 1504 2402 1519 ne
tri 2402 1504 2424 1526 sw
rect 2468 1517 2511 1527
rect 2526 1541 2528 1545
rect 2650 1555 2710 1569
tri 2764 1564 2777 1577 ne
rect 2777 1571 2786 1577
tri 2786 1571 2792 1577 sw
rect 2650 1545 2695 1555
rect 2526 1517 2600 1541
rect 2468 1513 2600 1517
tri 2600 1513 2628 1541 sw
rect 2650 1531 2652 1545
tri 2650 1529 2652 1531 ne
rect 2664 1527 2695 1545
rect 2664 1517 2710 1527
rect 2777 1556 2792 1571
tri 2402 1492 2414 1504 ne
rect 2414 1499 2424 1504
tri 2424 1499 2429 1504 sw
rect 2313 1153 2328 1381
rect 2414 1343 2429 1499
rect 2468 1457 2496 1513
tri 2588 1495 2606 1513 ne
rect 2606 1493 2628 1513
tri 2628 1493 2648 1513 sw
tri 2664 1499 2682 1517 ne
rect 2487 1423 2496 1457
rect 2530 1484 2572 1485
rect 2530 1450 2535 1484
rect 2565 1450 2572 1484
rect 2530 1441 2572 1450
rect 2606 1484 2648 1493
rect 2606 1450 2613 1484
rect 2643 1450 2648 1484
rect 2606 1445 2648 1450
rect 2682 1457 2710 1517
tri 2755 1504 2777 1526 se
rect 2777 1519 2792 1527
tri 2777 1504 2792 1519 nw
tri 2749 1498 2755 1504 se
rect 2755 1498 2764 1504
rect 2468 1413 2496 1423
tri 2496 1413 2520 1437 sw
rect 2468 1381 2510 1413
tri 2527 1405 2528 1406 sw
rect 2527 1381 2528 1405
tri 2530 1404 2567 1441 ne
rect 2567 1413 2572 1441
tri 2572 1413 2598 1439 sw
rect 2682 1423 2691 1457
rect 2682 1413 2710 1423
rect 2567 1404 2651 1413
tri 2567 1385 2586 1404 ne
rect 2586 1385 2651 1404
rect 2468 1359 2528 1381
rect 2650 1381 2651 1385
rect 2668 1381 2710 1413
rect 2650 1359 2710 1381
rect 2556 1343 2573 1357
rect 2605 1343 2622 1357
tri 2393 1307 2415 1329 se
rect 2415 1322 2430 1343
tri 2415 1307 2430 1322 nw
rect 2749 1322 2764 1498
tri 2764 1491 2777 1504 nw
rect 2850 1423 2865 1651
tri 2387 1301 2393 1307 se
rect 2393 1301 2402 1307
rect 2387 1285 2402 1301
tri 2402 1294 2415 1307 nw
rect 2556 1299 2573 1313
rect 2605 1299 2622 1313
tri 2749 1307 2764 1322 ne
tri 2764 1307 2786 1329 sw
rect 2387 1249 2402 1257
rect 2468 1285 2528 1299
rect 2483 1275 2528 1285
rect 2483 1257 2511 1275
tri 2387 1234 2402 1249 ne
tri 2402 1234 2424 1256 sw
rect 2468 1247 2511 1257
rect 2526 1271 2528 1275
rect 2650 1285 2710 1299
tri 2764 1294 2777 1307 ne
rect 2777 1301 2786 1307
tri 2786 1301 2792 1307 sw
rect 2650 1275 2695 1285
rect 2526 1247 2600 1271
rect 2468 1243 2600 1247
tri 2600 1243 2628 1271 sw
rect 2650 1261 2652 1275
tri 2650 1259 2652 1261 ne
rect 2664 1257 2695 1275
rect 2664 1247 2710 1257
rect 2777 1286 2792 1301
tri 2402 1222 2414 1234 ne
rect 2414 1229 2424 1234
tri 2424 1229 2429 1234 sw
rect 2313 883 2328 1111
rect 2414 1121 2429 1229
rect 2468 1187 2496 1243
tri 2588 1225 2606 1243 ne
rect 2606 1223 2628 1243
tri 2628 1223 2648 1243 sw
tri 2664 1229 2682 1247 ne
rect 2487 1153 2496 1187
rect 2530 1214 2572 1215
rect 2530 1180 2535 1214
rect 2565 1180 2572 1214
rect 2530 1171 2572 1180
rect 2606 1214 2648 1223
rect 2606 1180 2613 1214
rect 2643 1180 2648 1214
rect 2606 1175 2648 1180
rect 2682 1187 2710 1247
tri 2755 1234 2777 1256 se
rect 2777 1249 2792 1257
tri 2777 1234 2792 1249 nw
tri 2749 1228 2755 1234 se
rect 2755 1228 2764 1234
rect 2468 1143 2496 1153
tri 2496 1143 2520 1167 sw
rect 2414 1073 2430 1121
rect 2468 1111 2510 1143
tri 2527 1135 2528 1136 sw
rect 2527 1111 2528 1135
tri 2530 1134 2567 1171 ne
rect 2567 1143 2572 1171
tri 2572 1143 2598 1169 sw
rect 2682 1153 2691 1187
rect 2682 1143 2710 1153
rect 2567 1134 2651 1143
tri 2567 1115 2586 1134 ne
rect 2586 1115 2651 1134
rect 2468 1089 2528 1111
rect 2650 1111 2651 1115
rect 2668 1111 2710 1143
rect 2650 1089 2710 1111
rect 2556 1073 2573 1087
rect 2605 1073 2622 1087
tri 2393 1037 2415 1059 se
rect 2415 1052 2430 1073
tri 2415 1037 2430 1052 nw
rect 2749 1052 2764 1228
tri 2764 1221 2777 1234 nw
rect 2850 1153 2865 1381
tri 2387 1031 2393 1037 se
rect 2393 1031 2402 1037
rect 2387 1015 2402 1031
tri 2402 1024 2415 1037 nw
rect 2556 1029 2573 1043
rect 2605 1029 2622 1043
tri 2749 1037 2764 1052 ne
tri 2764 1037 2786 1059 sw
rect 2387 979 2402 987
rect 2468 1015 2528 1029
rect 2483 1005 2528 1015
rect 2483 987 2511 1005
tri 2387 964 2402 979 ne
tri 2402 964 2424 986 sw
rect 2468 977 2511 987
rect 2526 1001 2528 1005
rect 2650 1015 2710 1029
tri 2764 1024 2777 1037 ne
rect 2777 1031 2786 1037
tri 2786 1031 2792 1037 sw
rect 2650 1005 2695 1015
rect 2526 977 2600 1001
rect 2468 973 2600 977
tri 2600 973 2628 1001 sw
rect 2650 991 2652 1005
tri 2650 989 2652 991 ne
rect 2664 987 2695 1005
rect 2664 977 2710 987
rect 2777 1016 2792 1031
tri 2402 952 2414 964 ne
rect 2414 959 2424 964
tri 2424 959 2429 964 sw
rect 2313 613 2328 841
rect 2414 803 2429 959
rect 2468 917 2496 973
tri 2588 955 2606 973 ne
rect 2606 953 2628 973
tri 2628 953 2648 973 sw
tri 2664 959 2682 977 ne
rect 2487 883 2496 917
rect 2530 944 2572 945
rect 2530 910 2535 944
rect 2565 910 2572 944
rect 2530 901 2572 910
rect 2606 944 2648 953
rect 2606 910 2613 944
rect 2643 910 2648 944
rect 2606 905 2648 910
rect 2682 917 2710 977
tri 2755 964 2777 986 se
rect 2777 979 2792 987
tri 2777 964 2792 979 nw
tri 2749 958 2755 964 se
rect 2755 958 2764 964
rect 2468 873 2496 883
tri 2496 873 2520 897 sw
rect 2468 841 2510 873
tri 2527 865 2528 866 sw
rect 2527 841 2528 865
tri 2530 864 2567 901 ne
rect 2567 873 2572 901
tri 2572 873 2598 899 sw
rect 2682 883 2691 917
rect 2682 873 2710 883
rect 2567 864 2651 873
tri 2567 845 2586 864 ne
rect 2586 845 2651 864
rect 2468 819 2528 841
rect 2650 841 2651 845
rect 2668 841 2710 873
rect 2650 819 2710 841
rect 2556 803 2573 817
rect 2605 803 2622 817
tri 2393 767 2415 789 se
rect 2415 782 2430 803
tri 2415 767 2430 782 nw
rect 2749 782 2764 958
tri 2764 951 2777 964 nw
rect 2850 883 2865 1111
tri 2387 761 2393 767 se
rect 2393 761 2402 767
rect 2387 745 2402 761
tri 2402 754 2415 767 nw
rect 2556 759 2573 773
rect 2605 759 2622 773
tri 2749 767 2764 782 ne
tri 2764 767 2786 789 sw
rect 2387 709 2402 717
rect 2468 745 2528 759
rect 2483 735 2528 745
rect 2483 717 2511 735
tri 2387 694 2402 709 ne
tri 2402 694 2424 716 sw
rect 2468 707 2511 717
rect 2526 731 2528 735
rect 2650 745 2710 759
tri 2764 754 2777 767 ne
rect 2777 761 2786 767
tri 2786 761 2792 767 sw
rect 2650 735 2695 745
rect 2526 707 2600 731
rect 2468 703 2600 707
tri 2600 703 2628 731 sw
rect 2650 721 2652 735
tri 2650 719 2652 721 ne
rect 2664 717 2695 735
rect 2664 707 2710 717
rect 2777 746 2792 761
tri 2402 682 2414 694 ne
rect 2414 689 2424 694
tri 2424 689 2429 694 sw
rect 2313 343 2328 571
rect 2414 581 2429 689
rect 2468 647 2496 703
tri 2588 685 2606 703 ne
rect 2606 683 2628 703
tri 2628 683 2648 703 sw
tri 2664 689 2682 707 ne
rect 2487 613 2496 647
rect 2530 674 2572 675
rect 2530 640 2535 674
rect 2565 640 2572 674
rect 2530 631 2572 640
rect 2606 674 2648 683
rect 2606 640 2613 674
rect 2643 640 2648 674
rect 2606 635 2648 640
rect 2682 647 2710 707
tri 2755 694 2777 716 se
rect 2777 709 2792 717
tri 2777 694 2792 709 nw
tri 2749 688 2755 694 se
rect 2755 688 2764 694
rect 2468 603 2496 613
tri 2496 603 2520 627 sw
rect 2414 533 2430 581
rect 2468 571 2510 603
tri 2527 595 2528 596 sw
rect 2527 571 2528 595
tri 2530 594 2567 631 ne
rect 2567 603 2572 631
tri 2572 603 2598 629 sw
rect 2682 613 2691 647
rect 2682 603 2710 613
rect 2567 594 2651 603
tri 2567 575 2586 594 ne
rect 2586 575 2651 594
rect 2468 549 2528 571
rect 2650 571 2651 575
rect 2668 571 2710 603
rect 2650 549 2710 571
rect 2556 533 2573 547
rect 2605 533 2622 547
tri 2393 497 2415 519 se
rect 2415 512 2430 533
tri 2415 497 2430 512 nw
rect 2749 512 2764 688
tri 2764 681 2777 694 nw
rect 2850 613 2865 841
tri 2387 491 2393 497 se
rect 2393 491 2402 497
rect 2387 475 2402 491
tri 2402 484 2415 497 nw
rect 2556 489 2573 503
rect 2605 489 2622 503
tri 2749 497 2764 512 ne
tri 2764 497 2786 519 sw
rect 2387 439 2402 447
rect 2468 475 2528 489
rect 2483 465 2528 475
rect 2483 447 2511 465
tri 2387 424 2402 439 ne
tri 2402 424 2424 446 sw
rect 2468 437 2511 447
rect 2526 461 2528 465
rect 2650 475 2710 489
tri 2764 484 2777 497 ne
rect 2777 491 2786 497
tri 2786 491 2792 497 sw
rect 2650 465 2695 475
rect 2526 437 2600 461
rect 2468 433 2600 437
tri 2600 433 2628 461 sw
rect 2650 451 2652 465
tri 2650 449 2652 451 ne
rect 2664 447 2695 465
rect 2664 437 2710 447
rect 2777 476 2792 491
tri 2402 412 2414 424 ne
rect 2414 419 2424 424
tri 2424 419 2429 424 sw
rect 2313 73 2328 301
rect 2414 263 2429 419
rect 2468 377 2496 433
tri 2588 415 2606 433 ne
rect 2606 413 2628 433
tri 2628 413 2648 433 sw
tri 2664 419 2682 437 ne
rect 2487 343 2496 377
rect 2530 404 2572 405
rect 2530 370 2535 404
rect 2565 370 2572 404
rect 2530 361 2572 370
rect 2606 404 2648 413
rect 2606 370 2613 404
rect 2643 370 2648 404
rect 2606 365 2648 370
rect 2682 377 2710 437
tri 2755 424 2777 446 se
rect 2777 439 2792 447
tri 2777 424 2792 439 nw
tri 2749 418 2755 424 se
rect 2755 418 2764 424
rect 2468 333 2496 343
tri 2496 333 2520 357 sw
rect 2468 301 2510 333
tri 2527 325 2528 326 sw
rect 2527 301 2528 325
tri 2530 324 2567 361 ne
rect 2567 333 2572 361
tri 2572 333 2598 359 sw
rect 2682 343 2691 377
rect 2682 333 2710 343
rect 2567 324 2651 333
tri 2567 305 2586 324 ne
rect 2586 305 2651 324
rect 2468 279 2528 301
rect 2650 301 2651 305
rect 2668 301 2710 333
rect 2650 279 2710 301
rect 2556 263 2573 277
rect 2605 263 2622 277
tri 2393 227 2415 249 se
rect 2415 242 2430 263
tri 2415 227 2430 242 nw
rect 2749 242 2764 418
tri 2764 411 2777 424 nw
rect 2850 343 2865 571
tri 2387 221 2393 227 se
rect 2393 221 2402 227
rect 2387 205 2402 221
tri 2402 214 2415 227 nw
rect 2556 219 2573 233
rect 2605 219 2622 233
tri 2749 227 2764 242 ne
tri 2764 227 2786 249 sw
rect 2387 169 2402 177
rect 2468 205 2528 219
rect 2483 195 2528 205
rect 2483 177 2511 195
tri 2387 154 2402 169 ne
tri 2402 154 2424 176 sw
rect 2468 167 2511 177
rect 2526 191 2528 195
rect 2650 205 2710 219
tri 2764 214 2777 227 ne
rect 2777 221 2786 227
tri 2786 221 2792 227 sw
rect 2650 195 2695 205
rect 2526 167 2600 191
rect 2468 163 2600 167
tri 2600 163 2628 191 sw
rect 2650 181 2652 195
tri 2650 179 2652 181 ne
rect 2664 177 2695 195
rect 2664 167 2710 177
rect 2777 206 2792 221
tri 2402 142 2414 154 ne
rect 2414 149 2424 154
tri 2424 149 2429 154 sw
rect 2313 -55 2328 31
rect 2414 -55 2429 149
rect 2468 107 2496 163
tri 2588 145 2606 163 ne
rect 2606 143 2628 163
tri 2628 143 2648 163 sw
tri 2664 149 2682 167 ne
rect 2487 73 2496 107
rect 2530 134 2572 135
rect 2530 100 2535 134
rect 2565 100 2572 134
rect 2530 91 2572 100
rect 2606 134 2648 143
rect 2606 100 2613 134
rect 2643 100 2648 134
rect 2606 95 2648 100
rect 2682 107 2710 167
tri 2755 154 2777 176 se
rect 2777 169 2792 177
tri 2777 154 2792 169 nw
tri 2749 148 2755 154 se
rect 2755 148 2764 154
rect 2468 63 2496 73
tri 2496 63 2520 87 sw
rect 2468 31 2510 63
tri 2527 55 2528 56 sw
rect 2527 31 2528 55
tri 2530 54 2567 91 ne
rect 2567 63 2572 91
tri 2572 63 2598 89 sw
rect 2682 73 2691 107
rect 2682 63 2710 73
rect 2567 54 2651 63
tri 2567 35 2586 54 ne
rect 2586 35 2651 54
rect 2468 9 2528 31
rect 2650 31 2651 35
rect 2668 31 2710 63
rect 2650 9 2710 31
rect 2556 -7 2573 7
rect 2605 -7 2622 7
rect 2749 -55 2764 148
tri 2764 141 2777 154 nw
rect 2850 73 2865 301
rect 2850 -55 2865 31
rect 2893 4123 2908 4361
tri 2973 4277 2995 4299 se
rect 2995 4292 3010 4361
tri 2995 4277 3010 4292 nw
rect 3329 4292 3344 4361
tri 2967 4271 2973 4277 se
rect 2973 4271 2982 4277
rect 2967 4255 2982 4271
tri 2982 4264 2995 4277 nw
rect 3136 4269 3153 4283
rect 3185 4269 3202 4283
tri 3329 4277 3344 4292 ne
tri 3344 4277 3366 4299 sw
rect 2967 4219 2982 4227
rect 3048 4255 3108 4269
rect 3063 4245 3108 4255
rect 3063 4227 3091 4245
tri 2967 4204 2982 4219 ne
tri 2982 4204 3004 4226 sw
rect 3048 4217 3091 4227
rect 3106 4241 3108 4245
rect 3230 4255 3290 4269
tri 3344 4264 3357 4277 ne
rect 3357 4271 3366 4277
tri 3366 4271 3372 4277 sw
rect 3230 4245 3275 4255
rect 3106 4217 3180 4241
rect 3048 4213 3180 4217
tri 3180 4213 3208 4241 sw
rect 3230 4231 3232 4245
tri 3230 4229 3232 4231 ne
rect 3244 4227 3275 4245
rect 3244 4217 3290 4227
rect 3357 4256 3372 4271
tri 2982 4192 2994 4204 ne
rect 2994 4199 3004 4204
tri 3004 4199 3009 4204 sw
rect 2893 3853 2908 4081
rect 2994 4043 3009 4199
rect 3048 4157 3076 4213
tri 3168 4195 3186 4213 ne
rect 3186 4193 3208 4213
tri 3208 4193 3228 4213 sw
tri 3244 4199 3262 4217 ne
rect 3067 4123 3076 4157
rect 3110 4184 3152 4185
rect 3110 4150 3115 4184
rect 3145 4150 3152 4184
rect 3110 4141 3152 4150
rect 3186 4184 3228 4193
rect 3186 4150 3193 4184
rect 3223 4150 3228 4184
rect 3186 4145 3228 4150
rect 3262 4157 3290 4217
tri 3335 4204 3357 4226 se
rect 3357 4219 3372 4227
tri 3357 4204 3372 4219 nw
tri 3329 4198 3335 4204 se
rect 3335 4198 3344 4204
rect 3048 4113 3076 4123
tri 3076 4113 3100 4137 sw
rect 3048 4081 3090 4113
tri 3107 4105 3108 4106 sw
rect 3107 4081 3108 4105
tri 3110 4104 3147 4141 ne
rect 3147 4113 3152 4141
tri 3152 4113 3178 4139 sw
rect 3262 4123 3271 4157
rect 3262 4113 3290 4123
rect 3147 4104 3231 4113
tri 3147 4085 3166 4104 ne
rect 3166 4085 3231 4104
rect 3048 4059 3108 4081
rect 3230 4081 3231 4085
rect 3248 4081 3290 4113
rect 3230 4059 3290 4081
rect 3136 4043 3153 4057
rect 3185 4043 3202 4057
tri 2973 4007 2995 4029 se
rect 2995 4022 3010 4043
tri 2995 4007 3010 4022 nw
rect 3329 4022 3344 4198
tri 3344 4191 3357 4204 nw
rect 3430 4123 3445 4361
tri 2967 4001 2973 4007 se
rect 2973 4001 2982 4007
rect 2967 3985 2982 4001
tri 2982 3994 2995 4007 nw
rect 3136 3999 3153 4013
rect 3185 3999 3202 4013
tri 3329 4007 3344 4022 ne
tri 3344 4007 3366 4029 sw
rect 2967 3949 2982 3957
rect 3048 3985 3108 3999
rect 3063 3975 3108 3985
rect 3063 3957 3091 3975
tri 2967 3934 2982 3949 ne
tri 2982 3934 3004 3956 sw
rect 3048 3947 3091 3957
rect 3106 3971 3108 3975
rect 3230 3985 3290 3999
tri 3344 3994 3357 4007 ne
rect 3357 4001 3366 4007
tri 3366 4001 3372 4007 sw
rect 3230 3975 3275 3985
rect 3106 3947 3180 3971
rect 3048 3943 3180 3947
tri 3180 3943 3208 3971 sw
rect 3230 3961 3232 3975
tri 3230 3959 3232 3961 ne
rect 3244 3957 3275 3975
rect 3244 3947 3290 3957
rect 3357 3986 3372 4001
tri 2982 3922 2994 3934 ne
rect 2994 3929 3004 3934
tri 3004 3929 3009 3934 sw
rect 2893 3583 2908 3811
rect 2994 3821 3009 3929
rect 3048 3887 3076 3943
tri 3168 3925 3186 3943 ne
rect 3186 3923 3208 3943
tri 3208 3923 3228 3943 sw
tri 3244 3929 3262 3947 ne
rect 3067 3853 3076 3887
rect 3110 3914 3152 3915
rect 3110 3880 3115 3914
rect 3145 3880 3152 3914
rect 3110 3871 3152 3880
rect 3186 3914 3228 3923
rect 3186 3880 3193 3914
rect 3223 3880 3228 3914
rect 3186 3875 3228 3880
rect 3262 3887 3290 3947
tri 3335 3934 3357 3956 se
rect 3357 3949 3372 3957
tri 3357 3934 3372 3949 nw
tri 3329 3928 3335 3934 se
rect 3335 3928 3344 3934
rect 3048 3843 3076 3853
tri 3076 3843 3100 3867 sw
rect 2994 3773 3010 3821
rect 3048 3811 3090 3843
tri 3107 3835 3108 3836 sw
rect 3107 3811 3108 3835
tri 3110 3834 3147 3871 ne
rect 3147 3843 3152 3871
tri 3152 3843 3178 3869 sw
rect 3262 3853 3271 3887
rect 3262 3843 3290 3853
rect 3147 3834 3231 3843
tri 3147 3815 3166 3834 ne
rect 3166 3815 3231 3834
rect 3048 3789 3108 3811
rect 3230 3811 3231 3815
rect 3248 3811 3290 3843
rect 3230 3789 3290 3811
rect 3136 3773 3153 3787
rect 3185 3773 3202 3787
tri 2973 3737 2995 3759 se
rect 2995 3752 3010 3773
tri 2995 3737 3010 3752 nw
rect 3329 3752 3344 3928
tri 3344 3921 3357 3934 nw
rect 3430 3853 3445 4081
tri 2967 3731 2973 3737 se
rect 2973 3731 2982 3737
rect 2967 3715 2982 3731
tri 2982 3724 2995 3737 nw
rect 3136 3729 3153 3743
rect 3185 3729 3202 3743
tri 3329 3737 3344 3752 ne
tri 3344 3737 3366 3759 sw
rect 2967 3679 2982 3687
rect 3048 3715 3108 3729
rect 3063 3705 3108 3715
rect 3063 3687 3091 3705
tri 2967 3664 2982 3679 ne
tri 2982 3664 3004 3686 sw
rect 3048 3677 3091 3687
rect 3106 3701 3108 3705
rect 3230 3715 3290 3729
tri 3344 3724 3357 3737 ne
rect 3357 3731 3366 3737
tri 3366 3731 3372 3737 sw
rect 3230 3705 3275 3715
rect 3106 3677 3180 3701
rect 3048 3673 3180 3677
tri 3180 3673 3208 3701 sw
rect 3230 3691 3232 3705
tri 3230 3689 3232 3691 ne
rect 3244 3687 3275 3705
rect 3244 3677 3290 3687
rect 3357 3716 3372 3731
tri 2982 3652 2994 3664 ne
rect 2994 3659 3004 3664
tri 3004 3659 3009 3664 sw
rect 2893 3313 2908 3541
rect 2994 3503 3009 3659
rect 3048 3617 3076 3673
tri 3168 3655 3186 3673 ne
rect 3186 3653 3208 3673
tri 3208 3653 3228 3673 sw
tri 3244 3659 3262 3677 ne
rect 3067 3583 3076 3617
rect 3110 3644 3152 3645
rect 3110 3610 3115 3644
rect 3145 3610 3152 3644
rect 3110 3601 3152 3610
rect 3186 3644 3228 3653
rect 3186 3610 3193 3644
rect 3223 3610 3228 3644
rect 3186 3605 3228 3610
rect 3262 3617 3290 3677
tri 3335 3664 3357 3686 se
rect 3357 3679 3372 3687
tri 3357 3664 3372 3679 nw
tri 3329 3658 3335 3664 se
rect 3335 3658 3344 3664
rect 3048 3573 3076 3583
tri 3076 3573 3100 3597 sw
rect 3048 3541 3090 3573
tri 3107 3565 3108 3566 sw
rect 3107 3541 3108 3565
tri 3110 3564 3147 3601 ne
rect 3147 3573 3152 3601
tri 3152 3573 3178 3599 sw
rect 3262 3583 3271 3617
rect 3262 3573 3290 3583
rect 3147 3564 3231 3573
tri 3147 3545 3166 3564 ne
rect 3166 3545 3231 3564
rect 3048 3519 3108 3541
rect 3230 3541 3231 3545
rect 3248 3541 3290 3573
rect 3230 3519 3290 3541
rect 3136 3503 3153 3517
rect 3185 3503 3202 3517
tri 2973 3467 2995 3489 se
rect 2995 3482 3010 3503
tri 2995 3467 3010 3482 nw
rect 3329 3482 3344 3658
tri 3344 3651 3357 3664 nw
rect 3430 3583 3445 3811
tri 2967 3461 2973 3467 se
rect 2973 3461 2982 3467
rect 2967 3445 2982 3461
tri 2982 3454 2995 3467 nw
rect 3136 3459 3153 3473
rect 3185 3459 3202 3473
tri 3329 3467 3344 3482 ne
tri 3344 3467 3366 3489 sw
rect 2967 3409 2982 3417
rect 3048 3445 3108 3459
rect 3063 3435 3108 3445
rect 3063 3417 3091 3435
tri 2967 3394 2982 3409 ne
tri 2982 3394 3004 3416 sw
rect 3048 3407 3091 3417
rect 3106 3431 3108 3435
rect 3230 3445 3290 3459
tri 3344 3454 3357 3467 ne
rect 3357 3461 3366 3467
tri 3366 3461 3372 3467 sw
rect 3230 3435 3275 3445
rect 3106 3407 3180 3431
rect 3048 3403 3180 3407
tri 3180 3403 3208 3431 sw
rect 3230 3421 3232 3435
tri 3230 3419 3232 3421 ne
rect 3244 3417 3275 3435
rect 3244 3407 3290 3417
rect 3357 3446 3372 3461
tri 2982 3382 2994 3394 ne
rect 2994 3389 3004 3394
tri 3004 3389 3009 3394 sw
rect 2893 3043 2908 3271
rect 2994 3281 3009 3389
rect 3048 3347 3076 3403
tri 3168 3385 3186 3403 ne
rect 3186 3383 3208 3403
tri 3208 3383 3228 3403 sw
tri 3244 3389 3262 3407 ne
rect 3067 3313 3076 3347
rect 3110 3374 3152 3375
rect 3110 3340 3115 3374
rect 3145 3340 3152 3374
rect 3110 3331 3152 3340
rect 3186 3374 3228 3383
rect 3186 3340 3193 3374
rect 3223 3340 3228 3374
rect 3186 3335 3228 3340
rect 3262 3347 3290 3407
tri 3335 3394 3357 3416 se
rect 3357 3409 3372 3417
tri 3357 3394 3372 3409 nw
tri 3329 3388 3335 3394 se
rect 3335 3388 3344 3394
rect 3048 3303 3076 3313
tri 3076 3303 3100 3327 sw
rect 2994 3233 3010 3281
rect 3048 3271 3090 3303
tri 3107 3295 3108 3296 sw
rect 3107 3271 3108 3295
tri 3110 3294 3147 3331 ne
rect 3147 3303 3152 3331
tri 3152 3303 3178 3329 sw
rect 3262 3313 3271 3347
rect 3262 3303 3290 3313
rect 3147 3294 3231 3303
tri 3147 3275 3166 3294 ne
rect 3166 3275 3231 3294
rect 3048 3249 3108 3271
rect 3230 3271 3231 3275
rect 3248 3271 3290 3303
rect 3230 3249 3290 3271
rect 3136 3233 3153 3247
rect 3185 3233 3202 3247
tri 2973 3197 2995 3219 se
rect 2995 3212 3010 3233
tri 2995 3197 3010 3212 nw
rect 3329 3212 3344 3388
tri 3344 3381 3357 3394 nw
rect 3430 3313 3445 3541
tri 2967 3191 2973 3197 se
rect 2973 3191 2982 3197
rect 2967 3175 2982 3191
tri 2982 3184 2995 3197 nw
rect 3136 3189 3153 3203
rect 3185 3189 3202 3203
tri 3329 3197 3344 3212 ne
tri 3344 3197 3366 3219 sw
rect 2967 3139 2982 3147
rect 3048 3175 3108 3189
rect 3063 3165 3108 3175
rect 3063 3147 3091 3165
tri 2967 3124 2982 3139 ne
tri 2982 3124 3004 3146 sw
rect 3048 3137 3091 3147
rect 3106 3161 3108 3165
rect 3230 3175 3290 3189
tri 3344 3184 3357 3197 ne
rect 3357 3191 3366 3197
tri 3366 3191 3372 3197 sw
rect 3230 3165 3275 3175
rect 3106 3137 3180 3161
rect 3048 3133 3180 3137
tri 3180 3133 3208 3161 sw
rect 3230 3151 3232 3165
tri 3230 3149 3232 3151 ne
rect 3244 3147 3275 3165
rect 3244 3137 3290 3147
rect 3357 3176 3372 3191
tri 2982 3112 2994 3124 ne
rect 2994 3119 3004 3124
tri 3004 3119 3009 3124 sw
rect 2893 2773 2908 3001
rect 2994 2963 3009 3119
rect 3048 3077 3076 3133
tri 3168 3115 3186 3133 ne
rect 3186 3113 3208 3133
tri 3208 3113 3228 3133 sw
tri 3244 3119 3262 3137 ne
rect 3067 3043 3076 3077
rect 3110 3104 3152 3105
rect 3110 3070 3115 3104
rect 3145 3070 3152 3104
rect 3110 3061 3152 3070
rect 3186 3104 3228 3113
rect 3186 3070 3193 3104
rect 3223 3070 3228 3104
rect 3186 3065 3228 3070
rect 3262 3077 3290 3137
tri 3335 3124 3357 3146 se
rect 3357 3139 3372 3147
tri 3357 3124 3372 3139 nw
tri 3329 3118 3335 3124 se
rect 3335 3118 3344 3124
rect 3048 3033 3076 3043
tri 3076 3033 3100 3057 sw
rect 3048 3001 3090 3033
tri 3107 3025 3108 3026 sw
rect 3107 3001 3108 3025
tri 3110 3024 3147 3061 ne
rect 3147 3033 3152 3061
tri 3152 3033 3178 3059 sw
rect 3262 3043 3271 3077
rect 3262 3033 3290 3043
rect 3147 3024 3231 3033
tri 3147 3005 3166 3024 ne
rect 3166 3005 3231 3024
rect 3048 2979 3108 3001
rect 3230 3001 3231 3005
rect 3248 3001 3290 3033
rect 3230 2979 3290 3001
rect 3136 2963 3153 2977
rect 3185 2963 3202 2977
tri 2973 2927 2995 2949 se
rect 2995 2942 3010 2963
tri 2995 2927 3010 2942 nw
rect 3329 2942 3344 3118
tri 3344 3111 3357 3124 nw
rect 3430 3043 3445 3271
tri 2967 2921 2973 2927 se
rect 2973 2921 2982 2927
rect 2967 2905 2982 2921
tri 2982 2914 2995 2927 nw
rect 3136 2919 3153 2933
rect 3185 2919 3202 2933
tri 3329 2927 3344 2942 ne
tri 3344 2927 3366 2949 sw
rect 2967 2869 2982 2877
rect 3048 2905 3108 2919
rect 3063 2895 3108 2905
rect 3063 2877 3091 2895
tri 2967 2854 2982 2869 ne
tri 2982 2854 3004 2876 sw
rect 3048 2867 3091 2877
rect 3106 2891 3108 2895
rect 3230 2905 3290 2919
tri 3344 2914 3357 2927 ne
rect 3357 2921 3366 2927
tri 3366 2921 3372 2927 sw
rect 3230 2895 3275 2905
rect 3106 2867 3180 2891
rect 3048 2863 3180 2867
tri 3180 2863 3208 2891 sw
rect 3230 2881 3232 2895
tri 3230 2879 3232 2881 ne
rect 3244 2877 3275 2895
rect 3244 2867 3290 2877
rect 3357 2906 3372 2921
tri 2982 2842 2994 2854 ne
rect 2994 2849 3004 2854
tri 3004 2849 3009 2854 sw
rect 2893 2503 2908 2731
rect 2994 2741 3009 2849
rect 3048 2807 3076 2863
tri 3168 2845 3186 2863 ne
rect 3186 2843 3208 2863
tri 3208 2843 3228 2863 sw
tri 3244 2849 3262 2867 ne
rect 3067 2773 3076 2807
rect 3110 2834 3152 2835
rect 3110 2800 3115 2834
rect 3145 2800 3152 2834
rect 3110 2791 3152 2800
rect 3186 2834 3228 2843
rect 3186 2800 3193 2834
rect 3223 2800 3228 2834
rect 3186 2795 3228 2800
rect 3262 2807 3290 2867
tri 3335 2854 3357 2876 se
rect 3357 2869 3372 2877
tri 3357 2854 3372 2869 nw
tri 3329 2848 3335 2854 se
rect 3335 2848 3344 2854
rect 3048 2763 3076 2773
tri 3076 2763 3100 2787 sw
rect 2994 2693 3010 2741
rect 3048 2731 3090 2763
tri 3107 2755 3108 2756 sw
rect 3107 2731 3108 2755
tri 3110 2754 3147 2791 ne
rect 3147 2763 3152 2791
tri 3152 2763 3178 2789 sw
rect 3262 2773 3271 2807
rect 3262 2763 3290 2773
rect 3147 2754 3231 2763
tri 3147 2735 3166 2754 ne
rect 3166 2735 3231 2754
rect 3048 2709 3108 2731
rect 3230 2731 3231 2735
rect 3248 2731 3290 2763
rect 3230 2709 3290 2731
rect 3136 2693 3153 2707
rect 3185 2693 3202 2707
tri 2973 2657 2995 2679 se
rect 2995 2672 3010 2693
tri 2995 2657 3010 2672 nw
rect 3329 2672 3344 2848
tri 3344 2841 3357 2854 nw
rect 3430 2773 3445 3001
tri 2967 2651 2973 2657 se
rect 2973 2651 2982 2657
rect 2967 2635 2982 2651
tri 2982 2644 2995 2657 nw
rect 3136 2649 3153 2663
rect 3185 2649 3202 2663
tri 3329 2657 3344 2672 ne
tri 3344 2657 3366 2679 sw
rect 2967 2599 2982 2607
rect 3048 2635 3108 2649
rect 3063 2625 3108 2635
rect 3063 2607 3091 2625
tri 2967 2584 2982 2599 ne
tri 2982 2584 3004 2606 sw
rect 3048 2597 3091 2607
rect 3106 2621 3108 2625
rect 3230 2635 3290 2649
tri 3344 2644 3357 2657 ne
rect 3357 2651 3366 2657
tri 3366 2651 3372 2657 sw
rect 3230 2625 3275 2635
rect 3106 2597 3180 2621
rect 3048 2593 3180 2597
tri 3180 2593 3208 2621 sw
rect 3230 2611 3232 2625
tri 3230 2609 3232 2611 ne
rect 3244 2607 3275 2625
rect 3244 2597 3290 2607
rect 3357 2636 3372 2651
tri 2982 2572 2994 2584 ne
rect 2994 2579 3004 2584
tri 3004 2579 3009 2584 sw
rect 2893 2233 2908 2461
rect 2994 2423 3009 2579
rect 3048 2537 3076 2593
tri 3168 2575 3186 2593 ne
rect 3186 2573 3208 2593
tri 3208 2573 3228 2593 sw
tri 3244 2579 3262 2597 ne
rect 3067 2503 3076 2537
rect 3110 2564 3152 2565
rect 3110 2530 3115 2564
rect 3145 2530 3152 2564
rect 3110 2521 3152 2530
rect 3186 2564 3228 2573
rect 3186 2530 3193 2564
rect 3223 2530 3228 2564
rect 3186 2525 3228 2530
rect 3262 2537 3290 2597
tri 3335 2584 3357 2606 se
rect 3357 2599 3372 2607
tri 3357 2584 3372 2599 nw
tri 3329 2578 3335 2584 se
rect 3335 2578 3344 2584
rect 3048 2493 3076 2503
tri 3076 2493 3100 2517 sw
rect 3048 2461 3090 2493
tri 3107 2485 3108 2486 sw
rect 3107 2461 3108 2485
tri 3110 2484 3147 2521 ne
rect 3147 2493 3152 2521
tri 3152 2493 3178 2519 sw
rect 3262 2503 3271 2537
rect 3262 2493 3290 2503
rect 3147 2484 3231 2493
tri 3147 2465 3166 2484 ne
rect 3166 2465 3231 2484
rect 3048 2439 3108 2461
rect 3230 2461 3231 2465
rect 3248 2461 3290 2493
rect 3230 2439 3290 2461
rect 3136 2423 3153 2437
rect 3185 2423 3202 2437
tri 2973 2387 2995 2409 se
rect 2995 2402 3010 2423
tri 2995 2387 3010 2402 nw
rect 3329 2402 3344 2578
tri 3344 2571 3357 2584 nw
rect 3430 2503 3445 2731
tri 2967 2381 2973 2387 se
rect 2973 2381 2982 2387
rect 2967 2365 2982 2381
tri 2982 2374 2995 2387 nw
rect 3136 2379 3153 2393
rect 3185 2379 3202 2393
tri 3329 2387 3344 2402 ne
tri 3344 2387 3366 2409 sw
rect 2967 2329 2982 2337
rect 3048 2365 3108 2379
rect 3063 2355 3108 2365
rect 3063 2337 3091 2355
tri 2967 2314 2982 2329 ne
tri 2982 2314 3004 2336 sw
rect 3048 2327 3091 2337
rect 3106 2351 3108 2355
rect 3230 2365 3290 2379
tri 3344 2374 3357 2387 ne
rect 3357 2381 3366 2387
tri 3366 2381 3372 2387 sw
rect 3230 2355 3275 2365
rect 3106 2327 3180 2351
rect 3048 2323 3180 2327
tri 3180 2323 3208 2351 sw
rect 3230 2341 3232 2355
tri 3230 2339 3232 2341 ne
rect 3244 2337 3275 2355
rect 3244 2327 3290 2337
rect 3357 2366 3372 2381
tri 2982 2302 2994 2314 ne
rect 2994 2309 3004 2314
tri 3004 2309 3009 2314 sw
rect 2893 1963 2908 2191
rect 2994 2201 3009 2309
rect 3048 2267 3076 2323
tri 3168 2305 3186 2323 ne
rect 3186 2303 3208 2323
tri 3208 2303 3228 2323 sw
tri 3244 2309 3262 2327 ne
rect 3067 2233 3076 2267
rect 3110 2294 3152 2295
rect 3110 2260 3115 2294
rect 3145 2260 3152 2294
rect 3110 2251 3152 2260
rect 3186 2294 3228 2303
rect 3186 2260 3193 2294
rect 3223 2260 3228 2294
rect 3186 2255 3228 2260
rect 3262 2267 3290 2327
tri 3335 2314 3357 2336 se
rect 3357 2329 3372 2337
tri 3357 2314 3372 2329 nw
tri 3329 2308 3335 2314 se
rect 3335 2308 3344 2314
rect 3048 2223 3076 2233
tri 3076 2223 3100 2247 sw
rect 2994 2153 3010 2201
rect 3048 2191 3090 2223
tri 3107 2215 3108 2216 sw
rect 3107 2191 3108 2215
tri 3110 2214 3147 2251 ne
rect 3147 2223 3152 2251
tri 3152 2223 3178 2249 sw
rect 3262 2233 3271 2267
rect 3262 2223 3290 2233
rect 3147 2214 3231 2223
tri 3147 2195 3166 2214 ne
rect 3166 2195 3231 2214
rect 3048 2169 3108 2191
rect 3230 2191 3231 2195
rect 3248 2191 3290 2223
rect 3230 2169 3290 2191
rect 3136 2153 3153 2167
rect 3185 2153 3202 2167
tri 2973 2117 2995 2139 se
rect 2995 2132 3010 2153
tri 2995 2117 3010 2132 nw
rect 3329 2132 3344 2308
tri 3344 2301 3357 2314 nw
rect 3430 2233 3445 2461
tri 2967 2111 2973 2117 se
rect 2973 2111 2982 2117
rect 2967 2095 2982 2111
tri 2982 2104 2995 2117 nw
rect 3136 2109 3153 2123
rect 3185 2109 3202 2123
tri 3329 2117 3344 2132 ne
tri 3344 2117 3366 2139 sw
rect 2967 2059 2982 2067
rect 3048 2095 3108 2109
rect 3063 2085 3108 2095
rect 3063 2067 3091 2085
tri 2967 2044 2982 2059 ne
tri 2982 2044 3004 2066 sw
rect 3048 2057 3091 2067
rect 3106 2081 3108 2085
rect 3230 2095 3290 2109
tri 3344 2104 3357 2117 ne
rect 3357 2111 3366 2117
tri 3366 2111 3372 2117 sw
rect 3230 2085 3275 2095
rect 3106 2057 3180 2081
rect 3048 2053 3180 2057
tri 3180 2053 3208 2081 sw
rect 3230 2071 3232 2085
tri 3230 2069 3232 2071 ne
rect 3244 2067 3275 2085
rect 3244 2057 3290 2067
rect 3357 2096 3372 2111
tri 2982 2032 2994 2044 ne
rect 2994 2039 3004 2044
tri 3004 2039 3009 2044 sw
rect 2893 1693 2908 1921
rect 2994 1883 3009 2039
rect 3048 1997 3076 2053
tri 3168 2035 3186 2053 ne
rect 3186 2033 3208 2053
tri 3208 2033 3228 2053 sw
tri 3244 2039 3262 2057 ne
rect 3067 1963 3076 1997
rect 3110 2024 3152 2025
rect 3110 1990 3115 2024
rect 3145 1990 3152 2024
rect 3110 1981 3152 1990
rect 3186 2024 3228 2033
rect 3186 1990 3193 2024
rect 3223 1990 3228 2024
rect 3186 1985 3228 1990
rect 3262 1997 3290 2057
tri 3335 2044 3357 2066 se
rect 3357 2059 3372 2067
tri 3357 2044 3372 2059 nw
tri 3329 2038 3335 2044 se
rect 3335 2038 3344 2044
rect 3048 1953 3076 1963
tri 3076 1953 3100 1977 sw
rect 3048 1921 3090 1953
tri 3107 1945 3108 1946 sw
rect 3107 1921 3108 1945
tri 3110 1944 3147 1981 ne
rect 3147 1953 3152 1981
tri 3152 1953 3178 1979 sw
rect 3262 1963 3271 1997
rect 3262 1953 3290 1963
rect 3147 1944 3231 1953
tri 3147 1925 3166 1944 ne
rect 3166 1925 3231 1944
rect 3048 1899 3108 1921
rect 3230 1921 3231 1925
rect 3248 1921 3290 1953
rect 3230 1899 3290 1921
rect 3136 1883 3153 1897
rect 3185 1883 3202 1897
tri 2973 1847 2995 1869 se
rect 2995 1862 3010 1883
tri 2995 1847 3010 1862 nw
rect 3329 1862 3344 2038
tri 3344 2031 3357 2044 nw
rect 3430 1963 3445 2191
tri 2967 1841 2973 1847 se
rect 2973 1841 2982 1847
rect 2967 1825 2982 1841
tri 2982 1834 2995 1847 nw
rect 3136 1839 3153 1853
rect 3185 1839 3202 1853
tri 3329 1847 3344 1862 ne
tri 3344 1847 3366 1869 sw
rect 2967 1789 2982 1797
rect 3048 1825 3108 1839
rect 3063 1815 3108 1825
rect 3063 1797 3091 1815
tri 2967 1774 2982 1789 ne
tri 2982 1774 3004 1796 sw
rect 3048 1787 3091 1797
rect 3106 1811 3108 1815
rect 3230 1825 3290 1839
tri 3344 1834 3357 1847 ne
rect 3357 1841 3366 1847
tri 3366 1841 3372 1847 sw
rect 3230 1815 3275 1825
rect 3106 1787 3180 1811
rect 3048 1783 3180 1787
tri 3180 1783 3208 1811 sw
rect 3230 1801 3232 1815
tri 3230 1799 3232 1801 ne
rect 3244 1797 3275 1815
rect 3244 1787 3290 1797
rect 3357 1826 3372 1841
tri 2982 1762 2994 1774 ne
rect 2994 1769 3004 1774
tri 3004 1769 3009 1774 sw
rect 2893 1423 2908 1651
rect 2994 1661 3009 1769
rect 3048 1727 3076 1783
tri 3168 1765 3186 1783 ne
rect 3186 1763 3208 1783
tri 3208 1763 3228 1783 sw
tri 3244 1769 3262 1787 ne
rect 3067 1693 3076 1727
rect 3110 1754 3152 1755
rect 3110 1720 3115 1754
rect 3145 1720 3152 1754
rect 3110 1711 3152 1720
rect 3186 1754 3228 1763
rect 3186 1720 3193 1754
rect 3223 1720 3228 1754
rect 3186 1715 3228 1720
rect 3262 1727 3290 1787
tri 3335 1774 3357 1796 se
rect 3357 1789 3372 1797
tri 3357 1774 3372 1789 nw
tri 3329 1768 3335 1774 se
rect 3335 1768 3344 1774
rect 3048 1683 3076 1693
tri 3076 1683 3100 1707 sw
rect 2994 1613 3010 1661
rect 3048 1651 3090 1683
tri 3107 1675 3108 1676 sw
rect 3107 1651 3108 1675
tri 3110 1674 3147 1711 ne
rect 3147 1683 3152 1711
tri 3152 1683 3178 1709 sw
rect 3262 1693 3271 1727
rect 3262 1683 3290 1693
rect 3147 1674 3231 1683
tri 3147 1655 3166 1674 ne
rect 3166 1655 3231 1674
rect 3048 1629 3108 1651
rect 3230 1651 3231 1655
rect 3248 1651 3290 1683
rect 3230 1629 3290 1651
rect 3136 1613 3153 1627
rect 3185 1613 3202 1627
tri 2973 1577 2995 1599 se
rect 2995 1592 3010 1613
tri 2995 1577 3010 1592 nw
rect 3329 1592 3344 1768
tri 3344 1761 3357 1774 nw
rect 3430 1693 3445 1921
tri 2967 1571 2973 1577 se
rect 2973 1571 2982 1577
rect 2967 1555 2982 1571
tri 2982 1564 2995 1577 nw
rect 3136 1569 3153 1583
rect 3185 1569 3202 1583
tri 3329 1577 3344 1592 ne
tri 3344 1577 3366 1599 sw
rect 2967 1519 2982 1527
rect 3048 1555 3108 1569
rect 3063 1545 3108 1555
rect 3063 1527 3091 1545
tri 2967 1504 2982 1519 ne
tri 2982 1504 3004 1526 sw
rect 3048 1517 3091 1527
rect 3106 1541 3108 1545
rect 3230 1555 3290 1569
tri 3344 1564 3357 1577 ne
rect 3357 1571 3366 1577
tri 3366 1571 3372 1577 sw
rect 3230 1545 3275 1555
rect 3106 1517 3180 1541
rect 3048 1513 3180 1517
tri 3180 1513 3208 1541 sw
rect 3230 1531 3232 1545
tri 3230 1529 3232 1531 ne
rect 3244 1527 3275 1545
rect 3244 1517 3290 1527
rect 3357 1556 3372 1571
tri 2982 1492 2994 1504 ne
rect 2994 1499 3004 1504
tri 3004 1499 3009 1504 sw
rect 2893 1153 2908 1381
rect 2994 1343 3009 1499
rect 3048 1457 3076 1513
tri 3168 1495 3186 1513 ne
rect 3186 1493 3208 1513
tri 3208 1493 3228 1513 sw
tri 3244 1499 3262 1517 ne
rect 3067 1423 3076 1457
rect 3110 1484 3152 1485
rect 3110 1450 3115 1484
rect 3145 1450 3152 1484
rect 3110 1441 3152 1450
rect 3186 1484 3228 1493
rect 3186 1450 3193 1484
rect 3223 1450 3228 1484
rect 3186 1445 3228 1450
rect 3262 1457 3290 1517
tri 3335 1504 3357 1526 se
rect 3357 1519 3372 1527
tri 3357 1504 3372 1519 nw
tri 3329 1498 3335 1504 se
rect 3335 1498 3344 1504
rect 3048 1413 3076 1423
tri 3076 1413 3100 1437 sw
rect 3048 1381 3090 1413
tri 3107 1405 3108 1406 sw
rect 3107 1381 3108 1405
tri 3110 1404 3147 1441 ne
rect 3147 1413 3152 1441
tri 3152 1413 3178 1439 sw
rect 3262 1423 3271 1457
rect 3262 1413 3290 1423
rect 3147 1404 3231 1413
tri 3147 1385 3166 1404 ne
rect 3166 1385 3231 1404
rect 3048 1359 3108 1381
rect 3230 1381 3231 1385
rect 3248 1381 3290 1413
rect 3230 1359 3290 1381
rect 3136 1343 3153 1357
rect 3185 1343 3202 1357
tri 2973 1307 2995 1329 se
rect 2995 1322 3010 1343
tri 2995 1307 3010 1322 nw
rect 3329 1322 3344 1498
tri 3344 1491 3357 1504 nw
rect 3430 1423 3445 1651
tri 2967 1301 2973 1307 se
rect 2973 1301 2982 1307
rect 2967 1285 2982 1301
tri 2982 1294 2995 1307 nw
rect 3136 1299 3153 1313
rect 3185 1299 3202 1313
tri 3329 1307 3344 1322 ne
tri 3344 1307 3366 1329 sw
rect 2967 1249 2982 1257
rect 3048 1285 3108 1299
rect 3063 1275 3108 1285
rect 3063 1257 3091 1275
tri 2967 1234 2982 1249 ne
tri 2982 1234 3004 1256 sw
rect 3048 1247 3091 1257
rect 3106 1271 3108 1275
rect 3230 1285 3290 1299
tri 3344 1294 3357 1307 ne
rect 3357 1301 3366 1307
tri 3366 1301 3372 1307 sw
rect 3230 1275 3275 1285
rect 3106 1247 3180 1271
rect 3048 1243 3180 1247
tri 3180 1243 3208 1271 sw
rect 3230 1261 3232 1275
tri 3230 1259 3232 1261 ne
rect 3244 1257 3275 1275
rect 3244 1247 3290 1257
rect 3357 1286 3372 1301
tri 2982 1222 2994 1234 ne
rect 2994 1229 3004 1234
tri 3004 1229 3009 1234 sw
rect 2893 883 2908 1111
rect 2994 1121 3009 1229
rect 3048 1187 3076 1243
tri 3168 1225 3186 1243 ne
rect 3186 1223 3208 1243
tri 3208 1223 3228 1243 sw
tri 3244 1229 3262 1247 ne
rect 3067 1153 3076 1187
rect 3110 1214 3152 1215
rect 3110 1180 3115 1214
rect 3145 1180 3152 1214
rect 3110 1171 3152 1180
rect 3186 1214 3228 1223
rect 3186 1180 3193 1214
rect 3223 1180 3228 1214
rect 3186 1175 3228 1180
rect 3262 1187 3290 1247
tri 3335 1234 3357 1256 se
rect 3357 1249 3372 1257
tri 3357 1234 3372 1249 nw
tri 3329 1228 3335 1234 se
rect 3335 1228 3344 1234
rect 3048 1143 3076 1153
tri 3076 1143 3100 1167 sw
rect 2994 1073 3010 1121
rect 3048 1111 3090 1143
tri 3107 1135 3108 1136 sw
rect 3107 1111 3108 1135
tri 3110 1134 3147 1171 ne
rect 3147 1143 3152 1171
tri 3152 1143 3178 1169 sw
rect 3262 1153 3271 1187
rect 3262 1143 3290 1153
rect 3147 1134 3231 1143
tri 3147 1115 3166 1134 ne
rect 3166 1115 3231 1134
rect 3048 1089 3108 1111
rect 3230 1111 3231 1115
rect 3248 1111 3290 1143
rect 3230 1089 3290 1111
rect 3136 1073 3153 1087
rect 3185 1073 3202 1087
tri 2973 1037 2995 1059 se
rect 2995 1052 3010 1073
tri 2995 1037 3010 1052 nw
rect 3329 1052 3344 1228
tri 3344 1221 3357 1234 nw
rect 3430 1153 3445 1381
tri 2967 1031 2973 1037 se
rect 2973 1031 2982 1037
rect 2967 1015 2982 1031
tri 2982 1024 2995 1037 nw
rect 3136 1029 3153 1043
rect 3185 1029 3202 1043
tri 3329 1037 3344 1052 ne
tri 3344 1037 3366 1059 sw
rect 2967 979 2982 987
rect 3048 1015 3108 1029
rect 3063 1005 3108 1015
rect 3063 987 3091 1005
tri 2967 964 2982 979 ne
tri 2982 964 3004 986 sw
rect 3048 977 3091 987
rect 3106 1001 3108 1005
rect 3230 1015 3290 1029
tri 3344 1024 3357 1037 ne
rect 3357 1031 3366 1037
tri 3366 1031 3372 1037 sw
rect 3230 1005 3275 1015
rect 3106 977 3180 1001
rect 3048 973 3180 977
tri 3180 973 3208 1001 sw
rect 3230 991 3232 1005
tri 3230 989 3232 991 ne
rect 3244 987 3275 1005
rect 3244 977 3290 987
rect 3357 1016 3372 1031
tri 2982 952 2994 964 ne
rect 2994 959 3004 964
tri 3004 959 3009 964 sw
rect 2893 613 2908 841
rect 2994 803 3009 959
rect 3048 917 3076 973
tri 3168 955 3186 973 ne
rect 3186 953 3208 973
tri 3208 953 3228 973 sw
tri 3244 959 3262 977 ne
rect 3067 883 3076 917
rect 3110 944 3152 945
rect 3110 910 3115 944
rect 3145 910 3152 944
rect 3110 901 3152 910
rect 3186 944 3228 953
rect 3186 910 3193 944
rect 3223 910 3228 944
rect 3186 905 3228 910
rect 3262 917 3290 977
tri 3335 964 3357 986 se
rect 3357 979 3372 987
tri 3357 964 3372 979 nw
tri 3329 958 3335 964 se
rect 3335 958 3344 964
rect 3048 873 3076 883
tri 3076 873 3100 897 sw
rect 3048 841 3090 873
tri 3107 865 3108 866 sw
rect 3107 841 3108 865
tri 3110 864 3147 901 ne
rect 3147 873 3152 901
tri 3152 873 3178 899 sw
rect 3262 883 3271 917
rect 3262 873 3290 883
rect 3147 864 3231 873
tri 3147 845 3166 864 ne
rect 3166 845 3231 864
rect 3048 819 3108 841
rect 3230 841 3231 845
rect 3248 841 3290 873
rect 3230 819 3290 841
rect 3136 803 3153 817
rect 3185 803 3202 817
tri 2973 767 2995 789 se
rect 2995 782 3010 803
tri 2995 767 3010 782 nw
rect 3329 782 3344 958
tri 3344 951 3357 964 nw
rect 3430 883 3445 1111
tri 2967 761 2973 767 se
rect 2973 761 2982 767
rect 2967 745 2982 761
tri 2982 754 2995 767 nw
rect 3136 759 3153 773
rect 3185 759 3202 773
tri 3329 767 3344 782 ne
tri 3344 767 3366 789 sw
rect 2967 709 2982 717
rect 3048 745 3108 759
rect 3063 735 3108 745
rect 3063 717 3091 735
tri 2967 694 2982 709 ne
tri 2982 694 3004 716 sw
rect 3048 707 3091 717
rect 3106 731 3108 735
rect 3230 745 3290 759
tri 3344 754 3357 767 ne
rect 3357 761 3366 767
tri 3366 761 3372 767 sw
rect 3230 735 3275 745
rect 3106 707 3180 731
rect 3048 703 3180 707
tri 3180 703 3208 731 sw
rect 3230 721 3232 735
tri 3230 719 3232 721 ne
rect 3244 717 3275 735
rect 3244 707 3290 717
rect 3357 746 3372 761
tri 2982 682 2994 694 ne
rect 2994 689 3004 694
tri 3004 689 3009 694 sw
rect 2893 343 2908 571
rect 2994 581 3009 689
rect 3048 647 3076 703
tri 3168 685 3186 703 ne
rect 3186 683 3208 703
tri 3208 683 3228 703 sw
tri 3244 689 3262 707 ne
rect 3067 613 3076 647
rect 3110 674 3152 675
rect 3110 640 3115 674
rect 3145 640 3152 674
rect 3110 631 3152 640
rect 3186 674 3228 683
rect 3186 640 3193 674
rect 3223 640 3228 674
rect 3186 635 3228 640
rect 3262 647 3290 707
tri 3335 694 3357 716 se
rect 3357 709 3372 717
tri 3357 694 3372 709 nw
tri 3329 688 3335 694 se
rect 3335 688 3344 694
rect 3048 603 3076 613
tri 3076 603 3100 627 sw
rect 2994 533 3010 581
rect 3048 571 3090 603
tri 3107 595 3108 596 sw
rect 3107 571 3108 595
tri 3110 594 3147 631 ne
rect 3147 603 3152 631
tri 3152 603 3178 629 sw
rect 3262 613 3271 647
rect 3262 603 3290 613
rect 3147 594 3231 603
tri 3147 575 3166 594 ne
rect 3166 575 3231 594
rect 3048 549 3108 571
rect 3230 571 3231 575
rect 3248 571 3290 603
rect 3230 549 3290 571
rect 3136 533 3153 547
rect 3185 533 3202 547
tri 2973 497 2995 519 se
rect 2995 512 3010 533
tri 2995 497 3010 512 nw
rect 3329 512 3344 688
tri 3344 681 3357 694 nw
rect 3430 613 3445 841
tri 2967 491 2973 497 se
rect 2973 491 2982 497
rect 2967 475 2982 491
tri 2982 484 2995 497 nw
rect 3136 489 3153 503
rect 3185 489 3202 503
tri 3329 497 3344 512 ne
tri 3344 497 3366 519 sw
rect 2967 439 2982 447
rect 3048 475 3108 489
rect 3063 465 3108 475
rect 3063 447 3091 465
tri 2967 424 2982 439 ne
tri 2982 424 3004 446 sw
rect 3048 437 3091 447
rect 3106 461 3108 465
rect 3230 475 3290 489
tri 3344 484 3357 497 ne
rect 3357 491 3366 497
tri 3366 491 3372 497 sw
rect 3230 465 3275 475
rect 3106 437 3180 461
rect 3048 433 3180 437
tri 3180 433 3208 461 sw
rect 3230 451 3232 465
tri 3230 449 3232 451 ne
rect 3244 447 3275 465
rect 3244 437 3290 447
rect 3357 476 3372 491
tri 2982 412 2994 424 ne
rect 2994 419 3004 424
tri 3004 419 3009 424 sw
rect 2893 73 2908 301
rect 2994 263 3009 419
rect 3048 377 3076 433
tri 3168 415 3186 433 ne
rect 3186 413 3208 433
tri 3208 413 3228 433 sw
tri 3244 419 3262 437 ne
rect 3067 343 3076 377
rect 3110 404 3152 405
rect 3110 370 3115 404
rect 3145 370 3152 404
rect 3110 361 3152 370
rect 3186 404 3228 413
rect 3186 370 3193 404
rect 3223 370 3228 404
rect 3186 365 3228 370
rect 3262 377 3290 437
tri 3335 424 3357 446 se
rect 3357 439 3372 447
tri 3357 424 3372 439 nw
tri 3329 418 3335 424 se
rect 3335 418 3344 424
rect 3048 333 3076 343
tri 3076 333 3100 357 sw
rect 3048 301 3090 333
tri 3107 325 3108 326 sw
rect 3107 301 3108 325
tri 3110 324 3147 361 ne
rect 3147 333 3152 361
tri 3152 333 3178 359 sw
rect 3262 343 3271 377
rect 3262 333 3290 343
rect 3147 324 3231 333
tri 3147 305 3166 324 ne
rect 3166 305 3231 324
rect 3048 279 3108 301
rect 3230 301 3231 305
rect 3248 301 3290 333
rect 3230 279 3290 301
rect 3136 263 3153 277
rect 3185 263 3202 277
tri 2973 227 2995 249 se
rect 2995 242 3010 263
tri 2995 227 3010 242 nw
rect 3329 242 3344 418
tri 3344 411 3357 424 nw
rect 3430 343 3445 571
tri 2967 221 2973 227 se
rect 2973 221 2982 227
rect 2967 205 2982 221
tri 2982 214 2995 227 nw
rect 3136 219 3153 233
rect 3185 219 3202 233
tri 3329 227 3344 242 ne
tri 3344 227 3366 249 sw
rect 2967 169 2982 177
rect 3048 205 3108 219
rect 3063 195 3108 205
rect 3063 177 3091 195
tri 2967 154 2982 169 ne
tri 2982 154 3004 176 sw
rect 3048 167 3091 177
rect 3106 191 3108 195
rect 3230 205 3290 219
tri 3344 214 3357 227 ne
rect 3357 221 3366 227
tri 3366 221 3372 227 sw
rect 3230 195 3275 205
rect 3106 167 3180 191
rect 3048 163 3180 167
tri 3180 163 3208 191 sw
rect 3230 181 3232 195
tri 3230 179 3232 181 ne
rect 3244 177 3275 195
rect 3244 167 3290 177
rect 3357 206 3372 221
tri 2982 142 2994 154 ne
rect 2994 149 3004 154
tri 3004 149 3009 154 sw
rect 2893 -55 2908 31
rect 2994 -55 3009 149
rect 3048 107 3076 163
tri 3168 145 3186 163 ne
rect 3186 143 3208 163
tri 3208 143 3228 163 sw
tri 3244 149 3262 167 ne
rect 3067 73 3076 107
rect 3110 134 3152 135
rect 3110 100 3115 134
rect 3145 100 3152 134
rect 3110 91 3152 100
rect 3186 134 3228 143
rect 3186 100 3193 134
rect 3223 100 3228 134
rect 3186 95 3228 100
rect 3262 107 3290 167
tri 3335 154 3357 176 se
rect 3357 169 3372 177
tri 3357 154 3372 169 nw
tri 3329 148 3335 154 se
rect 3335 148 3344 154
rect 3048 63 3076 73
tri 3076 63 3100 87 sw
rect 3048 31 3090 63
tri 3107 55 3108 56 sw
rect 3107 31 3108 55
tri 3110 54 3147 91 ne
rect 3147 63 3152 91
tri 3152 63 3178 89 sw
rect 3262 73 3271 107
rect 3262 63 3290 73
rect 3147 54 3231 63
tri 3147 35 3166 54 ne
rect 3166 35 3231 54
rect 3048 9 3108 31
rect 3230 31 3231 35
rect 3248 31 3290 63
rect 3230 9 3290 31
rect 3136 -7 3153 7
rect 3185 -7 3202 7
rect 3329 -55 3344 148
tri 3344 141 3357 154 nw
rect 3430 73 3445 301
rect 3430 -55 3445 31
rect 3473 4123 3488 4361
tri 3553 4277 3575 4299 se
rect 3575 4292 3590 4361
tri 3575 4277 3590 4292 nw
rect 3909 4292 3924 4361
tri 3547 4271 3553 4277 se
rect 3553 4271 3562 4277
rect 3547 4255 3562 4271
tri 3562 4264 3575 4277 nw
rect 3716 4269 3733 4283
rect 3765 4269 3782 4283
tri 3909 4277 3924 4292 ne
tri 3924 4277 3946 4299 sw
rect 3547 4219 3562 4227
rect 3628 4255 3688 4269
rect 3643 4245 3688 4255
rect 3643 4227 3671 4245
tri 3547 4204 3562 4219 ne
tri 3562 4204 3584 4226 sw
rect 3628 4217 3671 4227
rect 3686 4241 3688 4245
rect 3810 4255 3870 4269
tri 3924 4264 3937 4277 ne
rect 3937 4271 3946 4277
tri 3946 4271 3952 4277 sw
rect 3810 4245 3855 4255
rect 3686 4217 3760 4241
rect 3628 4213 3760 4217
tri 3760 4213 3788 4241 sw
rect 3810 4231 3812 4245
tri 3810 4229 3812 4231 ne
rect 3824 4227 3855 4245
rect 3824 4217 3870 4227
rect 3937 4256 3952 4271
tri 3562 4192 3574 4204 ne
rect 3574 4199 3584 4204
tri 3584 4199 3589 4204 sw
rect 3473 3853 3488 4081
rect 3574 4043 3589 4199
rect 3628 4157 3656 4213
tri 3748 4195 3766 4213 ne
rect 3766 4193 3788 4213
tri 3788 4193 3808 4213 sw
tri 3824 4199 3842 4217 ne
rect 3647 4123 3656 4157
rect 3690 4184 3732 4185
rect 3690 4150 3695 4184
rect 3725 4150 3732 4184
rect 3690 4141 3732 4150
rect 3766 4184 3808 4193
rect 3766 4150 3773 4184
rect 3803 4150 3808 4184
rect 3766 4145 3808 4150
rect 3842 4157 3870 4217
tri 3915 4204 3937 4226 se
rect 3937 4219 3952 4227
tri 3937 4204 3952 4219 nw
tri 3909 4198 3915 4204 se
rect 3915 4198 3924 4204
rect 3628 4113 3656 4123
tri 3656 4113 3680 4137 sw
rect 3628 4081 3670 4113
tri 3687 4105 3688 4106 sw
rect 3687 4081 3688 4105
tri 3690 4104 3727 4141 ne
rect 3727 4113 3732 4141
tri 3732 4113 3758 4139 sw
rect 3842 4123 3851 4157
rect 3842 4113 3870 4123
rect 3727 4104 3811 4113
tri 3727 4085 3746 4104 ne
rect 3746 4085 3811 4104
rect 3628 4059 3688 4081
rect 3810 4081 3811 4085
rect 3828 4081 3870 4113
rect 3810 4059 3870 4081
rect 3716 4043 3733 4057
rect 3765 4043 3782 4057
tri 3553 4007 3575 4029 se
rect 3575 4022 3590 4043
tri 3575 4007 3590 4022 nw
rect 3909 4022 3924 4198
tri 3924 4191 3937 4204 nw
rect 4010 4123 4025 4361
tri 3547 4001 3553 4007 se
rect 3553 4001 3562 4007
rect 3547 3985 3562 4001
tri 3562 3994 3575 4007 nw
rect 3716 3999 3733 4013
rect 3765 3999 3782 4013
tri 3909 4007 3924 4022 ne
tri 3924 4007 3946 4029 sw
rect 3547 3949 3562 3957
rect 3628 3985 3688 3999
rect 3643 3975 3688 3985
rect 3643 3957 3671 3975
tri 3547 3934 3562 3949 ne
tri 3562 3934 3584 3956 sw
rect 3628 3947 3671 3957
rect 3686 3971 3688 3975
rect 3810 3985 3870 3999
tri 3924 3994 3937 4007 ne
rect 3937 4001 3946 4007
tri 3946 4001 3952 4007 sw
rect 3810 3975 3855 3985
rect 3686 3947 3760 3971
rect 3628 3943 3760 3947
tri 3760 3943 3788 3971 sw
rect 3810 3961 3812 3975
tri 3810 3959 3812 3961 ne
rect 3824 3957 3855 3975
rect 3824 3947 3870 3957
rect 3937 3986 3952 4001
tri 3562 3922 3574 3934 ne
rect 3574 3929 3584 3934
tri 3584 3929 3589 3934 sw
rect 3473 3583 3488 3811
rect 3574 3821 3589 3929
rect 3628 3887 3656 3943
tri 3748 3925 3766 3943 ne
rect 3766 3923 3788 3943
tri 3788 3923 3808 3943 sw
tri 3824 3929 3842 3947 ne
rect 3647 3853 3656 3887
rect 3690 3914 3732 3915
rect 3690 3880 3695 3914
rect 3725 3880 3732 3914
rect 3690 3871 3732 3880
rect 3766 3914 3808 3923
rect 3766 3880 3773 3914
rect 3803 3880 3808 3914
rect 3766 3875 3808 3880
rect 3842 3887 3870 3947
tri 3915 3934 3937 3956 se
rect 3937 3949 3952 3957
tri 3937 3934 3952 3949 nw
tri 3909 3928 3915 3934 se
rect 3915 3928 3924 3934
rect 3628 3843 3656 3853
tri 3656 3843 3680 3867 sw
rect 3574 3773 3590 3821
rect 3628 3811 3670 3843
tri 3687 3835 3688 3836 sw
rect 3687 3811 3688 3835
tri 3690 3834 3727 3871 ne
rect 3727 3843 3732 3871
tri 3732 3843 3758 3869 sw
rect 3842 3853 3851 3887
rect 3842 3843 3870 3853
rect 3727 3834 3811 3843
tri 3727 3815 3746 3834 ne
rect 3746 3815 3811 3834
rect 3628 3789 3688 3811
rect 3810 3811 3811 3815
rect 3828 3811 3870 3843
rect 3810 3789 3870 3811
rect 3716 3773 3733 3787
rect 3765 3773 3782 3787
tri 3553 3737 3575 3759 se
rect 3575 3752 3590 3773
tri 3575 3737 3590 3752 nw
rect 3909 3752 3924 3928
tri 3924 3921 3937 3934 nw
rect 4010 3853 4025 4081
tri 3547 3731 3553 3737 se
rect 3553 3731 3562 3737
rect 3547 3715 3562 3731
tri 3562 3724 3575 3737 nw
rect 3716 3729 3733 3743
rect 3765 3729 3782 3743
tri 3909 3737 3924 3752 ne
tri 3924 3737 3946 3759 sw
rect 3547 3679 3562 3687
rect 3628 3715 3688 3729
rect 3643 3705 3688 3715
rect 3643 3687 3671 3705
tri 3547 3664 3562 3679 ne
tri 3562 3664 3584 3686 sw
rect 3628 3677 3671 3687
rect 3686 3701 3688 3705
rect 3810 3715 3870 3729
tri 3924 3724 3937 3737 ne
rect 3937 3731 3946 3737
tri 3946 3731 3952 3737 sw
rect 3810 3705 3855 3715
rect 3686 3677 3760 3701
rect 3628 3673 3760 3677
tri 3760 3673 3788 3701 sw
rect 3810 3691 3812 3705
tri 3810 3689 3812 3691 ne
rect 3824 3687 3855 3705
rect 3824 3677 3870 3687
rect 3937 3716 3952 3731
tri 3562 3652 3574 3664 ne
rect 3574 3659 3584 3664
tri 3584 3659 3589 3664 sw
rect 3473 3313 3488 3541
rect 3574 3503 3589 3659
rect 3628 3617 3656 3673
tri 3748 3655 3766 3673 ne
rect 3766 3653 3788 3673
tri 3788 3653 3808 3673 sw
tri 3824 3659 3842 3677 ne
rect 3647 3583 3656 3617
rect 3690 3644 3732 3645
rect 3690 3610 3695 3644
rect 3725 3610 3732 3644
rect 3690 3601 3732 3610
rect 3766 3644 3808 3653
rect 3766 3610 3773 3644
rect 3803 3610 3808 3644
rect 3766 3605 3808 3610
rect 3842 3617 3870 3677
tri 3915 3664 3937 3686 se
rect 3937 3679 3952 3687
tri 3937 3664 3952 3679 nw
tri 3909 3658 3915 3664 se
rect 3915 3658 3924 3664
rect 3628 3573 3656 3583
tri 3656 3573 3680 3597 sw
rect 3628 3541 3670 3573
tri 3687 3565 3688 3566 sw
rect 3687 3541 3688 3565
tri 3690 3564 3727 3601 ne
rect 3727 3573 3732 3601
tri 3732 3573 3758 3599 sw
rect 3842 3583 3851 3617
rect 3842 3573 3870 3583
rect 3727 3564 3811 3573
tri 3727 3545 3746 3564 ne
rect 3746 3545 3811 3564
rect 3628 3519 3688 3541
rect 3810 3541 3811 3545
rect 3828 3541 3870 3573
rect 3810 3519 3870 3541
rect 3716 3503 3733 3517
rect 3765 3503 3782 3517
tri 3553 3467 3575 3489 se
rect 3575 3482 3590 3503
tri 3575 3467 3590 3482 nw
rect 3909 3482 3924 3658
tri 3924 3651 3937 3664 nw
rect 4010 3583 4025 3811
tri 3547 3461 3553 3467 se
rect 3553 3461 3562 3467
rect 3547 3445 3562 3461
tri 3562 3454 3575 3467 nw
rect 3716 3459 3733 3473
rect 3765 3459 3782 3473
tri 3909 3467 3924 3482 ne
tri 3924 3467 3946 3489 sw
rect 3547 3409 3562 3417
rect 3628 3445 3688 3459
rect 3643 3435 3688 3445
rect 3643 3417 3671 3435
tri 3547 3394 3562 3409 ne
tri 3562 3394 3584 3416 sw
rect 3628 3407 3671 3417
rect 3686 3431 3688 3435
rect 3810 3445 3870 3459
tri 3924 3454 3937 3467 ne
rect 3937 3461 3946 3467
tri 3946 3461 3952 3467 sw
rect 3810 3435 3855 3445
rect 3686 3407 3760 3431
rect 3628 3403 3760 3407
tri 3760 3403 3788 3431 sw
rect 3810 3421 3812 3435
tri 3810 3419 3812 3421 ne
rect 3824 3417 3855 3435
rect 3824 3407 3870 3417
rect 3937 3446 3952 3461
tri 3562 3382 3574 3394 ne
rect 3574 3389 3584 3394
tri 3584 3389 3589 3394 sw
rect 3473 3043 3488 3271
rect 3574 3281 3589 3389
rect 3628 3347 3656 3403
tri 3748 3385 3766 3403 ne
rect 3766 3383 3788 3403
tri 3788 3383 3808 3403 sw
tri 3824 3389 3842 3407 ne
rect 3647 3313 3656 3347
rect 3690 3374 3732 3375
rect 3690 3340 3695 3374
rect 3725 3340 3732 3374
rect 3690 3331 3732 3340
rect 3766 3374 3808 3383
rect 3766 3340 3773 3374
rect 3803 3340 3808 3374
rect 3766 3335 3808 3340
rect 3842 3347 3870 3407
tri 3915 3394 3937 3416 se
rect 3937 3409 3952 3417
tri 3937 3394 3952 3409 nw
tri 3909 3388 3915 3394 se
rect 3915 3388 3924 3394
rect 3628 3303 3656 3313
tri 3656 3303 3680 3327 sw
rect 3574 3233 3590 3281
rect 3628 3271 3670 3303
tri 3687 3295 3688 3296 sw
rect 3687 3271 3688 3295
tri 3690 3294 3727 3331 ne
rect 3727 3303 3732 3331
tri 3732 3303 3758 3329 sw
rect 3842 3313 3851 3347
rect 3842 3303 3870 3313
rect 3727 3294 3811 3303
tri 3727 3275 3746 3294 ne
rect 3746 3275 3811 3294
rect 3628 3249 3688 3271
rect 3810 3271 3811 3275
rect 3828 3271 3870 3303
rect 3810 3249 3870 3271
rect 3716 3233 3733 3247
rect 3765 3233 3782 3247
tri 3553 3197 3575 3219 se
rect 3575 3212 3590 3233
tri 3575 3197 3590 3212 nw
rect 3909 3212 3924 3388
tri 3924 3381 3937 3394 nw
rect 4010 3313 4025 3541
tri 3547 3191 3553 3197 se
rect 3553 3191 3562 3197
rect 3547 3175 3562 3191
tri 3562 3184 3575 3197 nw
rect 3716 3189 3733 3203
rect 3765 3189 3782 3203
tri 3909 3197 3924 3212 ne
tri 3924 3197 3946 3219 sw
rect 3547 3139 3562 3147
rect 3628 3175 3688 3189
rect 3643 3165 3688 3175
rect 3643 3147 3671 3165
tri 3547 3124 3562 3139 ne
tri 3562 3124 3584 3146 sw
rect 3628 3137 3671 3147
rect 3686 3161 3688 3165
rect 3810 3175 3870 3189
tri 3924 3184 3937 3197 ne
rect 3937 3191 3946 3197
tri 3946 3191 3952 3197 sw
rect 3810 3165 3855 3175
rect 3686 3137 3760 3161
rect 3628 3133 3760 3137
tri 3760 3133 3788 3161 sw
rect 3810 3151 3812 3165
tri 3810 3149 3812 3151 ne
rect 3824 3147 3855 3165
rect 3824 3137 3870 3147
rect 3937 3176 3952 3191
tri 3562 3112 3574 3124 ne
rect 3574 3119 3584 3124
tri 3584 3119 3589 3124 sw
rect 3473 2773 3488 3001
rect 3574 2963 3589 3119
rect 3628 3077 3656 3133
tri 3748 3115 3766 3133 ne
rect 3766 3113 3788 3133
tri 3788 3113 3808 3133 sw
tri 3824 3119 3842 3137 ne
rect 3647 3043 3656 3077
rect 3690 3104 3732 3105
rect 3690 3070 3695 3104
rect 3725 3070 3732 3104
rect 3690 3061 3732 3070
rect 3766 3104 3808 3113
rect 3766 3070 3773 3104
rect 3803 3070 3808 3104
rect 3766 3065 3808 3070
rect 3842 3077 3870 3137
tri 3915 3124 3937 3146 se
rect 3937 3139 3952 3147
tri 3937 3124 3952 3139 nw
tri 3909 3118 3915 3124 se
rect 3915 3118 3924 3124
rect 3628 3033 3656 3043
tri 3656 3033 3680 3057 sw
rect 3628 3001 3670 3033
tri 3687 3025 3688 3026 sw
rect 3687 3001 3688 3025
tri 3690 3024 3727 3061 ne
rect 3727 3033 3732 3061
tri 3732 3033 3758 3059 sw
rect 3842 3043 3851 3077
rect 3842 3033 3870 3043
rect 3727 3024 3811 3033
tri 3727 3005 3746 3024 ne
rect 3746 3005 3811 3024
rect 3628 2979 3688 3001
rect 3810 3001 3811 3005
rect 3828 3001 3870 3033
rect 3810 2979 3870 3001
rect 3716 2963 3733 2977
rect 3765 2963 3782 2977
tri 3553 2927 3575 2949 se
rect 3575 2942 3590 2963
tri 3575 2927 3590 2942 nw
rect 3909 2942 3924 3118
tri 3924 3111 3937 3124 nw
rect 4010 3043 4025 3271
tri 3547 2921 3553 2927 se
rect 3553 2921 3562 2927
rect 3547 2905 3562 2921
tri 3562 2914 3575 2927 nw
rect 3716 2919 3733 2933
rect 3765 2919 3782 2933
tri 3909 2927 3924 2942 ne
tri 3924 2927 3946 2949 sw
rect 3547 2869 3562 2877
rect 3628 2905 3688 2919
rect 3643 2895 3688 2905
rect 3643 2877 3671 2895
tri 3547 2854 3562 2869 ne
tri 3562 2854 3584 2876 sw
rect 3628 2867 3671 2877
rect 3686 2891 3688 2895
rect 3810 2905 3870 2919
tri 3924 2914 3937 2927 ne
rect 3937 2921 3946 2927
tri 3946 2921 3952 2927 sw
rect 3810 2895 3855 2905
rect 3686 2867 3760 2891
rect 3628 2863 3760 2867
tri 3760 2863 3788 2891 sw
rect 3810 2881 3812 2895
tri 3810 2879 3812 2881 ne
rect 3824 2877 3855 2895
rect 3824 2867 3870 2877
rect 3937 2906 3952 2921
tri 3562 2842 3574 2854 ne
rect 3574 2849 3584 2854
tri 3584 2849 3589 2854 sw
rect 3473 2503 3488 2731
rect 3574 2741 3589 2849
rect 3628 2807 3656 2863
tri 3748 2845 3766 2863 ne
rect 3766 2843 3788 2863
tri 3788 2843 3808 2863 sw
tri 3824 2849 3842 2867 ne
rect 3647 2773 3656 2807
rect 3690 2834 3732 2835
rect 3690 2800 3695 2834
rect 3725 2800 3732 2834
rect 3690 2791 3732 2800
rect 3766 2834 3808 2843
rect 3766 2800 3773 2834
rect 3803 2800 3808 2834
rect 3766 2795 3808 2800
rect 3842 2807 3870 2867
tri 3915 2854 3937 2876 se
rect 3937 2869 3952 2877
tri 3937 2854 3952 2869 nw
tri 3909 2848 3915 2854 se
rect 3915 2848 3924 2854
rect 3628 2763 3656 2773
tri 3656 2763 3680 2787 sw
rect 3574 2693 3590 2741
rect 3628 2731 3670 2763
tri 3687 2755 3688 2756 sw
rect 3687 2731 3688 2755
tri 3690 2754 3727 2791 ne
rect 3727 2763 3732 2791
tri 3732 2763 3758 2789 sw
rect 3842 2773 3851 2807
rect 3842 2763 3870 2773
rect 3727 2754 3811 2763
tri 3727 2735 3746 2754 ne
rect 3746 2735 3811 2754
rect 3628 2709 3688 2731
rect 3810 2731 3811 2735
rect 3828 2731 3870 2763
rect 3810 2709 3870 2731
rect 3716 2693 3733 2707
rect 3765 2693 3782 2707
tri 3553 2657 3575 2679 se
rect 3575 2672 3590 2693
tri 3575 2657 3590 2672 nw
rect 3909 2672 3924 2848
tri 3924 2841 3937 2854 nw
rect 4010 2773 4025 3001
tri 3547 2651 3553 2657 se
rect 3553 2651 3562 2657
rect 3547 2635 3562 2651
tri 3562 2644 3575 2657 nw
rect 3716 2649 3733 2663
rect 3765 2649 3782 2663
tri 3909 2657 3924 2672 ne
tri 3924 2657 3946 2679 sw
rect 3547 2599 3562 2607
rect 3628 2635 3688 2649
rect 3643 2625 3688 2635
rect 3643 2607 3671 2625
tri 3547 2584 3562 2599 ne
tri 3562 2584 3584 2606 sw
rect 3628 2597 3671 2607
rect 3686 2621 3688 2625
rect 3810 2635 3870 2649
tri 3924 2644 3937 2657 ne
rect 3937 2651 3946 2657
tri 3946 2651 3952 2657 sw
rect 3810 2625 3855 2635
rect 3686 2597 3760 2621
rect 3628 2593 3760 2597
tri 3760 2593 3788 2621 sw
rect 3810 2611 3812 2625
tri 3810 2609 3812 2611 ne
rect 3824 2607 3855 2625
rect 3824 2597 3870 2607
rect 3937 2636 3952 2651
tri 3562 2572 3574 2584 ne
rect 3574 2579 3584 2584
tri 3584 2579 3589 2584 sw
rect 3473 2233 3488 2461
rect 3574 2423 3589 2579
rect 3628 2537 3656 2593
tri 3748 2575 3766 2593 ne
rect 3766 2573 3788 2593
tri 3788 2573 3808 2593 sw
tri 3824 2579 3842 2597 ne
rect 3647 2503 3656 2537
rect 3690 2564 3732 2565
rect 3690 2530 3695 2564
rect 3725 2530 3732 2564
rect 3690 2521 3732 2530
rect 3766 2564 3808 2573
rect 3766 2530 3773 2564
rect 3803 2530 3808 2564
rect 3766 2525 3808 2530
rect 3842 2537 3870 2597
tri 3915 2584 3937 2606 se
rect 3937 2599 3952 2607
tri 3937 2584 3952 2599 nw
tri 3909 2578 3915 2584 se
rect 3915 2578 3924 2584
rect 3628 2493 3656 2503
tri 3656 2493 3680 2517 sw
rect 3628 2461 3670 2493
tri 3687 2485 3688 2486 sw
rect 3687 2461 3688 2485
tri 3690 2484 3727 2521 ne
rect 3727 2493 3732 2521
tri 3732 2493 3758 2519 sw
rect 3842 2503 3851 2537
rect 3842 2493 3870 2503
rect 3727 2484 3811 2493
tri 3727 2465 3746 2484 ne
rect 3746 2465 3811 2484
rect 3628 2439 3688 2461
rect 3810 2461 3811 2465
rect 3828 2461 3870 2493
rect 3810 2439 3870 2461
rect 3716 2423 3733 2437
rect 3765 2423 3782 2437
tri 3553 2387 3575 2409 se
rect 3575 2402 3590 2423
tri 3575 2387 3590 2402 nw
rect 3909 2402 3924 2578
tri 3924 2571 3937 2584 nw
rect 4010 2503 4025 2731
tri 3547 2381 3553 2387 se
rect 3553 2381 3562 2387
rect 3547 2365 3562 2381
tri 3562 2374 3575 2387 nw
rect 3716 2379 3733 2393
rect 3765 2379 3782 2393
tri 3909 2387 3924 2402 ne
tri 3924 2387 3946 2409 sw
rect 3547 2329 3562 2337
rect 3628 2365 3688 2379
rect 3643 2355 3688 2365
rect 3643 2337 3671 2355
tri 3547 2314 3562 2329 ne
tri 3562 2314 3584 2336 sw
rect 3628 2327 3671 2337
rect 3686 2351 3688 2355
rect 3810 2365 3870 2379
tri 3924 2374 3937 2387 ne
rect 3937 2381 3946 2387
tri 3946 2381 3952 2387 sw
rect 3810 2355 3855 2365
rect 3686 2327 3760 2351
rect 3628 2323 3760 2327
tri 3760 2323 3788 2351 sw
rect 3810 2341 3812 2355
tri 3810 2339 3812 2341 ne
rect 3824 2337 3855 2355
rect 3824 2327 3870 2337
rect 3937 2366 3952 2381
tri 3562 2302 3574 2314 ne
rect 3574 2309 3584 2314
tri 3584 2309 3589 2314 sw
rect 3473 1963 3488 2191
rect 3574 2201 3589 2309
rect 3628 2267 3656 2323
tri 3748 2305 3766 2323 ne
rect 3766 2303 3788 2323
tri 3788 2303 3808 2323 sw
tri 3824 2309 3842 2327 ne
rect 3647 2233 3656 2267
rect 3690 2294 3732 2295
rect 3690 2260 3695 2294
rect 3725 2260 3732 2294
rect 3690 2251 3732 2260
rect 3766 2294 3808 2303
rect 3766 2260 3773 2294
rect 3803 2260 3808 2294
rect 3766 2255 3808 2260
rect 3842 2267 3870 2327
tri 3915 2314 3937 2336 se
rect 3937 2329 3952 2337
tri 3937 2314 3952 2329 nw
tri 3909 2308 3915 2314 se
rect 3915 2308 3924 2314
rect 3628 2223 3656 2233
tri 3656 2223 3680 2247 sw
rect 3574 2153 3590 2201
rect 3628 2191 3670 2223
tri 3687 2215 3688 2216 sw
rect 3687 2191 3688 2215
tri 3690 2214 3727 2251 ne
rect 3727 2223 3732 2251
tri 3732 2223 3758 2249 sw
rect 3842 2233 3851 2267
rect 3842 2223 3870 2233
rect 3727 2214 3811 2223
tri 3727 2195 3746 2214 ne
rect 3746 2195 3811 2214
rect 3628 2169 3688 2191
rect 3810 2191 3811 2195
rect 3828 2191 3870 2223
rect 3810 2169 3870 2191
rect 3716 2153 3733 2167
rect 3765 2153 3782 2167
tri 3553 2117 3575 2139 se
rect 3575 2132 3590 2153
tri 3575 2117 3590 2132 nw
rect 3909 2132 3924 2308
tri 3924 2301 3937 2314 nw
rect 4010 2233 4025 2461
tri 3547 2111 3553 2117 se
rect 3553 2111 3562 2117
rect 3547 2095 3562 2111
tri 3562 2104 3575 2117 nw
rect 3716 2109 3733 2123
rect 3765 2109 3782 2123
tri 3909 2117 3924 2132 ne
tri 3924 2117 3946 2139 sw
rect 3547 2059 3562 2067
rect 3628 2095 3688 2109
rect 3643 2085 3688 2095
rect 3643 2067 3671 2085
tri 3547 2044 3562 2059 ne
tri 3562 2044 3584 2066 sw
rect 3628 2057 3671 2067
rect 3686 2081 3688 2085
rect 3810 2095 3870 2109
tri 3924 2104 3937 2117 ne
rect 3937 2111 3946 2117
tri 3946 2111 3952 2117 sw
rect 3810 2085 3855 2095
rect 3686 2057 3760 2081
rect 3628 2053 3760 2057
tri 3760 2053 3788 2081 sw
rect 3810 2071 3812 2085
tri 3810 2069 3812 2071 ne
rect 3824 2067 3855 2085
rect 3824 2057 3870 2067
rect 3937 2096 3952 2111
tri 3562 2032 3574 2044 ne
rect 3574 2039 3584 2044
tri 3584 2039 3589 2044 sw
rect 3473 1693 3488 1921
rect 3574 1883 3589 2039
rect 3628 1997 3656 2053
tri 3748 2035 3766 2053 ne
rect 3766 2033 3788 2053
tri 3788 2033 3808 2053 sw
tri 3824 2039 3842 2057 ne
rect 3647 1963 3656 1997
rect 3690 2024 3732 2025
rect 3690 1990 3695 2024
rect 3725 1990 3732 2024
rect 3690 1981 3732 1990
rect 3766 2024 3808 2033
rect 3766 1990 3773 2024
rect 3803 1990 3808 2024
rect 3766 1985 3808 1990
rect 3842 1997 3870 2057
tri 3915 2044 3937 2066 se
rect 3937 2059 3952 2067
tri 3937 2044 3952 2059 nw
tri 3909 2038 3915 2044 se
rect 3915 2038 3924 2044
rect 3628 1953 3656 1963
tri 3656 1953 3680 1977 sw
rect 3628 1921 3670 1953
tri 3687 1945 3688 1946 sw
rect 3687 1921 3688 1945
tri 3690 1944 3727 1981 ne
rect 3727 1953 3732 1981
tri 3732 1953 3758 1979 sw
rect 3842 1963 3851 1997
rect 3842 1953 3870 1963
rect 3727 1944 3811 1953
tri 3727 1925 3746 1944 ne
rect 3746 1925 3811 1944
rect 3628 1899 3688 1921
rect 3810 1921 3811 1925
rect 3828 1921 3870 1953
rect 3810 1899 3870 1921
rect 3716 1883 3733 1897
rect 3765 1883 3782 1897
tri 3553 1847 3575 1869 se
rect 3575 1862 3590 1883
tri 3575 1847 3590 1862 nw
rect 3909 1862 3924 2038
tri 3924 2031 3937 2044 nw
rect 4010 1963 4025 2191
tri 3547 1841 3553 1847 se
rect 3553 1841 3562 1847
rect 3547 1825 3562 1841
tri 3562 1834 3575 1847 nw
rect 3716 1839 3733 1853
rect 3765 1839 3782 1853
tri 3909 1847 3924 1862 ne
tri 3924 1847 3946 1869 sw
rect 3547 1789 3562 1797
rect 3628 1825 3688 1839
rect 3643 1815 3688 1825
rect 3643 1797 3671 1815
tri 3547 1774 3562 1789 ne
tri 3562 1774 3584 1796 sw
rect 3628 1787 3671 1797
rect 3686 1811 3688 1815
rect 3810 1825 3870 1839
tri 3924 1834 3937 1847 ne
rect 3937 1841 3946 1847
tri 3946 1841 3952 1847 sw
rect 3810 1815 3855 1825
rect 3686 1787 3760 1811
rect 3628 1783 3760 1787
tri 3760 1783 3788 1811 sw
rect 3810 1801 3812 1815
tri 3810 1799 3812 1801 ne
rect 3824 1797 3855 1815
rect 3824 1787 3870 1797
rect 3937 1826 3952 1841
tri 3562 1762 3574 1774 ne
rect 3574 1769 3584 1774
tri 3584 1769 3589 1774 sw
rect 3473 1423 3488 1651
rect 3574 1661 3589 1769
rect 3628 1727 3656 1783
tri 3748 1765 3766 1783 ne
rect 3766 1763 3788 1783
tri 3788 1763 3808 1783 sw
tri 3824 1769 3842 1787 ne
rect 3647 1693 3656 1727
rect 3690 1754 3732 1755
rect 3690 1720 3695 1754
rect 3725 1720 3732 1754
rect 3690 1711 3732 1720
rect 3766 1754 3808 1763
rect 3766 1720 3773 1754
rect 3803 1720 3808 1754
rect 3766 1715 3808 1720
rect 3842 1727 3870 1787
tri 3915 1774 3937 1796 se
rect 3937 1789 3952 1797
tri 3937 1774 3952 1789 nw
tri 3909 1768 3915 1774 se
rect 3915 1768 3924 1774
rect 3628 1683 3656 1693
tri 3656 1683 3680 1707 sw
rect 3574 1613 3590 1661
rect 3628 1651 3670 1683
tri 3687 1675 3688 1676 sw
rect 3687 1651 3688 1675
tri 3690 1674 3727 1711 ne
rect 3727 1683 3732 1711
tri 3732 1683 3758 1709 sw
rect 3842 1693 3851 1727
rect 3842 1683 3870 1693
rect 3727 1674 3811 1683
tri 3727 1655 3746 1674 ne
rect 3746 1655 3811 1674
rect 3628 1629 3688 1651
rect 3810 1651 3811 1655
rect 3828 1651 3870 1683
rect 3810 1629 3870 1651
rect 3716 1613 3733 1627
rect 3765 1613 3782 1627
tri 3553 1577 3575 1599 se
rect 3575 1592 3590 1613
tri 3575 1577 3590 1592 nw
rect 3909 1592 3924 1768
tri 3924 1761 3937 1774 nw
rect 4010 1693 4025 1921
tri 3547 1571 3553 1577 se
rect 3553 1571 3562 1577
rect 3547 1555 3562 1571
tri 3562 1564 3575 1577 nw
rect 3716 1569 3733 1583
rect 3765 1569 3782 1583
tri 3909 1577 3924 1592 ne
tri 3924 1577 3946 1599 sw
rect 3547 1519 3562 1527
rect 3628 1555 3688 1569
rect 3643 1545 3688 1555
rect 3643 1527 3671 1545
tri 3547 1504 3562 1519 ne
tri 3562 1504 3584 1526 sw
rect 3628 1517 3671 1527
rect 3686 1541 3688 1545
rect 3810 1555 3870 1569
tri 3924 1564 3937 1577 ne
rect 3937 1571 3946 1577
tri 3946 1571 3952 1577 sw
rect 3810 1545 3855 1555
rect 3686 1517 3760 1541
rect 3628 1513 3760 1517
tri 3760 1513 3788 1541 sw
rect 3810 1531 3812 1545
tri 3810 1529 3812 1531 ne
rect 3824 1527 3855 1545
rect 3824 1517 3870 1527
rect 3937 1556 3952 1571
tri 3562 1492 3574 1504 ne
rect 3574 1499 3584 1504
tri 3584 1499 3589 1504 sw
rect 3473 1153 3488 1381
rect 3574 1343 3589 1499
rect 3628 1457 3656 1513
tri 3748 1495 3766 1513 ne
rect 3766 1493 3788 1513
tri 3788 1493 3808 1513 sw
tri 3824 1499 3842 1517 ne
rect 3647 1423 3656 1457
rect 3690 1484 3732 1485
rect 3690 1450 3695 1484
rect 3725 1450 3732 1484
rect 3690 1441 3732 1450
rect 3766 1484 3808 1493
rect 3766 1450 3773 1484
rect 3803 1450 3808 1484
rect 3766 1445 3808 1450
rect 3842 1457 3870 1517
tri 3915 1504 3937 1526 se
rect 3937 1519 3952 1527
tri 3937 1504 3952 1519 nw
tri 3909 1498 3915 1504 se
rect 3915 1498 3924 1504
rect 3628 1413 3656 1423
tri 3656 1413 3680 1437 sw
rect 3628 1381 3670 1413
tri 3687 1405 3688 1406 sw
rect 3687 1381 3688 1405
tri 3690 1404 3727 1441 ne
rect 3727 1413 3732 1441
tri 3732 1413 3758 1439 sw
rect 3842 1423 3851 1457
rect 3842 1413 3870 1423
rect 3727 1404 3811 1413
tri 3727 1385 3746 1404 ne
rect 3746 1385 3811 1404
rect 3628 1359 3688 1381
rect 3810 1381 3811 1385
rect 3828 1381 3870 1413
rect 3810 1359 3870 1381
rect 3716 1343 3733 1357
rect 3765 1343 3782 1357
tri 3553 1307 3575 1329 se
rect 3575 1322 3590 1343
tri 3575 1307 3590 1322 nw
rect 3909 1322 3924 1498
tri 3924 1491 3937 1504 nw
rect 4010 1423 4025 1651
tri 3547 1301 3553 1307 se
rect 3553 1301 3562 1307
rect 3547 1285 3562 1301
tri 3562 1294 3575 1307 nw
rect 3716 1299 3733 1313
rect 3765 1299 3782 1313
tri 3909 1307 3924 1322 ne
tri 3924 1307 3946 1329 sw
rect 3547 1249 3562 1257
rect 3628 1285 3688 1299
rect 3643 1275 3688 1285
rect 3643 1257 3671 1275
tri 3547 1234 3562 1249 ne
tri 3562 1234 3584 1256 sw
rect 3628 1247 3671 1257
rect 3686 1271 3688 1275
rect 3810 1285 3870 1299
tri 3924 1294 3937 1307 ne
rect 3937 1301 3946 1307
tri 3946 1301 3952 1307 sw
rect 3810 1275 3855 1285
rect 3686 1247 3760 1271
rect 3628 1243 3760 1247
tri 3760 1243 3788 1271 sw
rect 3810 1261 3812 1275
tri 3810 1259 3812 1261 ne
rect 3824 1257 3855 1275
rect 3824 1247 3870 1257
rect 3937 1286 3952 1301
tri 3562 1222 3574 1234 ne
rect 3574 1229 3584 1234
tri 3584 1229 3589 1234 sw
rect 3473 883 3488 1111
rect 3574 1121 3589 1229
rect 3628 1187 3656 1243
tri 3748 1225 3766 1243 ne
rect 3766 1223 3788 1243
tri 3788 1223 3808 1243 sw
tri 3824 1229 3842 1247 ne
rect 3647 1153 3656 1187
rect 3690 1214 3732 1215
rect 3690 1180 3695 1214
rect 3725 1180 3732 1214
rect 3690 1171 3732 1180
rect 3766 1214 3808 1223
rect 3766 1180 3773 1214
rect 3803 1180 3808 1214
rect 3766 1175 3808 1180
rect 3842 1187 3870 1247
tri 3915 1234 3937 1256 se
rect 3937 1249 3952 1257
tri 3937 1234 3952 1249 nw
tri 3909 1228 3915 1234 se
rect 3915 1228 3924 1234
rect 3628 1143 3656 1153
tri 3656 1143 3680 1167 sw
rect 3574 1073 3590 1121
rect 3628 1111 3670 1143
tri 3687 1135 3688 1136 sw
rect 3687 1111 3688 1135
tri 3690 1134 3727 1171 ne
rect 3727 1143 3732 1171
tri 3732 1143 3758 1169 sw
rect 3842 1153 3851 1187
rect 3842 1143 3870 1153
rect 3727 1134 3811 1143
tri 3727 1115 3746 1134 ne
rect 3746 1115 3811 1134
rect 3628 1089 3688 1111
rect 3810 1111 3811 1115
rect 3828 1111 3870 1143
rect 3810 1089 3870 1111
rect 3716 1073 3733 1087
rect 3765 1073 3782 1087
tri 3553 1037 3575 1059 se
rect 3575 1052 3590 1073
tri 3575 1037 3590 1052 nw
rect 3909 1052 3924 1228
tri 3924 1221 3937 1234 nw
rect 4010 1153 4025 1381
tri 3547 1031 3553 1037 se
rect 3553 1031 3562 1037
rect 3547 1015 3562 1031
tri 3562 1024 3575 1037 nw
rect 3716 1029 3733 1043
rect 3765 1029 3782 1043
tri 3909 1037 3924 1052 ne
tri 3924 1037 3946 1059 sw
rect 3547 979 3562 987
rect 3628 1015 3688 1029
rect 3643 1005 3688 1015
rect 3643 987 3671 1005
tri 3547 964 3562 979 ne
tri 3562 964 3584 986 sw
rect 3628 977 3671 987
rect 3686 1001 3688 1005
rect 3810 1015 3870 1029
tri 3924 1024 3937 1037 ne
rect 3937 1031 3946 1037
tri 3946 1031 3952 1037 sw
rect 3810 1005 3855 1015
rect 3686 977 3760 1001
rect 3628 973 3760 977
tri 3760 973 3788 1001 sw
rect 3810 991 3812 1005
tri 3810 989 3812 991 ne
rect 3824 987 3855 1005
rect 3824 977 3870 987
rect 3937 1016 3952 1031
tri 3562 952 3574 964 ne
rect 3574 959 3584 964
tri 3584 959 3589 964 sw
rect 3473 613 3488 841
rect 3574 803 3589 959
rect 3628 917 3656 973
tri 3748 955 3766 973 ne
rect 3766 953 3788 973
tri 3788 953 3808 973 sw
tri 3824 959 3842 977 ne
rect 3647 883 3656 917
rect 3690 944 3732 945
rect 3690 910 3695 944
rect 3725 910 3732 944
rect 3690 901 3732 910
rect 3766 944 3808 953
rect 3766 910 3773 944
rect 3803 910 3808 944
rect 3766 905 3808 910
rect 3842 917 3870 977
tri 3915 964 3937 986 se
rect 3937 979 3952 987
tri 3937 964 3952 979 nw
tri 3909 958 3915 964 se
rect 3915 958 3924 964
rect 3628 873 3656 883
tri 3656 873 3680 897 sw
rect 3628 841 3670 873
tri 3687 865 3688 866 sw
rect 3687 841 3688 865
tri 3690 864 3727 901 ne
rect 3727 873 3732 901
tri 3732 873 3758 899 sw
rect 3842 883 3851 917
rect 3842 873 3870 883
rect 3727 864 3811 873
tri 3727 845 3746 864 ne
rect 3746 845 3811 864
rect 3628 819 3688 841
rect 3810 841 3811 845
rect 3828 841 3870 873
rect 3810 819 3870 841
rect 3716 803 3733 817
rect 3765 803 3782 817
tri 3553 767 3575 789 se
rect 3575 782 3590 803
tri 3575 767 3590 782 nw
rect 3909 782 3924 958
tri 3924 951 3937 964 nw
rect 4010 883 4025 1111
tri 3547 761 3553 767 se
rect 3553 761 3562 767
rect 3547 745 3562 761
tri 3562 754 3575 767 nw
rect 3716 759 3733 773
rect 3765 759 3782 773
tri 3909 767 3924 782 ne
tri 3924 767 3946 789 sw
rect 3547 709 3562 717
rect 3628 745 3688 759
rect 3643 735 3688 745
rect 3643 717 3671 735
tri 3547 694 3562 709 ne
tri 3562 694 3584 716 sw
rect 3628 707 3671 717
rect 3686 731 3688 735
rect 3810 745 3870 759
tri 3924 754 3937 767 ne
rect 3937 761 3946 767
tri 3946 761 3952 767 sw
rect 3810 735 3855 745
rect 3686 707 3760 731
rect 3628 703 3760 707
tri 3760 703 3788 731 sw
rect 3810 721 3812 735
tri 3810 719 3812 721 ne
rect 3824 717 3855 735
rect 3824 707 3870 717
rect 3937 746 3952 761
tri 3562 682 3574 694 ne
rect 3574 689 3584 694
tri 3584 689 3589 694 sw
rect 3473 343 3488 571
rect 3574 581 3589 689
rect 3628 647 3656 703
tri 3748 685 3766 703 ne
rect 3766 683 3788 703
tri 3788 683 3808 703 sw
tri 3824 689 3842 707 ne
rect 3647 613 3656 647
rect 3690 674 3732 675
rect 3690 640 3695 674
rect 3725 640 3732 674
rect 3690 631 3732 640
rect 3766 674 3808 683
rect 3766 640 3773 674
rect 3803 640 3808 674
rect 3766 635 3808 640
rect 3842 647 3870 707
tri 3915 694 3937 716 se
rect 3937 709 3952 717
tri 3937 694 3952 709 nw
tri 3909 688 3915 694 se
rect 3915 688 3924 694
rect 3628 603 3656 613
tri 3656 603 3680 627 sw
rect 3574 533 3590 581
rect 3628 571 3670 603
tri 3687 595 3688 596 sw
rect 3687 571 3688 595
tri 3690 594 3727 631 ne
rect 3727 603 3732 631
tri 3732 603 3758 629 sw
rect 3842 613 3851 647
rect 3842 603 3870 613
rect 3727 594 3811 603
tri 3727 575 3746 594 ne
rect 3746 575 3811 594
rect 3628 549 3688 571
rect 3810 571 3811 575
rect 3828 571 3870 603
rect 3810 549 3870 571
rect 3716 533 3733 547
rect 3765 533 3782 547
tri 3553 497 3575 519 se
rect 3575 512 3590 533
tri 3575 497 3590 512 nw
rect 3909 512 3924 688
tri 3924 681 3937 694 nw
rect 4010 613 4025 841
tri 3547 491 3553 497 se
rect 3553 491 3562 497
rect 3547 475 3562 491
tri 3562 484 3575 497 nw
rect 3716 489 3733 503
rect 3765 489 3782 503
tri 3909 497 3924 512 ne
tri 3924 497 3946 519 sw
rect 3547 439 3562 447
rect 3628 475 3688 489
rect 3643 465 3688 475
rect 3643 447 3671 465
tri 3547 424 3562 439 ne
tri 3562 424 3584 446 sw
rect 3628 437 3671 447
rect 3686 461 3688 465
rect 3810 475 3870 489
tri 3924 484 3937 497 ne
rect 3937 491 3946 497
tri 3946 491 3952 497 sw
rect 3810 465 3855 475
rect 3686 437 3760 461
rect 3628 433 3760 437
tri 3760 433 3788 461 sw
rect 3810 451 3812 465
tri 3810 449 3812 451 ne
rect 3824 447 3855 465
rect 3824 437 3870 447
rect 3937 476 3952 491
tri 3562 412 3574 424 ne
rect 3574 419 3584 424
tri 3584 419 3589 424 sw
rect 3473 73 3488 301
rect 3574 263 3589 419
rect 3628 377 3656 433
tri 3748 415 3766 433 ne
rect 3766 413 3788 433
tri 3788 413 3808 433 sw
tri 3824 419 3842 437 ne
rect 3647 343 3656 377
rect 3690 404 3732 405
rect 3690 370 3695 404
rect 3725 370 3732 404
rect 3690 361 3732 370
rect 3766 404 3808 413
rect 3766 370 3773 404
rect 3803 370 3808 404
rect 3766 365 3808 370
rect 3842 377 3870 437
tri 3915 424 3937 446 se
rect 3937 439 3952 447
tri 3937 424 3952 439 nw
tri 3909 418 3915 424 se
rect 3915 418 3924 424
rect 3628 333 3656 343
tri 3656 333 3680 357 sw
rect 3628 301 3670 333
tri 3687 325 3688 326 sw
rect 3687 301 3688 325
tri 3690 324 3727 361 ne
rect 3727 333 3732 361
tri 3732 333 3758 359 sw
rect 3842 343 3851 377
rect 3842 333 3870 343
rect 3727 324 3811 333
tri 3727 305 3746 324 ne
rect 3746 305 3811 324
rect 3628 279 3688 301
rect 3810 301 3811 305
rect 3828 301 3870 333
rect 3810 279 3870 301
rect 3716 263 3733 277
rect 3765 263 3782 277
tri 3553 227 3575 249 se
rect 3575 242 3590 263
tri 3575 227 3590 242 nw
rect 3909 242 3924 418
tri 3924 411 3937 424 nw
rect 4010 343 4025 571
tri 3547 221 3553 227 se
rect 3553 221 3562 227
rect 3547 205 3562 221
tri 3562 214 3575 227 nw
rect 3716 219 3733 233
rect 3765 219 3782 233
tri 3909 227 3924 242 ne
tri 3924 227 3946 249 sw
rect 3547 169 3562 177
rect 3628 205 3688 219
rect 3643 195 3688 205
rect 3643 177 3671 195
tri 3547 154 3562 169 ne
tri 3562 154 3584 176 sw
rect 3628 167 3671 177
rect 3686 191 3688 195
rect 3810 205 3870 219
tri 3924 214 3937 227 ne
rect 3937 221 3946 227
tri 3946 221 3952 227 sw
rect 3810 195 3855 205
rect 3686 167 3760 191
rect 3628 163 3760 167
tri 3760 163 3788 191 sw
rect 3810 181 3812 195
tri 3810 179 3812 181 ne
rect 3824 177 3855 195
rect 3824 167 3870 177
rect 3937 206 3952 221
tri 3562 142 3574 154 ne
rect 3574 149 3584 154
tri 3584 149 3589 154 sw
rect 3473 -55 3488 31
rect 3574 -55 3589 149
rect 3628 107 3656 163
tri 3748 145 3766 163 ne
rect 3766 143 3788 163
tri 3788 143 3808 163 sw
tri 3824 149 3842 167 ne
rect 3647 73 3656 107
rect 3690 134 3732 135
rect 3690 100 3695 134
rect 3725 100 3732 134
rect 3690 91 3732 100
rect 3766 134 3808 143
rect 3766 100 3773 134
rect 3803 100 3808 134
rect 3766 95 3808 100
rect 3842 107 3870 167
tri 3915 154 3937 176 se
rect 3937 169 3952 177
tri 3937 154 3952 169 nw
tri 3909 148 3915 154 se
rect 3915 148 3924 154
rect 3628 63 3656 73
tri 3656 63 3680 87 sw
rect 3628 31 3670 63
tri 3687 55 3688 56 sw
rect 3687 31 3688 55
tri 3690 54 3727 91 ne
rect 3727 63 3732 91
tri 3732 63 3758 89 sw
rect 3842 73 3851 107
rect 3842 63 3870 73
rect 3727 54 3811 63
tri 3727 35 3746 54 ne
rect 3746 35 3811 54
rect 3628 9 3688 31
rect 3810 31 3811 35
rect 3828 31 3870 63
rect 3810 9 3870 31
rect 3716 -7 3733 7
rect 3765 -7 3782 7
rect 3909 -55 3924 148
tri 3924 141 3937 154 nw
rect 4010 73 4025 301
rect 4010 -55 4025 31
rect 4053 4123 4068 4361
tri 4133 4277 4155 4299 se
rect 4155 4292 4170 4361
tri 4155 4277 4170 4292 nw
rect 4489 4292 4504 4361
tri 4127 4271 4133 4277 se
rect 4133 4271 4142 4277
rect 4127 4255 4142 4271
tri 4142 4264 4155 4277 nw
rect 4296 4269 4313 4283
rect 4345 4269 4362 4283
tri 4489 4277 4504 4292 ne
tri 4504 4277 4526 4299 sw
rect 4127 4219 4142 4227
rect 4208 4255 4268 4269
rect 4223 4245 4268 4255
rect 4223 4227 4251 4245
tri 4127 4204 4142 4219 ne
tri 4142 4204 4164 4226 sw
rect 4208 4217 4251 4227
rect 4266 4241 4268 4245
rect 4390 4255 4450 4269
tri 4504 4264 4517 4277 ne
rect 4517 4271 4526 4277
tri 4526 4271 4532 4277 sw
rect 4390 4245 4435 4255
rect 4266 4217 4340 4241
rect 4208 4213 4340 4217
tri 4340 4213 4368 4241 sw
rect 4390 4231 4392 4245
tri 4390 4229 4392 4231 ne
rect 4404 4227 4435 4245
rect 4404 4217 4450 4227
rect 4517 4256 4532 4271
tri 4142 4192 4154 4204 ne
rect 4154 4199 4164 4204
tri 4164 4199 4169 4204 sw
rect 4053 3853 4068 4081
rect 4154 4043 4169 4199
rect 4208 4157 4236 4213
tri 4328 4195 4346 4213 ne
rect 4346 4193 4368 4213
tri 4368 4193 4388 4213 sw
tri 4404 4199 4422 4217 ne
rect 4227 4123 4236 4157
rect 4270 4184 4312 4185
rect 4270 4150 4275 4184
rect 4305 4150 4312 4184
rect 4270 4141 4312 4150
rect 4346 4184 4388 4193
rect 4346 4150 4353 4184
rect 4383 4150 4388 4184
rect 4346 4145 4388 4150
rect 4422 4157 4450 4217
tri 4495 4204 4517 4226 se
rect 4517 4219 4532 4227
tri 4517 4204 4532 4219 nw
tri 4489 4198 4495 4204 se
rect 4495 4198 4504 4204
rect 4208 4113 4236 4123
tri 4236 4113 4260 4137 sw
rect 4208 4081 4250 4113
tri 4267 4105 4268 4106 sw
rect 4267 4081 4268 4105
tri 4270 4104 4307 4141 ne
rect 4307 4113 4312 4141
tri 4312 4113 4338 4139 sw
rect 4422 4123 4431 4157
rect 4422 4113 4450 4123
rect 4307 4104 4391 4113
tri 4307 4085 4326 4104 ne
rect 4326 4085 4391 4104
rect 4208 4059 4268 4081
rect 4390 4081 4391 4085
rect 4408 4081 4450 4113
rect 4390 4059 4450 4081
rect 4296 4043 4313 4057
rect 4345 4043 4362 4057
tri 4133 4007 4155 4029 se
rect 4155 4022 4170 4043
tri 4155 4007 4170 4022 nw
rect 4489 4022 4504 4198
tri 4504 4191 4517 4204 nw
rect 4590 4123 4605 4361
tri 4127 4001 4133 4007 se
rect 4133 4001 4142 4007
rect 4127 3985 4142 4001
tri 4142 3994 4155 4007 nw
rect 4296 3999 4313 4013
rect 4345 3999 4362 4013
tri 4489 4007 4504 4022 ne
tri 4504 4007 4526 4029 sw
rect 4127 3949 4142 3957
rect 4208 3985 4268 3999
rect 4223 3975 4268 3985
rect 4223 3957 4251 3975
tri 4127 3934 4142 3949 ne
tri 4142 3934 4164 3956 sw
rect 4208 3947 4251 3957
rect 4266 3971 4268 3975
rect 4390 3985 4450 3999
tri 4504 3994 4517 4007 ne
rect 4517 4001 4526 4007
tri 4526 4001 4532 4007 sw
rect 4390 3975 4435 3985
rect 4266 3947 4340 3971
rect 4208 3943 4340 3947
tri 4340 3943 4368 3971 sw
rect 4390 3961 4392 3975
tri 4390 3959 4392 3961 ne
rect 4404 3957 4435 3975
rect 4404 3947 4450 3957
rect 4517 3986 4532 4001
tri 4142 3922 4154 3934 ne
rect 4154 3929 4164 3934
tri 4164 3929 4169 3934 sw
rect 4053 3583 4068 3811
rect 4154 3821 4169 3929
rect 4208 3887 4236 3943
tri 4328 3925 4346 3943 ne
rect 4346 3923 4368 3943
tri 4368 3923 4388 3943 sw
tri 4404 3929 4422 3947 ne
rect 4227 3853 4236 3887
rect 4270 3914 4312 3915
rect 4270 3880 4275 3914
rect 4305 3880 4312 3914
rect 4270 3871 4312 3880
rect 4346 3914 4388 3923
rect 4346 3880 4353 3914
rect 4383 3880 4388 3914
rect 4346 3875 4388 3880
rect 4422 3887 4450 3947
tri 4495 3934 4517 3956 se
rect 4517 3949 4532 3957
tri 4517 3934 4532 3949 nw
tri 4489 3928 4495 3934 se
rect 4495 3928 4504 3934
rect 4208 3843 4236 3853
tri 4236 3843 4260 3867 sw
rect 4154 3773 4170 3821
rect 4208 3811 4250 3843
tri 4267 3835 4268 3836 sw
rect 4267 3811 4268 3835
tri 4270 3834 4307 3871 ne
rect 4307 3843 4312 3871
tri 4312 3843 4338 3869 sw
rect 4422 3853 4431 3887
rect 4422 3843 4450 3853
rect 4307 3834 4391 3843
tri 4307 3815 4326 3834 ne
rect 4326 3815 4391 3834
rect 4208 3789 4268 3811
rect 4390 3811 4391 3815
rect 4408 3811 4450 3843
rect 4390 3789 4450 3811
rect 4296 3773 4313 3787
rect 4345 3773 4362 3787
tri 4133 3737 4155 3759 se
rect 4155 3752 4170 3773
tri 4155 3737 4170 3752 nw
rect 4489 3752 4504 3928
tri 4504 3921 4517 3934 nw
rect 4590 3853 4605 4081
tri 4127 3731 4133 3737 se
rect 4133 3731 4142 3737
rect 4127 3715 4142 3731
tri 4142 3724 4155 3737 nw
rect 4296 3729 4313 3743
rect 4345 3729 4362 3743
tri 4489 3737 4504 3752 ne
tri 4504 3737 4526 3759 sw
rect 4127 3679 4142 3687
rect 4208 3715 4268 3729
rect 4223 3705 4268 3715
rect 4223 3687 4251 3705
tri 4127 3664 4142 3679 ne
tri 4142 3664 4164 3686 sw
rect 4208 3677 4251 3687
rect 4266 3701 4268 3705
rect 4390 3715 4450 3729
tri 4504 3724 4517 3737 ne
rect 4517 3731 4526 3737
tri 4526 3731 4532 3737 sw
rect 4390 3705 4435 3715
rect 4266 3677 4340 3701
rect 4208 3673 4340 3677
tri 4340 3673 4368 3701 sw
rect 4390 3691 4392 3705
tri 4390 3689 4392 3691 ne
rect 4404 3687 4435 3705
rect 4404 3677 4450 3687
rect 4517 3716 4532 3731
tri 4142 3652 4154 3664 ne
rect 4154 3659 4164 3664
tri 4164 3659 4169 3664 sw
rect 4053 3313 4068 3541
rect 4154 3503 4169 3659
rect 4208 3617 4236 3673
tri 4328 3655 4346 3673 ne
rect 4346 3653 4368 3673
tri 4368 3653 4388 3673 sw
tri 4404 3659 4422 3677 ne
rect 4227 3583 4236 3617
rect 4270 3644 4312 3645
rect 4270 3610 4275 3644
rect 4305 3610 4312 3644
rect 4270 3601 4312 3610
rect 4346 3644 4388 3653
rect 4346 3610 4353 3644
rect 4383 3610 4388 3644
rect 4346 3605 4388 3610
rect 4422 3617 4450 3677
tri 4495 3664 4517 3686 se
rect 4517 3679 4532 3687
tri 4517 3664 4532 3679 nw
tri 4489 3658 4495 3664 se
rect 4495 3658 4504 3664
rect 4208 3573 4236 3583
tri 4236 3573 4260 3597 sw
rect 4208 3541 4250 3573
tri 4267 3565 4268 3566 sw
rect 4267 3541 4268 3565
tri 4270 3564 4307 3601 ne
rect 4307 3573 4312 3601
tri 4312 3573 4338 3599 sw
rect 4422 3583 4431 3617
rect 4422 3573 4450 3583
rect 4307 3564 4391 3573
tri 4307 3545 4326 3564 ne
rect 4326 3545 4391 3564
rect 4208 3519 4268 3541
rect 4390 3541 4391 3545
rect 4408 3541 4450 3573
rect 4390 3519 4450 3541
rect 4296 3503 4313 3517
rect 4345 3503 4362 3517
tri 4133 3467 4155 3489 se
rect 4155 3482 4170 3503
tri 4155 3467 4170 3482 nw
rect 4489 3482 4504 3658
tri 4504 3651 4517 3664 nw
rect 4590 3583 4605 3811
tri 4127 3461 4133 3467 se
rect 4133 3461 4142 3467
rect 4127 3445 4142 3461
tri 4142 3454 4155 3467 nw
rect 4296 3459 4313 3473
rect 4345 3459 4362 3473
tri 4489 3467 4504 3482 ne
tri 4504 3467 4526 3489 sw
rect 4127 3409 4142 3417
rect 4208 3445 4268 3459
rect 4223 3435 4268 3445
rect 4223 3417 4251 3435
tri 4127 3394 4142 3409 ne
tri 4142 3394 4164 3416 sw
rect 4208 3407 4251 3417
rect 4266 3431 4268 3435
rect 4390 3445 4450 3459
tri 4504 3454 4517 3467 ne
rect 4517 3461 4526 3467
tri 4526 3461 4532 3467 sw
rect 4390 3435 4435 3445
rect 4266 3407 4340 3431
rect 4208 3403 4340 3407
tri 4340 3403 4368 3431 sw
rect 4390 3421 4392 3435
tri 4390 3419 4392 3421 ne
rect 4404 3417 4435 3435
rect 4404 3407 4450 3417
rect 4517 3446 4532 3461
tri 4142 3382 4154 3394 ne
rect 4154 3389 4164 3394
tri 4164 3389 4169 3394 sw
rect 4053 3043 4068 3271
rect 4154 3281 4169 3389
rect 4208 3347 4236 3403
tri 4328 3385 4346 3403 ne
rect 4346 3383 4368 3403
tri 4368 3383 4388 3403 sw
tri 4404 3389 4422 3407 ne
rect 4227 3313 4236 3347
rect 4270 3374 4312 3375
rect 4270 3340 4275 3374
rect 4305 3340 4312 3374
rect 4270 3331 4312 3340
rect 4346 3374 4388 3383
rect 4346 3340 4353 3374
rect 4383 3340 4388 3374
rect 4346 3335 4388 3340
rect 4422 3347 4450 3407
tri 4495 3394 4517 3416 se
rect 4517 3409 4532 3417
tri 4517 3394 4532 3409 nw
tri 4489 3388 4495 3394 se
rect 4495 3388 4504 3394
rect 4208 3303 4236 3313
tri 4236 3303 4260 3327 sw
rect 4154 3233 4170 3281
rect 4208 3271 4250 3303
tri 4267 3295 4268 3296 sw
rect 4267 3271 4268 3295
tri 4270 3294 4307 3331 ne
rect 4307 3303 4312 3331
tri 4312 3303 4338 3329 sw
rect 4422 3313 4431 3347
rect 4422 3303 4450 3313
rect 4307 3294 4391 3303
tri 4307 3275 4326 3294 ne
rect 4326 3275 4391 3294
rect 4208 3249 4268 3271
rect 4390 3271 4391 3275
rect 4408 3271 4450 3303
rect 4390 3249 4450 3271
rect 4296 3233 4313 3247
rect 4345 3233 4362 3247
tri 4133 3197 4155 3219 se
rect 4155 3212 4170 3233
tri 4155 3197 4170 3212 nw
rect 4489 3212 4504 3388
tri 4504 3381 4517 3394 nw
rect 4590 3313 4605 3541
tri 4127 3191 4133 3197 se
rect 4133 3191 4142 3197
rect 4127 3175 4142 3191
tri 4142 3184 4155 3197 nw
rect 4296 3189 4313 3203
rect 4345 3189 4362 3203
tri 4489 3197 4504 3212 ne
tri 4504 3197 4526 3219 sw
rect 4127 3139 4142 3147
rect 4208 3175 4268 3189
rect 4223 3165 4268 3175
rect 4223 3147 4251 3165
tri 4127 3124 4142 3139 ne
tri 4142 3124 4164 3146 sw
rect 4208 3137 4251 3147
rect 4266 3161 4268 3165
rect 4390 3175 4450 3189
tri 4504 3184 4517 3197 ne
rect 4517 3191 4526 3197
tri 4526 3191 4532 3197 sw
rect 4390 3165 4435 3175
rect 4266 3137 4340 3161
rect 4208 3133 4340 3137
tri 4340 3133 4368 3161 sw
rect 4390 3151 4392 3165
tri 4390 3149 4392 3151 ne
rect 4404 3147 4435 3165
rect 4404 3137 4450 3147
rect 4517 3176 4532 3191
tri 4142 3112 4154 3124 ne
rect 4154 3119 4164 3124
tri 4164 3119 4169 3124 sw
rect 4053 2773 4068 3001
rect 4154 2963 4169 3119
rect 4208 3077 4236 3133
tri 4328 3115 4346 3133 ne
rect 4346 3113 4368 3133
tri 4368 3113 4388 3133 sw
tri 4404 3119 4422 3137 ne
rect 4227 3043 4236 3077
rect 4270 3104 4312 3105
rect 4270 3070 4275 3104
rect 4305 3070 4312 3104
rect 4270 3061 4312 3070
rect 4346 3104 4388 3113
rect 4346 3070 4353 3104
rect 4383 3070 4388 3104
rect 4346 3065 4388 3070
rect 4422 3077 4450 3137
tri 4495 3124 4517 3146 se
rect 4517 3139 4532 3147
tri 4517 3124 4532 3139 nw
tri 4489 3118 4495 3124 se
rect 4495 3118 4504 3124
rect 4208 3033 4236 3043
tri 4236 3033 4260 3057 sw
rect 4208 3001 4250 3033
tri 4267 3025 4268 3026 sw
rect 4267 3001 4268 3025
tri 4270 3024 4307 3061 ne
rect 4307 3033 4312 3061
tri 4312 3033 4338 3059 sw
rect 4422 3043 4431 3077
rect 4422 3033 4450 3043
rect 4307 3024 4391 3033
tri 4307 3005 4326 3024 ne
rect 4326 3005 4391 3024
rect 4208 2979 4268 3001
rect 4390 3001 4391 3005
rect 4408 3001 4450 3033
rect 4390 2979 4450 3001
rect 4296 2963 4313 2977
rect 4345 2963 4362 2977
tri 4133 2927 4155 2949 se
rect 4155 2942 4170 2963
tri 4155 2927 4170 2942 nw
rect 4489 2942 4504 3118
tri 4504 3111 4517 3124 nw
rect 4590 3043 4605 3271
tri 4127 2921 4133 2927 se
rect 4133 2921 4142 2927
rect 4127 2905 4142 2921
tri 4142 2914 4155 2927 nw
rect 4296 2919 4313 2933
rect 4345 2919 4362 2933
tri 4489 2927 4504 2942 ne
tri 4504 2927 4526 2949 sw
rect 4127 2869 4142 2877
rect 4208 2905 4268 2919
rect 4223 2895 4268 2905
rect 4223 2877 4251 2895
tri 4127 2854 4142 2869 ne
tri 4142 2854 4164 2876 sw
rect 4208 2867 4251 2877
rect 4266 2891 4268 2895
rect 4390 2905 4450 2919
tri 4504 2914 4517 2927 ne
rect 4517 2921 4526 2927
tri 4526 2921 4532 2927 sw
rect 4390 2895 4435 2905
rect 4266 2867 4340 2891
rect 4208 2863 4340 2867
tri 4340 2863 4368 2891 sw
rect 4390 2881 4392 2895
tri 4390 2879 4392 2881 ne
rect 4404 2877 4435 2895
rect 4404 2867 4450 2877
rect 4517 2906 4532 2921
tri 4142 2842 4154 2854 ne
rect 4154 2849 4164 2854
tri 4164 2849 4169 2854 sw
rect 4053 2503 4068 2731
rect 4154 2741 4169 2849
rect 4208 2807 4236 2863
tri 4328 2845 4346 2863 ne
rect 4346 2843 4368 2863
tri 4368 2843 4388 2863 sw
tri 4404 2849 4422 2867 ne
rect 4227 2773 4236 2807
rect 4270 2834 4312 2835
rect 4270 2800 4275 2834
rect 4305 2800 4312 2834
rect 4270 2791 4312 2800
rect 4346 2834 4388 2843
rect 4346 2800 4353 2834
rect 4383 2800 4388 2834
rect 4346 2795 4388 2800
rect 4422 2807 4450 2867
tri 4495 2854 4517 2876 se
rect 4517 2869 4532 2877
tri 4517 2854 4532 2869 nw
tri 4489 2848 4495 2854 se
rect 4495 2848 4504 2854
rect 4208 2763 4236 2773
tri 4236 2763 4260 2787 sw
rect 4154 2693 4170 2741
rect 4208 2731 4250 2763
tri 4267 2755 4268 2756 sw
rect 4267 2731 4268 2755
tri 4270 2754 4307 2791 ne
rect 4307 2763 4312 2791
tri 4312 2763 4338 2789 sw
rect 4422 2773 4431 2807
rect 4422 2763 4450 2773
rect 4307 2754 4391 2763
tri 4307 2735 4326 2754 ne
rect 4326 2735 4391 2754
rect 4208 2709 4268 2731
rect 4390 2731 4391 2735
rect 4408 2731 4450 2763
rect 4390 2709 4450 2731
rect 4296 2693 4313 2707
rect 4345 2693 4362 2707
tri 4133 2657 4155 2679 se
rect 4155 2672 4170 2693
tri 4155 2657 4170 2672 nw
rect 4489 2672 4504 2848
tri 4504 2841 4517 2854 nw
rect 4590 2773 4605 3001
tri 4127 2651 4133 2657 se
rect 4133 2651 4142 2657
rect 4127 2635 4142 2651
tri 4142 2644 4155 2657 nw
rect 4296 2649 4313 2663
rect 4345 2649 4362 2663
tri 4489 2657 4504 2672 ne
tri 4504 2657 4526 2679 sw
rect 4127 2599 4142 2607
rect 4208 2635 4268 2649
rect 4223 2625 4268 2635
rect 4223 2607 4251 2625
tri 4127 2584 4142 2599 ne
tri 4142 2584 4164 2606 sw
rect 4208 2597 4251 2607
rect 4266 2621 4268 2625
rect 4390 2635 4450 2649
tri 4504 2644 4517 2657 ne
rect 4517 2651 4526 2657
tri 4526 2651 4532 2657 sw
rect 4390 2625 4435 2635
rect 4266 2597 4340 2621
rect 4208 2593 4340 2597
tri 4340 2593 4368 2621 sw
rect 4390 2611 4392 2625
tri 4390 2609 4392 2611 ne
rect 4404 2607 4435 2625
rect 4404 2597 4450 2607
rect 4517 2636 4532 2651
tri 4142 2572 4154 2584 ne
rect 4154 2579 4164 2584
tri 4164 2579 4169 2584 sw
rect 4053 2233 4068 2461
rect 4154 2423 4169 2579
rect 4208 2537 4236 2593
tri 4328 2575 4346 2593 ne
rect 4346 2573 4368 2593
tri 4368 2573 4388 2593 sw
tri 4404 2579 4422 2597 ne
rect 4227 2503 4236 2537
rect 4270 2564 4312 2565
rect 4270 2530 4275 2564
rect 4305 2530 4312 2564
rect 4270 2521 4312 2530
rect 4346 2564 4388 2573
rect 4346 2530 4353 2564
rect 4383 2530 4388 2564
rect 4346 2525 4388 2530
rect 4422 2537 4450 2597
tri 4495 2584 4517 2606 se
rect 4517 2599 4532 2607
tri 4517 2584 4532 2599 nw
tri 4489 2578 4495 2584 se
rect 4495 2578 4504 2584
rect 4208 2493 4236 2503
tri 4236 2493 4260 2517 sw
rect 4208 2461 4250 2493
tri 4267 2485 4268 2486 sw
rect 4267 2461 4268 2485
tri 4270 2484 4307 2521 ne
rect 4307 2493 4312 2521
tri 4312 2493 4338 2519 sw
rect 4422 2503 4431 2537
rect 4422 2493 4450 2503
rect 4307 2484 4391 2493
tri 4307 2465 4326 2484 ne
rect 4326 2465 4391 2484
rect 4208 2439 4268 2461
rect 4390 2461 4391 2465
rect 4408 2461 4450 2493
rect 4390 2439 4450 2461
rect 4296 2423 4313 2437
rect 4345 2423 4362 2437
tri 4133 2387 4155 2409 se
rect 4155 2402 4170 2423
tri 4155 2387 4170 2402 nw
rect 4489 2402 4504 2578
tri 4504 2571 4517 2584 nw
rect 4590 2503 4605 2731
tri 4127 2381 4133 2387 se
rect 4133 2381 4142 2387
rect 4127 2365 4142 2381
tri 4142 2374 4155 2387 nw
rect 4296 2379 4313 2393
rect 4345 2379 4362 2393
tri 4489 2387 4504 2402 ne
tri 4504 2387 4526 2409 sw
rect 4127 2329 4142 2337
rect 4208 2365 4268 2379
rect 4223 2355 4268 2365
rect 4223 2337 4251 2355
tri 4127 2314 4142 2329 ne
tri 4142 2314 4164 2336 sw
rect 4208 2327 4251 2337
rect 4266 2351 4268 2355
rect 4390 2365 4450 2379
tri 4504 2374 4517 2387 ne
rect 4517 2381 4526 2387
tri 4526 2381 4532 2387 sw
rect 4390 2355 4435 2365
rect 4266 2327 4340 2351
rect 4208 2323 4340 2327
tri 4340 2323 4368 2351 sw
rect 4390 2341 4392 2355
tri 4390 2339 4392 2341 ne
rect 4404 2337 4435 2355
rect 4404 2327 4450 2337
rect 4517 2366 4532 2381
tri 4142 2302 4154 2314 ne
rect 4154 2309 4164 2314
tri 4164 2309 4169 2314 sw
rect 4053 1963 4068 2191
rect 4154 2201 4169 2309
rect 4208 2267 4236 2323
tri 4328 2305 4346 2323 ne
rect 4346 2303 4368 2323
tri 4368 2303 4388 2323 sw
tri 4404 2309 4422 2327 ne
rect 4227 2233 4236 2267
rect 4270 2294 4312 2295
rect 4270 2260 4275 2294
rect 4305 2260 4312 2294
rect 4270 2251 4312 2260
rect 4346 2294 4388 2303
rect 4346 2260 4353 2294
rect 4383 2260 4388 2294
rect 4346 2255 4388 2260
rect 4422 2267 4450 2327
tri 4495 2314 4517 2336 se
rect 4517 2329 4532 2337
tri 4517 2314 4532 2329 nw
tri 4489 2308 4495 2314 se
rect 4495 2308 4504 2314
rect 4208 2223 4236 2233
tri 4236 2223 4260 2247 sw
rect 4154 2153 4170 2201
rect 4208 2191 4250 2223
tri 4267 2215 4268 2216 sw
rect 4267 2191 4268 2215
tri 4270 2214 4307 2251 ne
rect 4307 2223 4312 2251
tri 4312 2223 4338 2249 sw
rect 4422 2233 4431 2267
rect 4422 2223 4450 2233
rect 4307 2214 4391 2223
tri 4307 2195 4326 2214 ne
rect 4326 2195 4391 2214
rect 4208 2169 4268 2191
rect 4390 2191 4391 2195
rect 4408 2191 4450 2223
rect 4390 2169 4450 2191
rect 4296 2153 4313 2167
rect 4345 2153 4362 2167
tri 4133 2117 4155 2139 se
rect 4155 2132 4170 2153
tri 4155 2117 4170 2132 nw
rect 4489 2132 4504 2308
tri 4504 2301 4517 2314 nw
rect 4590 2233 4605 2461
tri 4127 2111 4133 2117 se
rect 4133 2111 4142 2117
rect 4127 2095 4142 2111
tri 4142 2104 4155 2117 nw
rect 4296 2109 4313 2123
rect 4345 2109 4362 2123
tri 4489 2117 4504 2132 ne
tri 4504 2117 4526 2139 sw
rect 4127 2059 4142 2067
rect 4208 2095 4268 2109
rect 4223 2085 4268 2095
rect 4223 2067 4251 2085
tri 4127 2044 4142 2059 ne
tri 4142 2044 4164 2066 sw
rect 4208 2057 4251 2067
rect 4266 2081 4268 2085
rect 4390 2095 4450 2109
tri 4504 2104 4517 2117 ne
rect 4517 2111 4526 2117
tri 4526 2111 4532 2117 sw
rect 4390 2085 4435 2095
rect 4266 2057 4340 2081
rect 4208 2053 4340 2057
tri 4340 2053 4368 2081 sw
rect 4390 2071 4392 2085
tri 4390 2069 4392 2071 ne
rect 4404 2067 4435 2085
rect 4404 2057 4450 2067
rect 4517 2096 4532 2111
tri 4142 2032 4154 2044 ne
rect 4154 2039 4164 2044
tri 4164 2039 4169 2044 sw
rect 4053 1693 4068 1921
rect 4154 1883 4169 2039
rect 4208 1997 4236 2053
tri 4328 2035 4346 2053 ne
rect 4346 2033 4368 2053
tri 4368 2033 4388 2053 sw
tri 4404 2039 4422 2057 ne
rect 4227 1963 4236 1997
rect 4270 2024 4312 2025
rect 4270 1990 4275 2024
rect 4305 1990 4312 2024
rect 4270 1981 4312 1990
rect 4346 2024 4388 2033
rect 4346 1990 4353 2024
rect 4383 1990 4388 2024
rect 4346 1985 4388 1990
rect 4422 1997 4450 2057
tri 4495 2044 4517 2066 se
rect 4517 2059 4532 2067
tri 4517 2044 4532 2059 nw
tri 4489 2038 4495 2044 se
rect 4495 2038 4504 2044
rect 4208 1953 4236 1963
tri 4236 1953 4260 1977 sw
rect 4208 1921 4250 1953
tri 4267 1945 4268 1946 sw
rect 4267 1921 4268 1945
tri 4270 1944 4307 1981 ne
rect 4307 1953 4312 1981
tri 4312 1953 4338 1979 sw
rect 4422 1963 4431 1997
rect 4422 1953 4450 1963
rect 4307 1944 4391 1953
tri 4307 1925 4326 1944 ne
rect 4326 1925 4391 1944
rect 4208 1899 4268 1921
rect 4390 1921 4391 1925
rect 4408 1921 4450 1953
rect 4390 1899 4450 1921
rect 4296 1883 4313 1897
rect 4345 1883 4362 1897
tri 4133 1847 4155 1869 se
rect 4155 1862 4170 1883
tri 4155 1847 4170 1862 nw
rect 4489 1862 4504 2038
tri 4504 2031 4517 2044 nw
rect 4590 1963 4605 2191
tri 4127 1841 4133 1847 se
rect 4133 1841 4142 1847
rect 4127 1825 4142 1841
tri 4142 1834 4155 1847 nw
rect 4296 1839 4313 1853
rect 4345 1839 4362 1853
tri 4489 1847 4504 1862 ne
tri 4504 1847 4526 1869 sw
rect 4127 1789 4142 1797
rect 4208 1825 4268 1839
rect 4223 1815 4268 1825
rect 4223 1797 4251 1815
tri 4127 1774 4142 1789 ne
tri 4142 1774 4164 1796 sw
rect 4208 1787 4251 1797
rect 4266 1811 4268 1815
rect 4390 1825 4450 1839
tri 4504 1834 4517 1847 ne
rect 4517 1841 4526 1847
tri 4526 1841 4532 1847 sw
rect 4390 1815 4435 1825
rect 4266 1787 4340 1811
rect 4208 1783 4340 1787
tri 4340 1783 4368 1811 sw
rect 4390 1801 4392 1815
tri 4390 1799 4392 1801 ne
rect 4404 1797 4435 1815
rect 4404 1787 4450 1797
rect 4517 1826 4532 1841
tri 4142 1762 4154 1774 ne
rect 4154 1769 4164 1774
tri 4164 1769 4169 1774 sw
rect 4053 1423 4068 1651
rect 4154 1661 4169 1769
rect 4208 1727 4236 1783
tri 4328 1765 4346 1783 ne
rect 4346 1763 4368 1783
tri 4368 1763 4388 1783 sw
tri 4404 1769 4422 1787 ne
rect 4227 1693 4236 1727
rect 4270 1754 4312 1755
rect 4270 1720 4275 1754
rect 4305 1720 4312 1754
rect 4270 1711 4312 1720
rect 4346 1754 4388 1763
rect 4346 1720 4353 1754
rect 4383 1720 4388 1754
rect 4346 1715 4388 1720
rect 4422 1727 4450 1787
tri 4495 1774 4517 1796 se
rect 4517 1789 4532 1797
tri 4517 1774 4532 1789 nw
tri 4489 1768 4495 1774 se
rect 4495 1768 4504 1774
rect 4208 1683 4236 1693
tri 4236 1683 4260 1707 sw
rect 4154 1613 4170 1661
rect 4208 1651 4250 1683
tri 4267 1675 4268 1676 sw
rect 4267 1651 4268 1675
tri 4270 1674 4307 1711 ne
rect 4307 1683 4312 1711
tri 4312 1683 4338 1709 sw
rect 4422 1693 4431 1727
rect 4422 1683 4450 1693
rect 4307 1674 4391 1683
tri 4307 1655 4326 1674 ne
rect 4326 1655 4391 1674
rect 4208 1629 4268 1651
rect 4390 1651 4391 1655
rect 4408 1651 4450 1683
rect 4390 1629 4450 1651
rect 4296 1613 4313 1627
rect 4345 1613 4362 1627
tri 4133 1577 4155 1599 se
rect 4155 1592 4170 1613
tri 4155 1577 4170 1592 nw
rect 4489 1592 4504 1768
tri 4504 1761 4517 1774 nw
rect 4590 1693 4605 1921
tri 4127 1571 4133 1577 se
rect 4133 1571 4142 1577
rect 4127 1555 4142 1571
tri 4142 1564 4155 1577 nw
rect 4296 1569 4313 1583
rect 4345 1569 4362 1583
tri 4489 1577 4504 1592 ne
tri 4504 1577 4526 1599 sw
rect 4127 1519 4142 1527
rect 4208 1555 4268 1569
rect 4223 1545 4268 1555
rect 4223 1527 4251 1545
tri 4127 1504 4142 1519 ne
tri 4142 1504 4164 1526 sw
rect 4208 1517 4251 1527
rect 4266 1541 4268 1545
rect 4390 1555 4450 1569
tri 4504 1564 4517 1577 ne
rect 4517 1571 4526 1577
tri 4526 1571 4532 1577 sw
rect 4390 1545 4435 1555
rect 4266 1517 4340 1541
rect 4208 1513 4340 1517
tri 4340 1513 4368 1541 sw
rect 4390 1531 4392 1545
tri 4390 1529 4392 1531 ne
rect 4404 1527 4435 1545
rect 4404 1517 4450 1527
rect 4517 1556 4532 1571
tri 4142 1492 4154 1504 ne
rect 4154 1499 4164 1504
tri 4164 1499 4169 1504 sw
rect 4053 1153 4068 1381
rect 4154 1343 4169 1499
rect 4208 1457 4236 1513
tri 4328 1495 4346 1513 ne
rect 4346 1493 4368 1513
tri 4368 1493 4388 1513 sw
tri 4404 1499 4422 1517 ne
rect 4227 1423 4236 1457
rect 4270 1484 4312 1485
rect 4270 1450 4275 1484
rect 4305 1450 4312 1484
rect 4270 1441 4312 1450
rect 4346 1484 4388 1493
rect 4346 1450 4353 1484
rect 4383 1450 4388 1484
rect 4346 1445 4388 1450
rect 4422 1457 4450 1517
tri 4495 1504 4517 1526 se
rect 4517 1519 4532 1527
tri 4517 1504 4532 1519 nw
tri 4489 1498 4495 1504 se
rect 4495 1498 4504 1504
rect 4208 1413 4236 1423
tri 4236 1413 4260 1437 sw
rect 4208 1381 4250 1413
tri 4267 1405 4268 1406 sw
rect 4267 1381 4268 1405
tri 4270 1404 4307 1441 ne
rect 4307 1413 4312 1441
tri 4312 1413 4338 1439 sw
rect 4422 1423 4431 1457
rect 4422 1413 4450 1423
rect 4307 1404 4391 1413
tri 4307 1385 4326 1404 ne
rect 4326 1385 4391 1404
rect 4208 1359 4268 1381
rect 4390 1381 4391 1385
rect 4408 1381 4450 1413
rect 4390 1359 4450 1381
rect 4296 1343 4313 1357
rect 4345 1343 4362 1357
tri 4133 1307 4155 1329 se
rect 4155 1322 4170 1343
tri 4155 1307 4170 1322 nw
rect 4489 1322 4504 1498
tri 4504 1491 4517 1504 nw
rect 4590 1423 4605 1651
tri 4127 1301 4133 1307 se
rect 4133 1301 4142 1307
rect 4127 1285 4142 1301
tri 4142 1294 4155 1307 nw
rect 4296 1299 4313 1313
rect 4345 1299 4362 1313
tri 4489 1307 4504 1322 ne
tri 4504 1307 4526 1329 sw
rect 4127 1249 4142 1257
rect 4208 1285 4268 1299
rect 4223 1275 4268 1285
rect 4223 1257 4251 1275
tri 4127 1234 4142 1249 ne
tri 4142 1234 4164 1256 sw
rect 4208 1247 4251 1257
rect 4266 1271 4268 1275
rect 4390 1285 4450 1299
tri 4504 1294 4517 1307 ne
rect 4517 1301 4526 1307
tri 4526 1301 4532 1307 sw
rect 4390 1275 4435 1285
rect 4266 1247 4340 1271
rect 4208 1243 4340 1247
tri 4340 1243 4368 1271 sw
rect 4390 1261 4392 1275
tri 4390 1259 4392 1261 ne
rect 4404 1257 4435 1275
rect 4404 1247 4450 1257
rect 4517 1286 4532 1301
tri 4142 1222 4154 1234 ne
rect 4154 1229 4164 1234
tri 4164 1229 4169 1234 sw
rect 4053 883 4068 1111
rect 4154 1121 4169 1229
rect 4208 1187 4236 1243
tri 4328 1225 4346 1243 ne
rect 4346 1223 4368 1243
tri 4368 1223 4388 1243 sw
tri 4404 1229 4422 1247 ne
rect 4227 1153 4236 1187
rect 4270 1214 4312 1215
rect 4270 1180 4275 1214
rect 4305 1180 4312 1214
rect 4270 1171 4312 1180
rect 4346 1214 4388 1223
rect 4346 1180 4353 1214
rect 4383 1180 4388 1214
rect 4346 1175 4388 1180
rect 4422 1187 4450 1247
tri 4495 1234 4517 1256 se
rect 4517 1249 4532 1257
tri 4517 1234 4532 1249 nw
tri 4489 1228 4495 1234 se
rect 4495 1228 4504 1234
rect 4208 1143 4236 1153
tri 4236 1143 4260 1167 sw
rect 4154 1073 4170 1121
rect 4208 1111 4250 1143
tri 4267 1135 4268 1136 sw
rect 4267 1111 4268 1135
tri 4270 1134 4307 1171 ne
rect 4307 1143 4312 1171
tri 4312 1143 4338 1169 sw
rect 4422 1153 4431 1187
rect 4422 1143 4450 1153
rect 4307 1134 4391 1143
tri 4307 1115 4326 1134 ne
rect 4326 1115 4391 1134
rect 4208 1089 4268 1111
rect 4390 1111 4391 1115
rect 4408 1111 4450 1143
rect 4390 1089 4450 1111
rect 4296 1073 4313 1087
rect 4345 1073 4362 1087
tri 4133 1037 4155 1059 se
rect 4155 1052 4170 1073
tri 4155 1037 4170 1052 nw
rect 4489 1052 4504 1228
tri 4504 1221 4517 1234 nw
rect 4590 1153 4605 1381
tri 4127 1031 4133 1037 se
rect 4133 1031 4142 1037
rect 4127 1015 4142 1031
tri 4142 1024 4155 1037 nw
rect 4296 1029 4313 1043
rect 4345 1029 4362 1043
tri 4489 1037 4504 1052 ne
tri 4504 1037 4526 1059 sw
rect 4127 979 4142 987
rect 4208 1015 4268 1029
rect 4223 1005 4268 1015
rect 4223 987 4251 1005
tri 4127 964 4142 979 ne
tri 4142 964 4164 986 sw
rect 4208 977 4251 987
rect 4266 1001 4268 1005
rect 4390 1015 4450 1029
tri 4504 1024 4517 1037 ne
rect 4517 1031 4526 1037
tri 4526 1031 4532 1037 sw
rect 4390 1005 4435 1015
rect 4266 977 4340 1001
rect 4208 973 4340 977
tri 4340 973 4368 1001 sw
rect 4390 991 4392 1005
tri 4390 989 4392 991 ne
rect 4404 987 4435 1005
rect 4404 977 4450 987
rect 4517 1016 4532 1031
tri 4142 952 4154 964 ne
rect 4154 959 4164 964
tri 4164 959 4169 964 sw
rect 4053 613 4068 841
rect 4154 803 4169 959
rect 4208 917 4236 973
tri 4328 955 4346 973 ne
rect 4346 953 4368 973
tri 4368 953 4388 973 sw
tri 4404 959 4422 977 ne
rect 4227 883 4236 917
rect 4270 944 4312 945
rect 4270 910 4275 944
rect 4305 910 4312 944
rect 4270 901 4312 910
rect 4346 944 4388 953
rect 4346 910 4353 944
rect 4383 910 4388 944
rect 4346 905 4388 910
rect 4422 917 4450 977
tri 4495 964 4517 986 se
rect 4517 979 4532 987
tri 4517 964 4532 979 nw
tri 4489 958 4495 964 se
rect 4495 958 4504 964
rect 4208 873 4236 883
tri 4236 873 4260 897 sw
rect 4208 841 4250 873
tri 4267 865 4268 866 sw
rect 4267 841 4268 865
tri 4270 864 4307 901 ne
rect 4307 873 4312 901
tri 4312 873 4338 899 sw
rect 4422 883 4431 917
rect 4422 873 4450 883
rect 4307 864 4391 873
tri 4307 845 4326 864 ne
rect 4326 845 4391 864
rect 4208 819 4268 841
rect 4390 841 4391 845
rect 4408 841 4450 873
rect 4390 819 4450 841
rect 4296 803 4313 817
rect 4345 803 4362 817
tri 4133 767 4155 789 se
rect 4155 782 4170 803
tri 4155 767 4170 782 nw
rect 4489 782 4504 958
tri 4504 951 4517 964 nw
rect 4590 883 4605 1111
tri 4127 761 4133 767 se
rect 4133 761 4142 767
rect 4127 745 4142 761
tri 4142 754 4155 767 nw
rect 4296 759 4313 773
rect 4345 759 4362 773
tri 4489 767 4504 782 ne
tri 4504 767 4526 789 sw
rect 4127 709 4142 717
rect 4208 745 4268 759
rect 4223 735 4268 745
rect 4223 717 4251 735
tri 4127 694 4142 709 ne
tri 4142 694 4164 716 sw
rect 4208 707 4251 717
rect 4266 731 4268 735
rect 4390 745 4450 759
tri 4504 754 4517 767 ne
rect 4517 761 4526 767
tri 4526 761 4532 767 sw
rect 4390 735 4435 745
rect 4266 707 4340 731
rect 4208 703 4340 707
tri 4340 703 4368 731 sw
rect 4390 721 4392 735
tri 4390 719 4392 721 ne
rect 4404 717 4435 735
rect 4404 707 4450 717
rect 4517 746 4532 761
tri 4142 682 4154 694 ne
rect 4154 689 4164 694
tri 4164 689 4169 694 sw
rect 4053 343 4068 571
rect 4154 581 4169 689
rect 4208 647 4236 703
tri 4328 685 4346 703 ne
rect 4346 683 4368 703
tri 4368 683 4388 703 sw
tri 4404 689 4422 707 ne
rect 4227 613 4236 647
rect 4270 674 4312 675
rect 4270 640 4275 674
rect 4305 640 4312 674
rect 4270 631 4312 640
rect 4346 674 4388 683
rect 4346 640 4353 674
rect 4383 640 4388 674
rect 4346 635 4388 640
rect 4422 647 4450 707
tri 4495 694 4517 716 se
rect 4517 709 4532 717
tri 4517 694 4532 709 nw
tri 4489 688 4495 694 se
rect 4495 688 4504 694
rect 4208 603 4236 613
tri 4236 603 4260 627 sw
rect 4154 533 4170 581
rect 4208 571 4250 603
tri 4267 595 4268 596 sw
rect 4267 571 4268 595
tri 4270 594 4307 631 ne
rect 4307 603 4312 631
tri 4312 603 4338 629 sw
rect 4422 613 4431 647
rect 4422 603 4450 613
rect 4307 594 4391 603
tri 4307 575 4326 594 ne
rect 4326 575 4391 594
rect 4208 549 4268 571
rect 4390 571 4391 575
rect 4408 571 4450 603
rect 4390 549 4450 571
rect 4296 533 4313 547
rect 4345 533 4362 547
tri 4133 497 4155 519 se
rect 4155 512 4170 533
tri 4155 497 4170 512 nw
rect 4489 512 4504 688
tri 4504 681 4517 694 nw
rect 4590 613 4605 841
tri 4127 491 4133 497 se
rect 4133 491 4142 497
rect 4127 475 4142 491
tri 4142 484 4155 497 nw
rect 4296 489 4313 503
rect 4345 489 4362 503
tri 4489 497 4504 512 ne
tri 4504 497 4526 519 sw
rect 4127 439 4142 447
rect 4208 475 4268 489
rect 4223 465 4268 475
rect 4223 447 4251 465
tri 4127 424 4142 439 ne
tri 4142 424 4164 446 sw
rect 4208 437 4251 447
rect 4266 461 4268 465
rect 4390 475 4450 489
tri 4504 484 4517 497 ne
rect 4517 491 4526 497
tri 4526 491 4532 497 sw
rect 4390 465 4435 475
rect 4266 437 4340 461
rect 4208 433 4340 437
tri 4340 433 4368 461 sw
rect 4390 451 4392 465
tri 4390 449 4392 451 ne
rect 4404 447 4435 465
rect 4404 437 4450 447
rect 4517 476 4532 491
tri 4142 412 4154 424 ne
rect 4154 419 4164 424
tri 4164 419 4169 424 sw
rect 4053 73 4068 301
rect 4154 263 4169 419
rect 4208 377 4236 433
tri 4328 415 4346 433 ne
rect 4346 413 4368 433
tri 4368 413 4388 433 sw
tri 4404 419 4422 437 ne
rect 4227 343 4236 377
rect 4270 404 4312 405
rect 4270 370 4275 404
rect 4305 370 4312 404
rect 4270 361 4312 370
rect 4346 404 4388 413
rect 4346 370 4353 404
rect 4383 370 4388 404
rect 4346 365 4388 370
rect 4422 377 4450 437
tri 4495 424 4517 446 se
rect 4517 439 4532 447
tri 4517 424 4532 439 nw
tri 4489 418 4495 424 se
rect 4495 418 4504 424
rect 4208 333 4236 343
tri 4236 333 4260 357 sw
rect 4208 301 4250 333
tri 4267 325 4268 326 sw
rect 4267 301 4268 325
tri 4270 324 4307 361 ne
rect 4307 333 4312 361
tri 4312 333 4338 359 sw
rect 4422 343 4431 377
rect 4422 333 4450 343
rect 4307 324 4391 333
tri 4307 305 4326 324 ne
rect 4326 305 4391 324
rect 4208 279 4268 301
rect 4390 301 4391 305
rect 4408 301 4450 333
rect 4390 279 4450 301
rect 4296 263 4313 277
rect 4345 263 4362 277
tri 4133 227 4155 249 se
rect 4155 242 4170 263
tri 4155 227 4170 242 nw
rect 4489 242 4504 418
tri 4504 411 4517 424 nw
rect 4590 343 4605 571
tri 4127 221 4133 227 se
rect 4133 221 4142 227
rect 4127 205 4142 221
tri 4142 214 4155 227 nw
rect 4296 219 4313 233
rect 4345 219 4362 233
tri 4489 227 4504 242 ne
tri 4504 227 4526 249 sw
rect 4127 169 4142 177
rect 4208 205 4268 219
rect 4223 195 4268 205
rect 4223 177 4251 195
tri 4127 154 4142 169 ne
tri 4142 154 4164 176 sw
rect 4208 167 4251 177
rect 4266 191 4268 195
rect 4390 205 4450 219
tri 4504 214 4517 227 ne
rect 4517 221 4526 227
tri 4526 221 4532 227 sw
rect 4390 195 4435 205
rect 4266 167 4340 191
rect 4208 163 4340 167
tri 4340 163 4368 191 sw
rect 4390 181 4392 195
tri 4390 179 4392 181 ne
rect 4404 177 4435 195
rect 4404 167 4450 177
rect 4517 206 4532 221
tri 4142 142 4154 154 ne
rect 4154 149 4164 154
tri 4164 149 4169 154 sw
rect 4053 -55 4068 31
rect 4154 -55 4169 149
rect 4208 107 4236 163
tri 4328 145 4346 163 ne
rect 4346 143 4368 163
tri 4368 143 4388 163 sw
tri 4404 149 4422 167 ne
rect 4227 73 4236 107
rect 4270 134 4312 135
rect 4270 100 4275 134
rect 4305 100 4312 134
rect 4270 91 4312 100
rect 4346 134 4388 143
rect 4346 100 4353 134
rect 4383 100 4388 134
rect 4346 95 4388 100
rect 4422 107 4450 167
tri 4495 154 4517 176 se
rect 4517 169 4532 177
tri 4517 154 4532 169 nw
tri 4489 148 4495 154 se
rect 4495 148 4504 154
rect 4208 63 4236 73
tri 4236 63 4260 87 sw
rect 4208 31 4250 63
tri 4267 55 4268 56 sw
rect 4267 31 4268 55
tri 4270 54 4307 91 ne
rect 4307 63 4312 91
tri 4312 63 4338 89 sw
rect 4422 73 4431 107
rect 4422 63 4450 73
rect 4307 54 4391 63
tri 4307 35 4326 54 ne
rect 4326 35 4391 54
rect 4208 9 4268 31
rect 4390 31 4391 35
rect 4408 31 4450 63
rect 4390 9 4450 31
rect 4296 -7 4313 7
rect 4345 -7 4362 7
rect 4489 -55 4504 148
tri 4504 141 4517 154 nw
rect 4590 73 4605 301
rect 4590 -55 4605 31
rect 4633 4123 4648 4361
tri 4713 4277 4735 4299 se
rect 4735 4292 4750 4361
tri 4735 4277 4750 4292 nw
rect 5069 4292 5084 4361
tri 4707 4271 4713 4277 se
rect 4713 4271 4722 4277
rect 4707 4255 4722 4271
tri 4722 4264 4735 4277 nw
rect 4876 4269 4893 4283
rect 4925 4269 4942 4283
tri 5069 4277 5084 4292 ne
tri 5084 4277 5106 4299 sw
rect 4707 4219 4722 4227
rect 4788 4255 4848 4269
rect 4803 4245 4848 4255
rect 4803 4227 4831 4245
tri 4707 4204 4722 4219 ne
tri 4722 4204 4744 4226 sw
rect 4788 4217 4831 4227
rect 4846 4241 4848 4245
rect 4970 4255 5030 4269
tri 5084 4264 5097 4277 ne
rect 5097 4271 5106 4277
tri 5106 4271 5112 4277 sw
rect 4970 4245 5015 4255
rect 4846 4217 4920 4241
rect 4788 4213 4920 4217
tri 4920 4213 4948 4241 sw
rect 4970 4231 4972 4245
tri 4970 4229 4972 4231 ne
rect 4984 4227 5015 4245
rect 4984 4217 5030 4227
rect 5097 4256 5112 4271
tri 4722 4192 4734 4204 ne
rect 4734 4199 4744 4204
tri 4744 4199 4749 4204 sw
rect 4633 3853 4648 4081
rect 4734 4043 4749 4199
rect 4788 4157 4816 4213
tri 4908 4195 4926 4213 ne
rect 4926 4193 4948 4213
tri 4948 4193 4968 4213 sw
tri 4984 4199 5002 4217 ne
rect 4807 4123 4816 4157
rect 4850 4184 4892 4185
rect 4850 4150 4855 4184
rect 4885 4150 4892 4184
rect 4850 4141 4892 4150
rect 4926 4184 4968 4193
rect 4926 4150 4933 4184
rect 4963 4150 4968 4184
rect 4926 4145 4968 4150
rect 5002 4157 5030 4217
tri 5075 4204 5097 4226 se
rect 5097 4219 5112 4227
tri 5097 4204 5112 4219 nw
tri 5069 4198 5075 4204 se
rect 5075 4198 5084 4204
rect 4788 4113 4816 4123
tri 4816 4113 4840 4137 sw
rect 4788 4081 4830 4113
tri 4847 4105 4848 4106 sw
rect 4847 4081 4848 4105
tri 4850 4104 4887 4141 ne
rect 4887 4113 4892 4141
tri 4892 4113 4918 4139 sw
rect 5002 4123 5011 4157
rect 5002 4113 5030 4123
rect 4887 4104 4971 4113
tri 4887 4085 4906 4104 ne
rect 4906 4085 4971 4104
rect 4788 4059 4848 4081
rect 4970 4081 4971 4085
rect 4988 4081 5030 4113
rect 4970 4059 5030 4081
rect 4876 4043 4893 4057
rect 4925 4043 4942 4057
tri 4713 4007 4735 4029 se
rect 4735 4022 4750 4043
tri 4735 4007 4750 4022 nw
rect 5069 4022 5084 4198
tri 5084 4191 5097 4204 nw
rect 5170 4123 5185 4361
tri 4707 4001 4713 4007 se
rect 4713 4001 4722 4007
rect 4707 3985 4722 4001
tri 4722 3994 4735 4007 nw
rect 4876 3999 4893 4013
rect 4925 3999 4942 4013
tri 5069 4007 5084 4022 ne
tri 5084 4007 5106 4029 sw
rect 4707 3949 4722 3957
rect 4788 3985 4848 3999
rect 4803 3975 4848 3985
rect 4803 3957 4831 3975
tri 4707 3934 4722 3949 ne
tri 4722 3934 4744 3956 sw
rect 4788 3947 4831 3957
rect 4846 3971 4848 3975
rect 4970 3985 5030 3999
tri 5084 3994 5097 4007 ne
rect 5097 4001 5106 4007
tri 5106 4001 5112 4007 sw
rect 4970 3975 5015 3985
rect 4846 3947 4920 3971
rect 4788 3943 4920 3947
tri 4920 3943 4948 3971 sw
rect 4970 3961 4972 3975
tri 4970 3959 4972 3961 ne
rect 4984 3957 5015 3975
rect 4984 3947 5030 3957
rect 5097 3986 5112 4001
tri 4722 3922 4734 3934 ne
rect 4734 3929 4744 3934
tri 4744 3929 4749 3934 sw
rect 4633 3583 4648 3811
rect 4734 3821 4749 3929
rect 4788 3887 4816 3943
tri 4908 3925 4926 3943 ne
rect 4926 3923 4948 3943
tri 4948 3923 4968 3943 sw
tri 4984 3929 5002 3947 ne
rect 4807 3853 4816 3887
rect 4850 3914 4892 3915
rect 4850 3880 4855 3914
rect 4885 3880 4892 3914
rect 4850 3871 4892 3880
rect 4926 3914 4968 3923
rect 4926 3880 4933 3914
rect 4963 3880 4968 3914
rect 4926 3875 4968 3880
rect 5002 3887 5030 3947
tri 5075 3934 5097 3956 se
rect 5097 3949 5112 3957
tri 5097 3934 5112 3949 nw
tri 5069 3928 5075 3934 se
rect 5075 3928 5084 3934
rect 4788 3843 4816 3853
tri 4816 3843 4840 3867 sw
rect 4734 3773 4750 3821
rect 4788 3811 4830 3843
tri 4847 3835 4848 3836 sw
rect 4847 3811 4848 3835
tri 4850 3834 4887 3871 ne
rect 4887 3843 4892 3871
tri 4892 3843 4918 3869 sw
rect 5002 3853 5011 3887
rect 5002 3843 5030 3853
rect 4887 3834 4971 3843
tri 4887 3815 4906 3834 ne
rect 4906 3815 4971 3834
rect 4788 3789 4848 3811
rect 4970 3811 4971 3815
rect 4988 3811 5030 3843
rect 4970 3789 5030 3811
rect 4876 3773 4893 3787
rect 4925 3773 4942 3787
tri 4713 3737 4735 3759 se
rect 4735 3752 4750 3773
tri 4735 3737 4750 3752 nw
rect 5069 3752 5084 3928
tri 5084 3921 5097 3934 nw
rect 5170 3853 5185 4081
tri 4707 3731 4713 3737 se
rect 4713 3731 4722 3737
rect 4707 3715 4722 3731
tri 4722 3724 4735 3737 nw
rect 4876 3729 4893 3743
rect 4925 3729 4942 3743
tri 5069 3737 5084 3752 ne
tri 5084 3737 5106 3759 sw
rect 4707 3679 4722 3687
rect 4788 3715 4848 3729
rect 4803 3705 4848 3715
rect 4803 3687 4831 3705
tri 4707 3664 4722 3679 ne
tri 4722 3664 4744 3686 sw
rect 4788 3677 4831 3687
rect 4846 3701 4848 3705
rect 4970 3715 5030 3729
tri 5084 3724 5097 3737 ne
rect 5097 3731 5106 3737
tri 5106 3731 5112 3737 sw
rect 4970 3705 5015 3715
rect 4846 3677 4920 3701
rect 4788 3673 4920 3677
tri 4920 3673 4948 3701 sw
rect 4970 3691 4972 3705
tri 4970 3689 4972 3691 ne
rect 4984 3687 5015 3705
rect 4984 3677 5030 3687
rect 5097 3716 5112 3731
tri 4722 3652 4734 3664 ne
rect 4734 3659 4744 3664
tri 4744 3659 4749 3664 sw
rect 4633 3313 4648 3541
rect 4734 3503 4749 3659
rect 4788 3617 4816 3673
tri 4908 3655 4926 3673 ne
rect 4926 3653 4948 3673
tri 4948 3653 4968 3673 sw
tri 4984 3659 5002 3677 ne
rect 4807 3583 4816 3617
rect 4850 3644 4892 3645
rect 4850 3610 4855 3644
rect 4885 3610 4892 3644
rect 4850 3601 4892 3610
rect 4926 3644 4968 3653
rect 4926 3610 4933 3644
rect 4963 3610 4968 3644
rect 4926 3605 4968 3610
rect 5002 3617 5030 3677
tri 5075 3664 5097 3686 se
rect 5097 3679 5112 3687
tri 5097 3664 5112 3679 nw
tri 5069 3658 5075 3664 se
rect 5075 3658 5084 3664
rect 4788 3573 4816 3583
tri 4816 3573 4840 3597 sw
rect 4788 3541 4830 3573
tri 4847 3565 4848 3566 sw
rect 4847 3541 4848 3565
tri 4850 3564 4887 3601 ne
rect 4887 3573 4892 3601
tri 4892 3573 4918 3599 sw
rect 5002 3583 5011 3617
rect 5002 3573 5030 3583
rect 4887 3564 4971 3573
tri 4887 3545 4906 3564 ne
rect 4906 3545 4971 3564
rect 4788 3519 4848 3541
rect 4970 3541 4971 3545
rect 4988 3541 5030 3573
rect 4970 3519 5030 3541
rect 4876 3503 4893 3517
rect 4925 3503 4942 3517
tri 4713 3467 4735 3489 se
rect 4735 3482 4750 3503
tri 4735 3467 4750 3482 nw
rect 5069 3482 5084 3658
tri 5084 3651 5097 3664 nw
rect 5170 3583 5185 3811
tri 4707 3461 4713 3467 se
rect 4713 3461 4722 3467
rect 4707 3445 4722 3461
tri 4722 3454 4735 3467 nw
rect 4876 3459 4893 3473
rect 4925 3459 4942 3473
tri 5069 3467 5084 3482 ne
tri 5084 3467 5106 3489 sw
rect 4707 3409 4722 3417
rect 4788 3445 4848 3459
rect 4803 3435 4848 3445
rect 4803 3417 4831 3435
tri 4707 3394 4722 3409 ne
tri 4722 3394 4744 3416 sw
rect 4788 3407 4831 3417
rect 4846 3431 4848 3435
rect 4970 3445 5030 3459
tri 5084 3454 5097 3467 ne
rect 5097 3461 5106 3467
tri 5106 3461 5112 3467 sw
rect 4970 3435 5015 3445
rect 4846 3407 4920 3431
rect 4788 3403 4920 3407
tri 4920 3403 4948 3431 sw
rect 4970 3421 4972 3435
tri 4970 3419 4972 3421 ne
rect 4984 3417 5015 3435
rect 4984 3407 5030 3417
rect 5097 3446 5112 3461
tri 4722 3382 4734 3394 ne
rect 4734 3389 4744 3394
tri 4744 3389 4749 3394 sw
rect 4633 3043 4648 3271
rect 4734 3281 4749 3389
rect 4788 3347 4816 3403
tri 4908 3385 4926 3403 ne
rect 4926 3383 4948 3403
tri 4948 3383 4968 3403 sw
tri 4984 3389 5002 3407 ne
rect 4807 3313 4816 3347
rect 4850 3374 4892 3375
rect 4850 3340 4855 3374
rect 4885 3340 4892 3374
rect 4850 3331 4892 3340
rect 4926 3374 4968 3383
rect 4926 3340 4933 3374
rect 4963 3340 4968 3374
rect 4926 3335 4968 3340
rect 5002 3347 5030 3407
tri 5075 3394 5097 3416 se
rect 5097 3409 5112 3417
tri 5097 3394 5112 3409 nw
tri 5069 3388 5075 3394 se
rect 5075 3388 5084 3394
rect 4788 3303 4816 3313
tri 4816 3303 4840 3327 sw
rect 4734 3233 4750 3281
rect 4788 3271 4830 3303
tri 4847 3295 4848 3296 sw
rect 4847 3271 4848 3295
tri 4850 3294 4887 3331 ne
rect 4887 3303 4892 3331
tri 4892 3303 4918 3329 sw
rect 5002 3313 5011 3347
rect 5002 3303 5030 3313
rect 4887 3294 4971 3303
tri 4887 3275 4906 3294 ne
rect 4906 3275 4971 3294
rect 4788 3249 4848 3271
rect 4970 3271 4971 3275
rect 4988 3271 5030 3303
rect 4970 3249 5030 3271
rect 4876 3233 4893 3247
rect 4925 3233 4942 3247
tri 4713 3197 4735 3219 se
rect 4735 3212 4750 3233
tri 4735 3197 4750 3212 nw
rect 5069 3212 5084 3388
tri 5084 3381 5097 3394 nw
rect 5170 3313 5185 3541
tri 4707 3191 4713 3197 se
rect 4713 3191 4722 3197
rect 4707 3175 4722 3191
tri 4722 3184 4735 3197 nw
rect 4876 3189 4893 3203
rect 4925 3189 4942 3203
tri 5069 3197 5084 3212 ne
tri 5084 3197 5106 3219 sw
rect 4707 3139 4722 3147
rect 4788 3175 4848 3189
rect 4803 3165 4848 3175
rect 4803 3147 4831 3165
tri 4707 3124 4722 3139 ne
tri 4722 3124 4744 3146 sw
rect 4788 3137 4831 3147
rect 4846 3161 4848 3165
rect 4970 3175 5030 3189
tri 5084 3184 5097 3197 ne
rect 5097 3191 5106 3197
tri 5106 3191 5112 3197 sw
rect 4970 3165 5015 3175
rect 4846 3137 4920 3161
rect 4788 3133 4920 3137
tri 4920 3133 4948 3161 sw
rect 4970 3151 4972 3165
tri 4970 3149 4972 3151 ne
rect 4984 3147 5015 3165
rect 4984 3137 5030 3147
rect 5097 3176 5112 3191
tri 4722 3112 4734 3124 ne
rect 4734 3119 4744 3124
tri 4744 3119 4749 3124 sw
rect 4633 2773 4648 3001
rect 4734 2963 4749 3119
rect 4788 3077 4816 3133
tri 4908 3115 4926 3133 ne
rect 4926 3113 4948 3133
tri 4948 3113 4968 3133 sw
tri 4984 3119 5002 3137 ne
rect 4807 3043 4816 3077
rect 4850 3104 4892 3105
rect 4850 3070 4855 3104
rect 4885 3070 4892 3104
rect 4850 3061 4892 3070
rect 4926 3104 4968 3113
rect 4926 3070 4933 3104
rect 4963 3070 4968 3104
rect 4926 3065 4968 3070
rect 5002 3077 5030 3137
tri 5075 3124 5097 3146 se
rect 5097 3139 5112 3147
tri 5097 3124 5112 3139 nw
tri 5069 3118 5075 3124 se
rect 5075 3118 5084 3124
rect 4788 3033 4816 3043
tri 4816 3033 4840 3057 sw
rect 4788 3001 4830 3033
tri 4847 3025 4848 3026 sw
rect 4847 3001 4848 3025
tri 4850 3024 4887 3061 ne
rect 4887 3033 4892 3061
tri 4892 3033 4918 3059 sw
rect 5002 3043 5011 3077
rect 5002 3033 5030 3043
rect 4887 3024 4971 3033
tri 4887 3005 4906 3024 ne
rect 4906 3005 4971 3024
rect 4788 2979 4848 3001
rect 4970 3001 4971 3005
rect 4988 3001 5030 3033
rect 4970 2979 5030 3001
rect 4876 2963 4893 2977
rect 4925 2963 4942 2977
tri 4713 2927 4735 2949 se
rect 4735 2942 4750 2963
tri 4735 2927 4750 2942 nw
rect 5069 2942 5084 3118
tri 5084 3111 5097 3124 nw
rect 5170 3043 5185 3271
tri 4707 2921 4713 2927 se
rect 4713 2921 4722 2927
rect 4707 2905 4722 2921
tri 4722 2914 4735 2927 nw
rect 4876 2919 4893 2933
rect 4925 2919 4942 2933
tri 5069 2927 5084 2942 ne
tri 5084 2927 5106 2949 sw
rect 4707 2869 4722 2877
rect 4788 2905 4848 2919
rect 4803 2895 4848 2905
rect 4803 2877 4831 2895
tri 4707 2854 4722 2869 ne
tri 4722 2854 4744 2876 sw
rect 4788 2867 4831 2877
rect 4846 2891 4848 2895
rect 4970 2905 5030 2919
tri 5084 2914 5097 2927 ne
rect 5097 2921 5106 2927
tri 5106 2921 5112 2927 sw
rect 4970 2895 5015 2905
rect 4846 2867 4920 2891
rect 4788 2863 4920 2867
tri 4920 2863 4948 2891 sw
rect 4970 2881 4972 2895
tri 4970 2879 4972 2881 ne
rect 4984 2877 5015 2895
rect 4984 2867 5030 2877
rect 5097 2906 5112 2921
tri 4722 2842 4734 2854 ne
rect 4734 2849 4744 2854
tri 4744 2849 4749 2854 sw
rect 4633 2503 4648 2731
rect 4734 2741 4749 2849
rect 4788 2807 4816 2863
tri 4908 2845 4926 2863 ne
rect 4926 2843 4948 2863
tri 4948 2843 4968 2863 sw
tri 4984 2849 5002 2867 ne
rect 4807 2773 4816 2807
rect 4850 2834 4892 2835
rect 4850 2800 4855 2834
rect 4885 2800 4892 2834
rect 4850 2791 4892 2800
rect 4926 2834 4968 2843
rect 4926 2800 4933 2834
rect 4963 2800 4968 2834
rect 4926 2795 4968 2800
rect 5002 2807 5030 2867
tri 5075 2854 5097 2876 se
rect 5097 2869 5112 2877
tri 5097 2854 5112 2869 nw
tri 5069 2848 5075 2854 se
rect 5075 2848 5084 2854
rect 4788 2763 4816 2773
tri 4816 2763 4840 2787 sw
rect 4734 2693 4750 2741
rect 4788 2731 4830 2763
tri 4847 2755 4848 2756 sw
rect 4847 2731 4848 2755
tri 4850 2754 4887 2791 ne
rect 4887 2763 4892 2791
tri 4892 2763 4918 2789 sw
rect 5002 2773 5011 2807
rect 5002 2763 5030 2773
rect 4887 2754 4971 2763
tri 4887 2735 4906 2754 ne
rect 4906 2735 4971 2754
rect 4788 2709 4848 2731
rect 4970 2731 4971 2735
rect 4988 2731 5030 2763
rect 4970 2709 5030 2731
rect 4876 2693 4893 2707
rect 4925 2693 4942 2707
tri 4713 2657 4735 2679 se
rect 4735 2672 4750 2693
tri 4735 2657 4750 2672 nw
rect 5069 2672 5084 2848
tri 5084 2841 5097 2854 nw
rect 5170 2773 5185 3001
tri 4707 2651 4713 2657 se
rect 4713 2651 4722 2657
rect 4707 2635 4722 2651
tri 4722 2644 4735 2657 nw
rect 4876 2649 4893 2663
rect 4925 2649 4942 2663
tri 5069 2657 5084 2672 ne
tri 5084 2657 5106 2679 sw
rect 4707 2599 4722 2607
rect 4788 2635 4848 2649
rect 4803 2625 4848 2635
rect 4803 2607 4831 2625
tri 4707 2584 4722 2599 ne
tri 4722 2584 4744 2606 sw
rect 4788 2597 4831 2607
rect 4846 2621 4848 2625
rect 4970 2635 5030 2649
tri 5084 2644 5097 2657 ne
rect 5097 2651 5106 2657
tri 5106 2651 5112 2657 sw
rect 4970 2625 5015 2635
rect 4846 2597 4920 2621
rect 4788 2593 4920 2597
tri 4920 2593 4948 2621 sw
rect 4970 2611 4972 2625
tri 4970 2609 4972 2611 ne
rect 4984 2607 5015 2625
rect 4984 2597 5030 2607
rect 5097 2636 5112 2651
tri 4722 2572 4734 2584 ne
rect 4734 2579 4744 2584
tri 4744 2579 4749 2584 sw
rect 4633 2233 4648 2461
rect 4734 2423 4749 2579
rect 4788 2537 4816 2593
tri 4908 2575 4926 2593 ne
rect 4926 2573 4948 2593
tri 4948 2573 4968 2593 sw
tri 4984 2579 5002 2597 ne
rect 4807 2503 4816 2537
rect 4850 2564 4892 2565
rect 4850 2530 4855 2564
rect 4885 2530 4892 2564
rect 4850 2521 4892 2530
rect 4926 2564 4968 2573
rect 4926 2530 4933 2564
rect 4963 2530 4968 2564
rect 4926 2525 4968 2530
rect 5002 2537 5030 2597
tri 5075 2584 5097 2606 se
rect 5097 2599 5112 2607
tri 5097 2584 5112 2599 nw
tri 5069 2578 5075 2584 se
rect 5075 2578 5084 2584
rect 4788 2493 4816 2503
tri 4816 2493 4840 2517 sw
rect 4788 2461 4830 2493
tri 4847 2485 4848 2486 sw
rect 4847 2461 4848 2485
tri 4850 2484 4887 2521 ne
rect 4887 2493 4892 2521
tri 4892 2493 4918 2519 sw
rect 5002 2503 5011 2537
rect 5002 2493 5030 2503
rect 4887 2484 4971 2493
tri 4887 2465 4906 2484 ne
rect 4906 2465 4971 2484
rect 4788 2439 4848 2461
rect 4970 2461 4971 2465
rect 4988 2461 5030 2493
rect 4970 2439 5030 2461
rect 4876 2423 4893 2437
rect 4925 2423 4942 2437
tri 4713 2387 4735 2409 se
rect 4735 2402 4750 2423
tri 4735 2387 4750 2402 nw
rect 5069 2402 5084 2578
tri 5084 2571 5097 2584 nw
rect 5170 2503 5185 2731
tri 4707 2381 4713 2387 se
rect 4713 2381 4722 2387
rect 4707 2365 4722 2381
tri 4722 2374 4735 2387 nw
rect 4876 2379 4893 2393
rect 4925 2379 4942 2393
tri 5069 2387 5084 2402 ne
tri 5084 2387 5106 2409 sw
rect 4707 2329 4722 2337
rect 4788 2365 4848 2379
rect 4803 2355 4848 2365
rect 4803 2337 4831 2355
tri 4707 2314 4722 2329 ne
tri 4722 2314 4744 2336 sw
rect 4788 2327 4831 2337
rect 4846 2351 4848 2355
rect 4970 2365 5030 2379
tri 5084 2374 5097 2387 ne
rect 5097 2381 5106 2387
tri 5106 2381 5112 2387 sw
rect 4970 2355 5015 2365
rect 4846 2327 4920 2351
rect 4788 2323 4920 2327
tri 4920 2323 4948 2351 sw
rect 4970 2341 4972 2355
tri 4970 2339 4972 2341 ne
rect 4984 2337 5015 2355
rect 4984 2327 5030 2337
rect 5097 2366 5112 2381
tri 4722 2302 4734 2314 ne
rect 4734 2309 4744 2314
tri 4744 2309 4749 2314 sw
rect 4633 1963 4648 2191
rect 4734 2201 4749 2309
rect 4788 2267 4816 2323
tri 4908 2305 4926 2323 ne
rect 4926 2303 4948 2323
tri 4948 2303 4968 2323 sw
tri 4984 2309 5002 2327 ne
rect 4807 2233 4816 2267
rect 4850 2294 4892 2295
rect 4850 2260 4855 2294
rect 4885 2260 4892 2294
rect 4850 2251 4892 2260
rect 4926 2294 4968 2303
rect 4926 2260 4933 2294
rect 4963 2260 4968 2294
rect 4926 2255 4968 2260
rect 5002 2267 5030 2327
tri 5075 2314 5097 2336 se
rect 5097 2329 5112 2337
tri 5097 2314 5112 2329 nw
tri 5069 2308 5075 2314 se
rect 5075 2308 5084 2314
rect 4788 2223 4816 2233
tri 4816 2223 4840 2247 sw
rect 4734 2153 4750 2201
rect 4788 2191 4830 2223
tri 4847 2215 4848 2216 sw
rect 4847 2191 4848 2215
tri 4850 2214 4887 2251 ne
rect 4887 2223 4892 2251
tri 4892 2223 4918 2249 sw
rect 5002 2233 5011 2267
rect 5002 2223 5030 2233
rect 4887 2214 4971 2223
tri 4887 2195 4906 2214 ne
rect 4906 2195 4971 2214
rect 4788 2169 4848 2191
rect 4970 2191 4971 2195
rect 4988 2191 5030 2223
rect 4970 2169 5030 2191
rect 4876 2153 4893 2167
rect 4925 2153 4942 2167
tri 4713 2117 4735 2139 se
rect 4735 2132 4750 2153
tri 4735 2117 4750 2132 nw
rect 5069 2132 5084 2308
tri 5084 2301 5097 2314 nw
rect 5170 2233 5185 2461
tri 4707 2111 4713 2117 se
rect 4713 2111 4722 2117
rect 4707 2095 4722 2111
tri 4722 2104 4735 2117 nw
rect 4876 2109 4893 2123
rect 4925 2109 4942 2123
tri 5069 2117 5084 2132 ne
tri 5084 2117 5106 2139 sw
rect 4707 2059 4722 2067
rect 4788 2095 4848 2109
rect 4803 2085 4848 2095
rect 4803 2067 4831 2085
tri 4707 2044 4722 2059 ne
tri 4722 2044 4744 2066 sw
rect 4788 2057 4831 2067
rect 4846 2081 4848 2085
rect 4970 2095 5030 2109
tri 5084 2104 5097 2117 ne
rect 5097 2111 5106 2117
tri 5106 2111 5112 2117 sw
rect 4970 2085 5015 2095
rect 4846 2057 4920 2081
rect 4788 2053 4920 2057
tri 4920 2053 4948 2081 sw
rect 4970 2071 4972 2085
tri 4970 2069 4972 2071 ne
rect 4984 2067 5015 2085
rect 4984 2057 5030 2067
rect 5097 2096 5112 2111
tri 4722 2032 4734 2044 ne
rect 4734 2039 4744 2044
tri 4744 2039 4749 2044 sw
rect 4633 1693 4648 1921
rect 4734 1883 4749 2039
rect 4788 1997 4816 2053
tri 4908 2035 4926 2053 ne
rect 4926 2033 4948 2053
tri 4948 2033 4968 2053 sw
tri 4984 2039 5002 2057 ne
rect 4807 1963 4816 1997
rect 4850 2024 4892 2025
rect 4850 1990 4855 2024
rect 4885 1990 4892 2024
rect 4850 1981 4892 1990
rect 4926 2024 4968 2033
rect 4926 1990 4933 2024
rect 4963 1990 4968 2024
rect 4926 1985 4968 1990
rect 5002 1997 5030 2057
tri 5075 2044 5097 2066 se
rect 5097 2059 5112 2067
tri 5097 2044 5112 2059 nw
tri 5069 2038 5075 2044 se
rect 5075 2038 5084 2044
rect 4788 1953 4816 1963
tri 4816 1953 4840 1977 sw
rect 4788 1921 4830 1953
tri 4847 1945 4848 1946 sw
rect 4847 1921 4848 1945
tri 4850 1944 4887 1981 ne
rect 4887 1953 4892 1981
tri 4892 1953 4918 1979 sw
rect 5002 1963 5011 1997
rect 5002 1953 5030 1963
rect 4887 1944 4971 1953
tri 4887 1925 4906 1944 ne
rect 4906 1925 4971 1944
rect 4788 1899 4848 1921
rect 4970 1921 4971 1925
rect 4988 1921 5030 1953
rect 4970 1899 5030 1921
rect 4876 1883 4893 1897
rect 4925 1883 4942 1897
tri 4713 1847 4735 1869 se
rect 4735 1862 4750 1883
tri 4735 1847 4750 1862 nw
rect 5069 1862 5084 2038
tri 5084 2031 5097 2044 nw
rect 5170 1963 5185 2191
tri 4707 1841 4713 1847 se
rect 4713 1841 4722 1847
rect 4707 1825 4722 1841
tri 4722 1834 4735 1847 nw
rect 4876 1839 4893 1853
rect 4925 1839 4942 1853
tri 5069 1847 5084 1862 ne
tri 5084 1847 5106 1869 sw
rect 4707 1789 4722 1797
rect 4788 1825 4848 1839
rect 4803 1815 4848 1825
rect 4803 1797 4831 1815
tri 4707 1774 4722 1789 ne
tri 4722 1774 4744 1796 sw
rect 4788 1787 4831 1797
rect 4846 1811 4848 1815
rect 4970 1825 5030 1839
tri 5084 1834 5097 1847 ne
rect 5097 1841 5106 1847
tri 5106 1841 5112 1847 sw
rect 4970 1815 5015 1825
rect 4846 1787 4920 1811
rect 4788 1783 4920 1787
tri 4920 1783 4948 1811 sw
rect 4970 1801 4972 1815
tri 4970 1799 4972 1801 ne
rect 4984 1797 5015 1815
rect 4984 1787 5030 1797
rect 5097 1826 5112 1841
tri 4722 1762 4734 1774 ne
rect 4734 1769 4744 1774
tri 4744 1769 4749 1774 sw
rect 4633 1423 4648 1651
rect 4734 1661 4749 1769
rect 4788 1727 4816 1783
tri 4908 1765 4926 1783 ne
rect 4926 1763 4948 1783
tri 4948 1763 4968 1783 sw
tri 4984 1769 5002 1787 ne
rect 4807 1693 4816 1727
rect 4850 1754 4892 1755
rect 4850 1720 4855 1754
rect 4885 1720 4892 1754
rect 4850 1711 4892 1720
rect 4926 1754 4968 1763
rect 4926 1720 4933 1754
rect 4963 1720 4968 1754
rect 4926 1715 4968 1720
rect 5002 1727 5030 1787
tri 5075 1774 5097 1796 se
rect 5097 1789 5112 1797
tri 5097 1774 5112 1789 nw
tri 5069 1768 5075 1774 se
rect 5075 1768 5084 1774
rect 4788 1683 4816 1693
tri 4816 1683 4840 1707 sw
rect 4734 1613 4750 1661
rect 4788 1651 4830 1683
tri 4847 1675 4848 1676 sw
rect 4847 1651 4848 1675
tri 4850 1674 4887 1711 ne
rect 4887 1683 4892 1711
tri 4892 1683 4918 1709 sw
rect 5002 1693 5011 1727
rect 5002 1683 5030 1693
rect 4887 1674 4971 1683
tri 4887 1655 4906 1674 ne
rect 4906 1655 4971 1674
rect 4788 1629 4848 1651
rect 4970 1651 4971 1655
rect 4988 1651 5030 1683
rect 4970 1629 5030 1651
rect 4876 1613 4893 1627
rect 4925 1613 4942 1627
tri 4713 1577 4735 1599 se
rect 4735 1592 4750 1613
tri 4735 1577 4750 1592 nw
rect 5069 1592 5084 1768
tri 5084 1761 5097 1774 nw
rect 5170 1693 5185 1921
tri 4707 1571 4713 1577 se
rect 4713 1571 4722 1577
rect 4707 1555 4722 1571
tri 4722 1564 4735 1577 nw
rect 4876 1569 4893 1583
rect 4925 1569 4942 1583
tri 5069 1577 5084 1592 ne
tri 5084 1577 5106 1599 sw
rect 4707 1519 4722 1527
rect 4788 1555 4848 1569
rect 4803 1545 4848 1555
rect 4803 1527 4831 1545
tri 4707 1504 4722 1519 ne
tri 4722 1504 4744 1526 sw
rect 4788 1517 4831 1527
rect 4846 1541 4848 1545
rect 4970 1555 5030 1569
tri 5084 1564 5097 1577 ne
rect 5097 1571 5106 1577
tri 5106 1571 5112 1577 sw
rect 4970 1545 5015 1555
rect 4846 1517 4920 1541
rect 4788 1513 4920 1517
tri 4920 1513 4948 1541 sw
rect 4970 1531 4972 1545
tri 4970 1529 4972 1531 ne
rect 4984 1527 5015 1545
rect 4984 1517 5030 1527
rect 5097 1556 5112 1571
tri 4722 1492 4734 1504 ne
rect 4734 1499 4744 1504
tri 4744 1499 4749 1504 sw
rect 4633 1153 4648 1381
rect 4734 1343 4749 1499
rect 4788 1457 4816 1513
tri 4908 1495 4926 1513 ne
rect 4926 1493 4948 1513
tri 4948 1493 4968 1513 sw
tri 4984 1499 5002 1517 ne
rect 4807 1423 4816 1457
rect 4850 1484 4892 1485
rect 4850 1450 4855 1484
rect 4885 1450 4892 1484
rect 4850 1441 4892 1450
rect 4926 1484 4968 1493
rect 4926 1450 4933 1484
rect 4963 1450 4968 1484
rect 4926 1445 4968 1450
rect 5002 1457 5030 1517
tri 5075 1504 5097 1526 se
rect 5097 1519 5112 1527
tri 5097 1504 5112 1519 nw
tri 5069 1498 5075 1504 se
rect 5075 1498 5084 1504
rect 4788 1413 4816 1423
tri 4816 1413 4840 1437 sw
rect 4788 1381 4830 1413
tri 4847 1405 4848 1406 sw
rect 4847 1381 4848 1405
tri 4850 1404 4887 1441 ne
rect 4887 1413 4892 1441
tri 4892 1413 4918 1439 sw
rect 5002 1423 5011 1457
rect 5002 1413 5030 1423
rect 4887 1404 4971 1413
tri 4887 1385 4906 1404 ne
rect 4906 1385 4971 1404
rect 4788 1359 4848 1381
rect 4970 1381 4971 1385
rect 4988 1381 5030 1413
rect 4970 1359 5030 1381
rect 4876 1343 4893 1357
rect 4925 1343 4942 1357
tri 4713 1307 4735 1329 se
rect 4735 1322 4750 1343
tri 4735 1307 4750 1322 nw
rect 5069 1322 5084 1498
tri 5084 1491 5097 1504 nw
rect 5170 1423 5185 1651
tri 4707 1301 4713 1307 se
rect 4713 1301 4722 1307
rect 4707 1285 4722 1301
tri 4722 1294 4735 1307 nw
rect 4876 1299 4893 1313
rect 4925 1299 4942 1313
tri 5069 1307 5084 1322 ne
tri 5084 1307 5106 1329 sw
rect 4707 1249 4722 1257
rect 4788 1285 4848 1299
rect 4803 1275 4848 1285
rect 4803 1257 4831 1275
tri 4707 1234 4722 1249 ne
tri 4722 1234 4744 1256 sw
rect 4788 1247 4831 1257
rect 4846 1271 4848 1275
rect 4970 1285 5030 1299
tri 5084 1294 5097 1307 ne
rect 5097 1301 5106 1307
tri 5106 1301 5112 1307 sw
rect 4970 1275 5015 1285
rect 4846 1247 4920 1271
rect 4788 1243 4920 1247
tri 4920 1243 4948 1271 sw
rect 4970 1261 4972 1275
tri 4970 1259 4972 1261 ne
rect 4984 1257 5015 1275
rect 4984 1247 5030 1257
rect 5097 1286 5112 1301
tri 4722 1222 4734 1234 ne
rect 4734 1229 4744 1234
tri 4744 1229 4749 1234 sw
rect 4633 883 4648 1111
rect 4734 1121 4749 1229
rect 4788 1187 4816 1243
tri 4908 1225 4926 1243 ne
rect 4926 1223 4948 1243
tri 4948 1223 4968 1243 sw
tri 4984 1229 5002 1247 ne
rect 4807 1153 4816 1187
rect 4850 1214 4892 1215
rect 4850 1180 4855 1214
rect 4885 1180 4892 1214
rect 4850 1171 4892 1180
rect 4926 1214 4968 1223
rect 4926 1180 4933 1214
rect 4963 1180 4968 1214
rect 4926 1175 4968 1180
rect 5002 1187 5030 1247
tri 5075 1234 5097 1256 se
rect 5097 1249 5112 1257
tri 5097 1234 5112 1249 nw
tri 5069 1228 5075 1234 se
rect 5075 1228 5084 1234
rect 4788 1143 4816 1153
tri 4816 1143 4840 1167 sw
rect 4734 1073 4750 1121
rect 4788 1111 4830 1143
tri 4847 1135 4848 1136 sw
rect 4847 1111 4848 1135
tri 4850 1134 4887 1171 ne
rect 4887 1143 4892 1171
tri 4892 1143 4918 1169 sw
rect 5002 1153 5011 1187
rect 5002 1143 5030 1153
rect 4887 1134 4971 1143
tri 4887 1115 4906 1134 ne
rect 4906 1115 4971 1134
rect 4788 1089 4848 1111
rect 4970 1111 4971 1115
rect 4988 1111 5030 1143
rect 4970 1089 5030 1111
rect 4876 1073 4893 1087
rect 4925 1073 4942 1087
tri 4713 1037 4735 1059 se
rect 4735 1052 4750 1073
tri 4735 1037 4750 1052 nw
rect 5069 1052 5084 1228
tri 5084 1221 5097 1234 nw
rect 5170 1153 5185 1381
tri 4707 1031 4713 1037 se
rect 4713 1031 4722 1037
rect 4707 1015 4722 1031
tri 4722 1024 4735 1037 nw
rect 4876 1029 4893 1043
rect 4925 1029 4942 1043
tri 5069 1037 5084 1052 ne
tri 5084 1037 5106 1059 sw
rect 4707 979 4722 987
rect 4788 1015 4848 1029
rect 4803 1005 4848 1015
rect 4803 987 4831 1005
tri 4707 964 4722 979 ne
tri 4722 964 4744 986 sw
rect 4788 977 4831 987
rect 4846 1001 4848 1005
rect 4970 1015 5030 1029
tri 5084 1024 5097 1037 ne
rect 5097 1031 5106 1037
tri 5106 1031 5112 1037 sw
rect 4970 1005 5015 1015
rect 4846 977 4920 1001
rect 4788 973 4920 977
tri 4920 973 4948 1001 sw
rect 4970 991 4972 1005
tri 4970 989 4972 991 ne
rect 4984 987 5015 1005
rect 4984 977 5030 987
rect 5097 1016 5112 1031
tri 4722 952 4734 964 ne
rect 4734 959 4744 964
tri 4744 959 4749 964 sw
rect 4633 613 4648 841
rect 4734 803 4749 959
rect 4788 917 4816 973
tri 4908 955 4926 973 ne
rect 4926 953 4948 973
tri 4948 953 4968 973 sw
tri 4984 959 5002 977 ne
rect 4807 883 4816 917
rect 4850 944 4892 945
rect 4850 910 4855 944
rect 4885 910 4892 944
rect 4850 901 4892 910
rect 4926 944 4968 953
rect 4926 910 4933 944
rect 4963 910 4968 944
rect 4926 905 4968 910
rect 5002 917 5030 977
tri 5075 964 5097 986 se
rect 5097 979 5112 987
tri 5097 964 5112 979 nw
tri 5069 958 5075 964 se
rect 5075 958 5084 964
rect 4788 873 4816 883
tri 4816 873 4840 897 sw
rect 4788 841 4830 873
tri 4847 865 4848 866 sw
rect 4847 841 4848 865
tri 4850 864 4887 901 ne
rect 4887 873 4892 901
tri 4892 873 4918 899 sw
rect 5002 883 5011 917
rect 5002 873 5030 883
rect 4887 864 4971 873
tri 4887 845 4906 864 ne
rect 4906 845 4971 864
rect 4788 819 4848 841
rect 4970 841 4971 845
rect 4988 841 5030 873
rect 4970 819 5030 841
rect 4876 803 4893 817
rect 4925 803 4942 817
tri 4713 767 4735 789 se
rect 4735 782 4750 803
tri 4735 767 4750 782 nw
rect 5069 782 5084 958
tri 5084 951 5097 964 nw
rect 5170 883 5185 1111
tri 4707 761 4713 767 se
rect 4713 761 4722 767
rect 4707 745 4722 761
tri 4722 754 4735 767 nw
rect 4876 759 4893 773
rect 4925 759 4942 773
tri 5069 767 5084 782 ne
tri 5084 767 5106 789 sw
rect 4707 709 4722 717
rect 4788 745 4848 759
rect 4803 735 4848 745
rect 4803 717 4831 735
tri 4707 694 4722 709 ne
tri 4722 694 4744 716 sw
rect 4788 707 4831 717
rect 4846 731 4848 735
rect 4970 745 5030 759
tri 5084 754 5097 767 ne
rect 5097 761 5106 767
tri 5106 761 5112 767 sw
rect 4970 735 5015 745
rect 4846 707 4920 731
rect 4788 703 4920 707
tri 4920 703 4948 731 sw
rect 4970 721 4972 735
tri 4970 719 4972 721 ne
rect 4984 717 5015 735
rect 4984 707 5030 717
rect 5097 746 5112 761
tri 4722 682 4734 694 ne
rect 4734 689 4744 694
tri 4744 689 4749 694 sw
rect 4633 343 4648 571
rect 4734 581 4749 689
rect 4788 647 4816 703
tri 4908 685 4926 703 ne
rect 4926 683 4948 703
tri 4948 683 4968 703 sw
tri 4984 689 5002 707 ne
rect 4807 613 4816 647
rect 4850 674 4892 675
rect 4850 640 4855 674
rect 4885 640 4892 674
rect 4850 631 4892 640
rect 4926 674 4968 683
rect 4926 640 4933 674
rect 4963 640 4968 674
rect 4926 635 4968 640
rect 5002 647 5030 707
tri 5075 694 5097 716 se
rect 5097 709 5112 717
tri 5097 694 5112 709 nw
tri 5069 688 5075 694 se
rect 5075 688 5084 694
rect 4788 603 4816 613
tri 4816 603 4840 627 sw
rect 4734 533 4750 581
rect 4788 571 4830 603
tri 4847 595 4848 596 sw
rect 4847 571 4848 595
tri 4850 594 4887 631 ne
rect 4887 603 4892 631
tri 4892 603 4918 629 sw
rect 5002 613 5011 647
rect 5002 603 5030 613
rect 4887 594 4971 603
tri 4887 575 4906 594 ne
rect 4906 575 4971 594
rect 4788 549 4848 571
rect 4970 571 4971 575
rect 4988 571 5030 603
rect 4970 549 5030 571
rect 4876 533 4893 547
rect 4925 533 4942 547
tri 4713 497 4735 519 se
rect 4735 512 4750 533
tri 4735 497 4750 512 nw
rect 5069 512 5084 688
tri 5084 681 5097 694 nw
rect 5170 613 5185 841
tri 4707 491 4713 497 se
rect 4713 491 4722 497
rect 4707 475 4722 491
tri 4722 484 4735 497 nw
rect 4876 489 4893 503
rect 4925 489 4942 503
tri 5069 497 5084 512 ne
tri 5084 497 5106 519 sw
rect 4707 439 4722 447
rect 4788 475 4848 489
rect 4803 465 4848 475
rect 4803 447 4831 465
tri 4707 424 4722 439 ne
tri 4722 424 4744 446 sw
rect 4788 437 4831 447
rect 4846 461 4848 465
rect 4970 475 5030 489
tri 5084 484 5097 497 ne
rect 5097 491 5106 497
tri 5106 491 5112 497 sw
rect 4970 465 5015 475
rect 4846 437 4920 461
rect 4788 433 4920 437
tri 4920 433 4948 461 sw
rect 4970 451 4972 465
tri 4970 449 4972 451 ne
rect 4984 447 5015 465
rect 4984 437 5030 447
rect 5097 476 5112 491
tri 4722 412 4734 424 ne
rect 4734 419 4744 424
tri 4744 419 4749 424 sw
rect 4633 73 4648 301
rect 4734 263 4749 419
rect 4788 377 4816 433
tri 4908 415 4926 433 ne
rect 4926 413 4948 433
tri 4948 413 4968 433 sw
tri 4984 419 5002 437 ne
rect 4807 343 4816 377
rect 4850 404 4892 405
rect 4850 370 4855 404
rect 4885 370 4892 404
rect 4850 361 4892 370
rect 4926 404 4968 413
rect 4926 370 4933 404
rect 4963 370 4968 404
rect 4926 365 4968 370
rect 5002 377 5030 437
tri 5075 424 5097 446 se
rect 5097 439 5112 447
tri 5097 424 5112 439 nw
tri 5069 418 5075 424 se
rect 5075 418 5084 424
rect 4788 333 4816 343
tri 4816 333 4840 357 sw
rect 4788 301 4830 333
tri 4847 325 4848 326 sw
rect 4847 301 4848 325
tri 4850 324 4887 361 ne
rect 4887 333 4892 361
tri 4892 333 4918 359 sw
rect 5002 343 5011 377
rect 5002 333 5030 343
rect 4887 324 4971 333
tri 4887 305 4906 324 ne
rect 4906 305 4971 324
rect 4788 279 4848 301
rect 4970 301 4971 305
rect 4988 301 5030 333
rect 4970 279 5030 301
rect 4876 263 4893 277
rect 4925 263 4942 277
tri 4713 227 4735 249 se
rect 4735 242 4750 263
tri 4735 227 4750 242 nw
rect 5069 242 5084 418
tri 5084 411 5097 424 nw
rect 5170 343 5185 571
tri 4707 221 4713 227 se
rect 4713 221 4722 227
rect 4707 205 4722 221
tri 4722 214 4735 227 nw
rect 4876 219 4893 233
rect 4925 219 4942 233
tri 5069 227 5084 242 ne
tri 5084 227 5106 249 sw
rect 4707 169 4722 177
rect 4788 205 4848 219
rect 4803 195 4848 205
rect 4803 177 4831 195
tri 4707 154 4722 169 ne
tri 4722 154 4744 176 sw
rect 4788 167 4831 177
rect 4846 191 4848 195
rect 4970 205 5030 219
tri 5084 214 5097 227 ne
rect 5097 221 5106 227
tri 5106 221 5112 227 sw
rect 4970 195 5015 205
rect 4846 167 4920 191
rect 4788 163 4920 167
tri 4920 163 4948 191 sw
rect 4970 181 4972 195
tri 4970 179 4972 181 ne
rect 4984 177 5015 195
rect 4984 167 5030 177
rect 5097 206 5112 221
tri 4722 142 4734 154 ne
rect 4734 149 4744 154
tri 4744 149 4749 154 sw
rect 4633 -55 4648 31
rect 4734 -55 4749 149
rect 4788 107 4816 163
tri 4908 145 4926 163 ne
rect 4926 143 4948 163
tri 4948 143 4968 163 sw
tri 4984 149 5002 167 ne
rect 4807 73 4816 107
rect 4850 134 4892 135
rect 4850 100 4855 134
rect 4885 100 4892 134
rect 4850 91 4892 100
rect 4926 134 4968 143
rect 4926 100 4933 134
rect 4963 100 4968 134
rect 4926 95 4968 100
rect 5002 107 5030 167
tri 5075 154 5097 176 se
rect 5097 169 5112 177
tri 5097 154 5112 169 nw
tri 5069 148 5075 154 se
rect 5075 148 5084 154
rect 4788 63 4816 73
tri 4816 63 4840 87 sw
rect 4788 31 4830 63
tri 4847 55 4848 56 sw
rect 4847 31 4848 55
tri 4850 54 4887 91 ne
rect 4887 63 4892 91
tri 4892 63 4918 89 sw
rect 5002 73 5011 107
rect 5002 63 5030 73
rect 4887 54 4971 63
tri 4887 35 4906 54 ne
rect 4906 35 4971 54
rect 4788 9 4848 31
rect 4970 31 4971 35
rect 4988 31 5030 63
rect 4970 9 5030 31
rect 4876 -7 4893 7
rect 4925 -7 4942 7
rect 5069 -55 5084 148
tri 5084 141 5097 154 nw
rect 5170 73 5185 301
rect 5170 -55 5185 31
rect 5213 4123 5228 4361
tri 5293 4277 5315 4299 se
rect 5315 4292 5330 4361
tri 5315 4277 5330 4292 nw
rect 5649 4292 5664 4361
tri 5287 4271 5293 4277 se
rect 5293 4271 5302 4277
rect 5287 4255 5302 4271
tri 5302 4264 5315 4277 nw
rect 5456 4269 5473 4283
rect 5505 4269 5522 4283
tri 5649 4277 5664 4292 ne
tri 5664 4277 5686 4299 sw
rect 5287 4219 5302 4227
rect 5368 4255 5428 4269
rect 5383 4245 5428 4255
rect 5383 4227 5411 4245
tri 5287 4204 5302 4219 ne
tri 5302 4204 5324 4226 sw
rect 5368 4217 5411 4227
rect 5426 4241 5428 4245
rect 5550 4255 5610 4269
tri 5664 4264 5677 4277 ne
rect 5677 4271 5686 4277
tri 5686 4271 5692 4277 sw
rect 5550 4245 5595 4255
rect 5426 4217 5500 4241
rect 5368 4213 5500 4217
tri 5500 4213 5528 4241 sw
rect 5550 4231 5552 4245
tri 5550 4229 5552 4231 ne
rect 5564 4227 5595 4245
rect 5564 4217 5610 4227
rect 5677 4256 5692 4271
tri 5302 4192 5314 4204 ne
rect 5314 4199 5324 4204
tri 5324 4199 5329 4204 sw
rect 5213 3853 5228 4081
rect 5314 4043 5329 4199
rect 5368 4157 5396 4213
tri 5488 4195 5506 4213 ne
rect 5506 4193 5528 4213
tri 5528 4193 5548 4213 sw
tri 5564 4199 5582 4217 ne
rect 5387 4123 5396 4157
rect 5430 4184 5472 4185
rect 5430 4150 5435 4184
rect 5465 4150 5472 4184
rect 5430 4141 5472 4150
rect 5506 4184 5548 4193
rect 5506 4150 5513 4184
rect 5543 4150 5548 4184
rect 5506 4145 5548 4150
rect 5582 4157 5610 4217
tri 5655 4204 5677 4226 se
rect 5677 4219 5692 4227
tri 5677 4204 5692 4219 nw
tri 5649 4198 5655 4204 se
rect 5655 4198 5664 4204
rect 5368 4113 5396 4123
tri 5396 4113 5420 4137 sw
rect 5368 4081 5410 4113
tri 5427 4105 5428 4106 sw
rect 5427 4081 5428 4105
tri 5430 4104 5467 4141 ne
rect 5467 4113 5472 4141
tri 5472 4113 5498 4139 sw
rect 5582 4123 5591 4157
rect 5582 4113 5610 4123
rect 5467 4104 5551 4113
tri 5467 4085 5486 4104 ne
rect 5486 4085 5551 4104
rect 5368 4059 5428 4081
rect 5550 4081 5551 4085
rect 5568 4081 5610 4113
rect 5550 4059 5610 4081
rect 5456 4043 5473 4057
rect 5505 4043 5522 4057
tri 5293 4007 5315 4029 se
rect 5315 4022 5330 4043
tri 5315 4007 5330 4022 nw
rect 5649 4022 5664 4198
tri 5664 4191 5677 4204 nw
rect 5750 4123 5765 4361
tri 5287 4001 5293 4007 se
rect 5293 4001 5302 4007
rect 5287 3985 5302 4001
tri 5302 3994 5315 4007 nw
rect 5456 3999 5473 4013
rect 5505 3999 5522 4013
tri 5649 4007 5664 4022 ne
tri 5664 4007 5686 4029 sw
rect 5287 3949 5302 3957
rect 5368 3985 5428 3999
rect 5383 3975 5428 3985
rect 5383 3957 5411 3975
tri 5287 3934 5302 3949 ne
tri 5302 3934 5324 3956 sw
rect 5368 3947 5411 3957
rect 5426 3971 5428 3975
rect 5550 3985 5610 3999
tri 5664 3994 5677 4007 ne
rect 5677 4001 5686 4007
tri 5686 4001 5692 4007 sw
rect 5550 3975 5595 3985
rect 5426 3947 5500 3971
rect 5368 3943 5500 3947
tri 5500 3943 5528 3971 sw
rect 5550 3961 5552 3975
tri 5550 3959 5552 3961 ne
rect 5564 3957 5595 3975
rect 5564 3947 5610 3957
rect 5677 3986 5692 4001
tri 5302 3922 5314 3934 ne
rect 5314 3929 5324 3934
tri 5324 3929 5329 3934 sw
rect 5213 3583 5228 3811
rect 5314 3821 5329 3929
rect 5368 3887 5396 3943
tri 5488 3925 5506 3943 ne
rect 5506 3923 5528 3943
tri 5528 3923 5548 3943 sw
tri 5564 3929 5582 3947 ne
rect 5387 3853 5396 3887
rect 5430 3914 5472 3915
rect 5430 3880 5435 3914
rect 5465 3880 5472 3914
rect 5430 3871 5472 3880
rect 5506 3914 5548 3923
rect 5506 3880 5513 3914
rect 5543 3880 5548 3914
rect 5506 3875 5548 3880
rect 5582 3887 5610 3947
tri 5655 3934 5677 3956 se
rect 5677 3949 5692 3957
tri 5677 3934 5692 3949 nw
tri 5649 3928 5655 3934 se
rect 5655 3928 5664 3934
rect 5368 3843 5396 3853
tri 5396 3843 5420 3867 sw
rect 5314 3773 5330 3821
rect 5368 3811 5410 3843
tri 5427 3835 5428 3836 sw
rect 5427 3811 5428 3835
tri 5430 3834 5467 3871 ne
rect 5467 3843 5472 3871
tri 5472 3843 5498 3869 sw
rect 5582 3853 5591 3887
rect 5582 3843 5610 3853
rect 5467 3834 5551 3843
tri 5467 3815 5486 3834 ne
rect 5486 3815 5551 3834
rect 5368 3789 5428 3811
rect 5550 3811 5551 3815
rect 5568 3811 5610 3843
rect 5550 3789 5610 3811
rect 5456 3773 5473 3787
rect 5505 3773 5522 3787
tri 5293 3737 5315 3759 se
rect 5315 3752 5330 3773
tri 5315 3737 5330 3752 nw
rect 5649 3752 5664 3928
tri 5664 3921 5677 3934 nw
rect 5750 3853 5765 4081
tri 5287 3731 5293 3737 se
rect 5293 3731 5302 3737
rect 5287 3715 5302 3731
tri 5302 3724 5315 3737 nw
rect 5456 3729 5473 3743
rect 5505 3729 5522 3743
tri 5649 3737 5664 3752 ne
tri 5664 3737 5686 3759 sw
rect 5287 3679 5302 3687
rect 5368 3715 5428 3729
rect 5383 3705 5428 3715
rect 5383 3687 5411 3705
tri 5287 3664 5302 3679 ne
tri 5302 3664 5324 3686 sw
rect 5368 3677 5411 3687
rect 5426 3701 5428 3705
rect 5550 3715 5610 3729
tri 5664 3724 5677 3737 ne
rect 5677 3731 5686 3737
tri 5686 3731 5692 3737 sw
rect 5550 3705 5595 3715
rect 5426 3677 5500 3701
rect 5368 3673 5500 3677
tri 5500 3673 5528 3701 sw
rect 5550 3691 5552 3705
tri 5550 3689 5552 3691 ne
rect 5564 3687 5595 3705
rect 5564 3677 5610 3687
rect 5677 3716 5692 3731
tri 5302 3652 5314 3664 ne
rect 5314 3659 5324 3664
tri 5324 3659 5329 3664 sw
rect 5213 3313 5228 3541
rect 5314 3503 5329 3659
rect 5368 3617 5396 3673
tri 5488 3655 5506 3673 ne
rect 5506 3653 5528 3673
tri 5528 3653 5548 3673 sw
tri 5564 3659 5582 3677 ne
rect 5387 3583 5396 3617
rect 5430 3644 5472 3645
rect 5430 3610 5435 3644
rect 5465 3610 5472 3644
rect 5430 3601 5472 3610
rect 5506 3644 5548 3653
rect 5506 3610 5513 3644
rect 5543 3610 5548 3644
rect 5506 3605 5548 3610
rect 5582 3617 5610 3677
tri 5655 3664 5677 3686 se
rect 5677 3679 5692 3687
tri 5677 3664 5692 3679 nw
tri 5649 3658 5655 3664 se
rect 5655 3658 5664 3664
rect 5368 3573 5396 3583
tri 5396 3573 5420 3597 sw
rect 5368 3541 5410 3573
tri 5427 3565 5428 3566 sw
rect 5427 3541 5428 3565
tri 5430 3564 5467 3601 ne
rect 5467 3573 5472 3601
tri 5472 3573 5498 3599 sw
rect 5582 3583 5591 3617
rect 5582 3573 5610 3583
rect 5467 3564 5551 3573
tri 5467 3545 5486 3564 ne
rect 5486 3545 5551 3564
rect 5368 3519 5428 3541
rect 5550 3541 5551 3545
rect 5568 3541 5610 3573
rect 5550 3519 5610 3541
rect 5456 3503 5473 3517
rect 5505 3503 5522 3517
tri 5293 3467 5315 3489 se
rect 5315 3482 5330 3503
tri 5315 3467 5330 3482 nw
rect 5649 3482 5664 3658
tri 5664 3651 5677 3664 nw
rect 5750 3583 5765 3811
tri 5287 3461 5293 3467 se
rect 5293 3461 5302 3467
rect 5287 3445 5302 3461
tri 5302 3454 5315 3467 nw
rect 5456 3459 5473 3473
rect 5505 3459 5522 3473
tri 5649 3467 5664 3482 ne
tri 5664 3467 5686 3489 sw
rect 5287 3409 5302 3417
rect 5368 3445 5428 3459
rect 5383 3435 5428 3445
rect 5383 3417 5411 3435
tri 5287 3394 5302 3409 ne
tri 5302 3394 5324 3416 sw
rect 5368 3407 5411 3417
rect 5426 3431 5428 3435
rect 5550 3445 5610 3459
tri 5664 3454 5677 3467 ne
rect 5677 3461 5686 3467
tri 5686 3461 5692 3467 sw
rect 5550 3435 5595 3445
rect 5426 3407 5500 3431
rect 5368 3403 5500 3407
tri 5500 3403 5528 3431 sw
rect 5550 3421 5552 3435
tri 5550 3419 5552 3421 ne
rect 5564 3417 5595 3435
rect 5564 3407 5610 3417
rect 5677 3446 5692 3461
tri 5302 3382 5314 3394 ne
rect 5314 3389 5324 3394
tri 5324 3389 5329 3394 sw
rect 5213 3043 5228 3271
rect 5314 3281 5329 3389
rect 5368 3347 5396 3403
tri 5488 3385 5506 3403 ne
rect 5506 3383 5528 3403
tri 5528 3383 5548 3403 sw
tri 5564 3389 5582 3407 ne
rect 5387 3313 5396 3347
rect 5430 3374 5472 3375
rect 5430 3340 5435 3374
rect 5465 3340 5472 3374
rect 5430 3331 5472 3340
rect 5506 3374 5548 3383
rect 5506 3340 5513 3374
rect 5543 3340 5548 3374
rect 5506 3335 5548 3340
rect 5582 3347 5610 3407
tri 5655 3394 5677 3416 se
rect 5677 3409 5692 3417
tri 5677 3394 5692 3409 nw
tri 5649 3388 5655 3394 se
rect 5655 3388 5664 3394
rect 5368 3303 5396 3313
tri 5396 3303 5420 3327 sw
rect 5314 3233 5330 3281
rect 5368 3271 5410 3303
tri 5427 3295 5428 3296 sw
rect 5427 3271 5428 3295
tri 5430 3294 5467 3331 ne
rect 5467 3303 5472 3331
tri 5472 3303 5498 3329 sw
rect 5582 3313 5591 3347
rect 5582 3303 5610 3313
rect 5467 3294 5551 3303
tri 5467 3275 5486 3294 ne
rect 5486 3275 5551 3294
rect 5368 3249 5428 3271
rect 5550 3271 5551 3275
rect 5568 3271 5610 3303
rect 5550 3249 5610 3271
rect 5456 3233 5473 3247
rect 5505 3233 5522 3247
tri 5293 3197 5315 3219 se
rect 5315 3212 5330 3233
tri 5315 3197 5330 3212 nw
rect 5649 3212 5664 3388
tri 5664 3381 5677 3394 nw
rect 5750 3313 5765 3541
tri 5287 3191 5293 3197 se
rect 5293 3191 5302 3197
rect 5287 3175 5302 3191
tri 5302 3184 5315 3197 nw
rect 5456 3189 5473 3203
rect 5505 3189 5522 3203
tri 5649 3197 5664 3212 ne
tri 5664 3197 5686 3219 sw
rect 5287 3139 5302 3147
rect 5368 3175 5428 3189
rect 5383 3165 5428 3175
rect 5383 3147 5411 3165
tri 5287 3124 5302 3139 ne
tri 5302 3124 5324 3146 sw
rect 5368 3137 5411 3147
rect 5426 3161 5428 3165
rect 5550 3175 5610 3189
tri 5664 3184 5677 3197 ne
rect 5677 3191 5686 3197
tri 5686 3191 5692 3197 sw
rect 5550 3165 5595 3175
rect 5426 3137 5500 3161
rect 5368 3133 5500 3137
tri 5500 3133 5528 3161 sw
rect 5550 3151 5552 3165
tri 5550 3149 5552 3151 ne
rect 5564 3147 5595 3165
rect 5564 3137 5610 3147
rect 5677 3176 5692 3191
tri 5302 3112 5314 3124 ne
rect 5314 3119 5324 3124
tri 5324 3119 5329 3124 sw
rect 5213 2773 5228 3001
rect 5314 2963 5329 3119
rect 5368 3077 5396 3133
tri 5488 3115 5506 3133 ne
rect 5506 3113 5528 3133
tri 5528 3113 5548 3133 sw
tri 5564 3119 5582 3137 ne
rect 5387 3043 5396 3077
rect 5430 3104 5472 3105
rect 5430 3070 5435 3104
rect 5465 3070 5472 3104
rect 5430 3061 5472 3070
rect 5506 3104 5548 3113
rect 5506 3070 5513 3104
rect 5543 3070 5548 3104
rect 5506 3065 5548 3070
rect 5582 3077 5610 3137
tri 5655 3124 5677 3146 se
rect 5677 3139 5692 3147
tri 5677 3124 5692 3139 nw
tri 5649 3118 5655 3124 se
rect 5655 3118 5664 3124
rect 5368 3033 5396 3043
tri 5396 3033 5420 3057 sw
rect 5368 3001 5410 3033
tri 5427 3025 5428 3026 sw
rect 5427 3001 5428 3025
tri 5430 3024 5467 3061 ne
rect 5467 3033 5472 3061
tri 5472 3033 5498 3059 sw
rect 5582 3043 5591 3077
rect 5582 3033 5610 3043
rect 5467 3024 5551 3033
tri 5467 3005 5486 3024 ne
rect 5486 3005 5551 3024
rect 5368 2979 5428 3001
rect 5550 3001 5551 3005
rect 5568 3001 5610 3033
rect 5550 2979 5610 3001
rect 5456 2963 5473 2977
rect 5505 2963 5522 2977
tri 5293 2927 5315 2949 se
rect 5315 2942 5330 2963
tri 5315 2927 5330 2942 nw
rect 5649 2942 5664 3118
tri 5664 3111 5677 3124 nw
rect 5750 3043 5765 3271
tri 5287 2921 5293 2927 se
rect 5293 2921 5302 2927
rect 5287 2905 5302 2921
tri 5302 2914 5315 2927 nw
rect 5456 2919 5473 2933
rect 5505 2919 5522 2933
tri 5649 2927 5664 2942 ne
tri 5664 2927 5686 2949 sw
rect 5287 2869 5302 2877
rect 5368 2905 5428 2919
rect 5383 2895 5428 2905
rect 5383 2877 5411 2895
tri 5287 2854 5302 2869 ne
tri 5302 2854 5324 2876 sw
rect 5368 2867 5411 2877
rect 5426 2891 5428 2895
rect 5550 2905 5610 2919
tri 5664 2914 5677 2927 ne
rect 5677 2921 5686 2927
tri 5686 2921 5692 2927 sw
rect 5550 2895 5595 2905
rect 5426 2867 5500 2891
rect 5368 2863 5500 2867
tri 5500 2863 5528 2891 sw
rect 5550 2881 5552 2895
tri 5550 2879 5552 2881 ne
rect 5564 2877 5595 2895
rect 5564 2867 5610 2877
rect 5677 2906 5692 2921
tri 5302 2842 5314 2854 ne
rect 5314 2849 5324 2854
tri 5324 2849 5329 2854 sw
rect 5213 2503 5228 2731
rect 5314 2741 5329 2849
rect 5368 2807 5396 2863
tri 5488 2845 5506 2863 ne
rect 5506 2843 5528 2863
tri 5528 2843 5548 2863 sw
tri 5564 2849 5582 2867 ne
rect 5387 2773 5396 2807
rect 5430 2834 5472 2835
rect 5430 2800 5435 2834
rect 5465 2800 5472 2834
rect 5430 2791 5472 2800
rect 5506 2834 5548 2843
rect 5506 2800 5513 2834
rect 5543 2800 5548 2834
rect 5506 2795 5548 2800
rect 5582 2807 5610 2867
tri 5655 2854 5677 2876 se
rect 5677 2869 5692 2877
tri 5677 2854 5692 2869 nw
tri 5649 2848 5655 2854 se
rect 5655 2848 5664 2854
rect 5368 2763 5396 2773
tri 5396 2763 5420 2787 sw
rect 5314 2693 5330 2741
rect 5368 2731 5410 2763
tri 5427 2755 5428 2756 sw
rect 5427 2731 5428 2755
tri 5430 2754 5467 2791 ne
rect 5467 2763 5472 2791
tri 5472 2763 5498 2789 sw
rect 5582 2773 5591 2807
rect 5582 2763 5610 2773
rect 5467 2754 5551 2763
tri 5467 2735 5486 2754 ne
rect 5486 2735 5551 2754
rect 5368 2709 5428 2731
rect 5550 2731 5551 2735
rect 5568 2731 5610 2763
rect 5550 2709 5610 2731
rect 5456 2693 5473 2707
rect 5505 2693 5522 2707
tri 5293 2657 5315 2679 se
rect 5315 2672 5330 2693
tri 5315 2657 5330 2672 nw
rect 5649 2672 5664 2848
tri 5664 2841 5677 2854 nw
rect 5750 2773 5765 3001
tri 5287 2651 5293 2657 se
rect 5293 2651 5302 2657
rect 5287 2635 5302 2651
tri 5302 2644 5315 2657 nw
rect 5456 2649 5473 2663
rect 5505 2649 5522 2663
tri 5649 2657 5664 2672 ne
tri 5664 2657 5686 2679 sw
rect 5287 2599 5302 2607
rect 5368 2635 5428 2649
rect 5383 2625 5428 2635
rect 5383 2607 5411 2625
tri 5287 2584 5302 2599 ne
tri 5302 2584 5324 2606 sw
rect 5368 2597 5411 2607
rect 5426 2621 5428 2625
rect 5550 2635 5610 2649
tri 5664 2644 5677 2657 ne
rect 5677 2651 5686 2657
tri 5686 2651 5692 2657 sw
rect 5550 2625 5595 2635
rect 5426 2597 5500 2621
rect 5368 2593 5500 2597
tri 5500 2593 5528 2621 sw
rect 5550 2611 5552 2625
tri 5550 2609 5552 2611 ne
rect 5564 2607 5595 2625
rect 5564 2597 5610 2607
rect 5677 2636 5692 2651
tri 5302 2572 5314 2584 ne
rect 5314 2579 5324 2584
tri 5324 2579 5329 2584 sw
rect 5213 2233 5228 2461
rect 5314 2423 5329 2579
rect 5368 2537 5396 2593
tri 5488 2575 5506 2593 ne
rect 5506 2573 5528 2593
tri 5528 2573 5548 2593 sw
tri 5564 2579 5582 2597 ne
rect 5387 2503 5396 2537
rect 5430 2564 5472 2565
rect 5430 2530 5435 2564
rect 5465 2530 5472 2564
rect 5430 2521 5472 2530
rect 5506 2564 5548 2573
rect 5506 2530 5513 2564
rect 5543 2530 5548 2564
rect 5506 2525 5548 2530
rect 5582 2537 5610 2597
tri 5655 2584 5677 2606 se
rect 5677 2599 5692 2607
tri 5677 2584 5692 2599 nw
tri 5649 2578 5655 2584 se
rect 5655 2578 5664 2584
rect 5368 2493 5396 2503
tri 5396 2493 5420 2517 sw
rect 5368 2461 5410 2493
tri 5427 2485 5428 2486 sw
rect 5427 2461 5428 2485
tri 5430 2484 5467 2521 ne
rect 5467 2493 5472 2521
tri 5472 2493 5498 2519 sw
rect 5582 2503 5591 2537
rect 5582 2493 5610 2503
rect 5467 2484 5551 2493
tri 5467 2465 5486 2484 ne
rect 5486 2465 5551 2484
rect 5368 2439 5428 2461
rect 5550 2461 5551 2465
rect 5568 2461 5610 2493
rect 5550 2439 5610 2461
rect 5456 2423 5473 2437
rect 5505 2423 5522 2437
tri 5293 2387 5315 2409 se
rect 5315 2402 5330 2423
tri 5315 2387 5330 2402 nw
rect 5649 2402 5664 2578
tri 5664 2571 5677 2584 nw
rect 5750 2503 5765 2731
tri 5287 2381 5293 2387 se
rect 5293 2381 5302 2387
rect 5287 2365 5302 2381
tri 5302 2374 5315 2387 nw
rect 5456 2379 5473 2393
rect 5505 2379 5522 2393
tri 5649 2387 5664 2402 ne
tri 5664 2387 5686 2409 sw
rect 5287 2329 5302 2337
rect 5368 2365 5428 2379
rect 5383 2355 5428 2365
rect 5383 2337 5411 2355
tri 5287 2314 5302 2329 ne
tri 5302 2314 5324 2336 sw
rect 5368 2327 5411 2337
rect 5426 2351 5428 2355
rect 5550 2365 5610 2379
tri 5664 2374 5677 2387 ne
rect 5677 2381 5686 2387
tri 5686 2381 5692 2387 sw
rect 5550 2355 5595 2365
rect 5426 2327 5500 2351
rect 5368 2323 5500 2327
tri 5500 2323 5528 2351 sw
rect 5550 2341 5552 2355
tri 5550 2339 5552 2341 ne
rect 5564 2337 5595 2355
rect 5564 2327 5610 2337
rect 5677 2366 5692 2381
tri 5302 2302 5314 2314 ne
rect 5314 2309 5324 2314
tri 5324 2309 5329 2314 sw
rect 5213 1963 5228 2191
rect 5314 2201 5329 2309
rect 5368 2267 5396 2323
tri 5488 2305 5506 2323 ne
rect 5506 2303 5528 2323
tri 5528 2303 5548 2323 sw
tri 5564 2309 5582 2327 ne
rect 5387 2233 5396 2267
rect 5430 2294 5472 2295
rect 5430 2260 5435 2294
rect 5465 2260 5472 2294
rect 5430 2251 5472 2260
rect 5506 2294 5548 2303
rect 5506 2260 5513 2294
rect 5543 2260 5548 2294
rect 5506 2255 5548 2260
rect 5582 2267 5610 2327
tri 5655 2314 5677 2336 se
rect 5677 2329 5692 2337
tri 5677 2314 5692 2329 nw
tri 5649 2308 5655 2314 se
rect 5655 2308 5664 2314
rect 5368 2223 5396 2233
tri 5396 2223 5420 2247 sw
rect 5314 2153 5330 2201
rect 5368 2191 5410 2223
tri 5427 2215 5428 2216 sw
rect 5427 2191 5428 2215
tri 5430 2214 5467 2251 ne
rect 5467 2223 5472 2251
tri 5472 2223 5498 2249 sw
rect 5582 2233 5591 2267
rect 5582 2223 5610 2233
rect 5467 2214 5551 2223
tri 5467 2195 5486 2214 ne
rect 5486 2195 5551 2214
rect 5368 2169 5428 2191
rect 5550 2191 5551 2195
rect 5568 2191 5610 2223
rect 5550 2169 5610 2191
rect 5456 2153 5473 2167
rect 5505 2153 5522 2167
tri 5293 2117 5315 2139 se
rect 5315 2132 5330 2153
tri 5315 2117 5330 2132 nw
rect 5649 2132 5664 2308
tri 5664 2301 5677 2314 nw
rect 5750 2233 5765 2461
tri 5287 2111 5293 2117 se
rect 5293 2111 5302 2117
rect 5287 2095 5302 2111
tri 5302 2104 5315 2117 nw
rect 5456 2109 5473 2123
rect 5505 2109 5522 2123
tri 5649 2117 5664 2132 ne
tri 5664 2117 5686 2139 sw
rect 5287 2059 5302 2067
rect 5368 2095 5428 2109
rect 5383 2085 5428 2095
rect 5383 2067 5411 2085
tri 5287 2044 5302 2059 ne
tri 5302 2044 5324 2066 sw
rect 5368 2057 5411 2067
rect 5426 2081 5428 2085
rect 5550 2095 5610 2109
tri 5664 2104 5677 2117 ne
rect 5677 2111 5686 2117
tri 5686 2111 5692 2117 sw
rect 5550 2085 5595 2095
rect 5426 2057 5500 2081
rect 5368 2053 5500 2057
tri 5500 2053 5528 2081 sw
rect 5550 2071 5552 2085
tri 5550 2069 5552 2071 ne
rect 5564 2067 5595 2085
rect 5564 2057 5610 2067
rect 5677 2096 5692 2111
tri 5302 2032 5314 2044 ne
rect 5314 2039 5324 2044
tri 5324 2039 5329 2044 sw
rect 5213 1693 5228 1921
rect 5314 1883 5329 2039
rect 5368 1997 5396 2053
tri 5488 2035 5506 2053 ne
rect 5506 2033 5528 2053
tri 5528 2033 5548 2053 sw
tri 5564 2039 5582 2057 ne
rect 5387 1963 5396 1997
rect 5430 2024 5472 2025
rect 5430 1990 5435 2024
rect 5465 1990 5472 2024
rect 5430 1981 5472 1990
rect 5506 2024 5548 2033
rect 5506 1990 5513 2024
rect 5543 1990 5548 2024
rect 5506 1985 5548 1990
rect 5582 1997 5610 2057
tri 5655 2044 5677 2066 se
rect 5677 2059 5692 2067
tri 5677 2044 5692 2059 nw
tri 5649 2038 5655 2044 se
rect 5655 2038 5664 2044
rect 5368 1953 5396 1963
tri 5396 1953 5420 1977 sw
rect 5368 1921 5410 1953
tri 5427 1945 5428 1946 sw
rect 5427 1921 5428 1945
tri 5430 1944 5467 1981 ne
rect 5467 1953 5472 1981
tri 5472 1953 5498 1979 sw
rect 5582 1963 5591 1997
rect 5582 1953 5610 1963
rect 5467 1944 5551 1953
tri 5467 1925 5486 1944 ne
rect 5486 1925 5551 1944
rect 5368 1899 5428 1921
rect 5550 1921 5551 1925
rect 5568 1921 5610 1953
rect 5550 1899 5610 1921
rect 5456 1883 5473 1897
rect 5505 1883 5522 1897
tri 5293 1847 5315 1869 se
rect 5315 1862 5330 1883
tri 5315 1847 5330 1862 nw
rect 5649 1862 5664 2038
tri 5664 2031 5677 2044 nw
rect 5750 1963 5765 2191
tri 5287 1841 5293 1847 se
rect 5293 1841 5302 1847
rect 5287 1825 5302 1841
tri 5302 1834 5315 1847 nw
rect 5456 1839 5473 1853
rect 5505 1839 5522 1853
tri 5649 1847 5664 1862 ne
tri 5664 1847 5686 1869 sw
rect 5287 1789 5302 1797
rect 5368 1825 5428 1839
rect 5383 1815 5428 1825
rect 5383 1797 5411 1815
tri 5287 1774 5302 1789 ne
tri 5302 1774 5324 1796 sw
rect 5368 1787 5411 1797
rect 5426 1811 5428 1815
rect 5550 1825 5610 1839
tri 5664 1834 5677 1847 ne
rect 5677 1841 5686 1847
tri 5686 1841 5692 1847 sw
rect 5550 1815 5595 1825
rect 5426 1787 5500 1811
rect 5368 1783 5500 1787
tri 5500 1783 5528 1811 sw
rect 5550 1801 5552 1815
tri 5550 1799 5552 1801 ne
rect 5564 1797 5595 1815
rect 5564 1787 5610 1797
rect 5677 1826 5692 1841
tri 5302 1762 5314 1774 ne
rect 5314 1769 5324 1774
tri 5324 1769 5329 1774 sw
rect 5213 1423 5228 1651
rect 5314 1661 5329 1769
rect 5368 1727 5396 1783
tri 5488 1765 5506 1783 ne
rect 5506 1763 5528 1783
tri 5528 1763 5548 1783 sw
tri 5564 1769 5582 1787 ne
rect 5387 1693 5396 1727
rect 5430 1754 5472 1755
rect 5430 1720 5435 1754
rect 5465 1720 5472 1754
rect 5430 1711 5472 1720
rect 5506 1754 5548 1763
rect 5506 1720 5513 1754
rect 5543 1720 5548 1754
rect 5506 1715 5548 1720
rect 5582 1727 5610 1787
tri 5655 1774 5677 1796 se
rect 5677 1789 5692 1797
tri 5677 1774 5692 1789 nw
tri 5649 1768 5655 1774 se
rect 5655 1768 5664 1774
rect 5368 1683 5396 1693
tri 5396 1683 5420 1707 sw
rect 5314 1613 5330 1661
rect 5368 1651 5410 1683
tri 5427 1675 5428 1676 sw
rect 5427 1651 5428 1675
tri 5430 1674 5467 1711 ne
rect 5467 1683 5472 1711
tri 5472 1683 5498 1709 sw
rect 5582 1693 5591 1727
rect 5582 1683 5610 1693
rect 5467 1674 5551 1683
tri 5467 1655 5486 1674 ne
rect 5486 1655 5551 1674
rect 5368 1629 5428 1651
rect 5550 1651 5551 1655
rect 5568 1651 5610 1683
rect 5550 1629 5610 1651
rect 5456 1613 5473 1627
rect 5505 1613 5522 1627
tri 5293 1577 5315 1599 se
rect 5315 1592 5330 1613
tri 5315 1577 5330 1592 nw
rect 5649 1592 5664 1768
tri 5664 1761 5677 1774 nw
rect 5750 1693 5765 1921
tri 5287 1571 5293 1577 se
rect 5293 1571 5302 1577
rect 5287 1555 5302 1571
tri 5302 1564 5315 1577 nw
rect 5456 1569 5473 1583
rect 5505 1569 5522 1583
tri 5649 1577 5664 1592 ne
tri 5664 1577 5686 1599 sw
rect 5287 1519 5302 1527
rect 5368 1555 5428 1569
rect 5383 1545 5428 1555
rect 5383 1527 5411 1545
tri 5287 1504 5302 1519 ne
tri 5302 1504 5324 1526 sw
rect 5368 1517 5411 1527
rect 5426 1541 5428 1545
rect 5550 1555 5610 1569
tri 5664 1564 5677 1577 ne
rect 5677 1571 5686 1577
tri 5686 1571 5692 1577 sw
rect 5550 1545 5595 1555
rect 5426 1517 5500 1541
rect 5368 1513 5500 1517
tri 5500 1513 5528 1541 sw
rect 5550 1531 5552 1545
tri 5550 1529 5552 1531 ne
rect 5564 1527 5595 1545
rect 5564 1517 5610 1527
rect 5677 1556 5692 1571
tri 5302 1492 5314 1504 ne
rect 5314 1499 5324 1504
tri 5324 1499 5329 1504 sw
rect 5213 1153 5228 1381
rect 5314 1343 5329 1499
rect 5368 1457 5396 1513
tri 5488 1495 5506 1513 ne
rect 5506 1493 5528 1513
tri 5528 1493 5548 1513 sw
tri 5564 1499 5582 1517 ne
rect 5387 1423 5396 1457
rect 5430 1484 5472 1485
rect 5430 1450 5435 1484
rect 5465 1450 5472 1484
rect 5430 1441 5472 1450
rect 5506 1484 5548 1493
rect 5506 1450 5513 1484
rect 5543 1450 5548 1484
rect 5506 1445 5548 1450
rect 5582 1457 5610 1517
tri 5655 1504 5677 1526 se
rect 5677 1519 5692 1527
tri 5677 1504 5692 1519 nw
tri 5649 1498 5655 1504 se
rect 5655 1498 5664 1504
rect 5368 1413 5396 1423
tri 5396 1413 5420 1437 sw
rect 5368 1381 5410 1413
tri 5427 1405 5428 1406 sw
rect 5427 1381 5428 1405
tri 5430 1404 5467 1441 ne
rect 5467 1413 5472 1441
tri 5472 1413 5498 1439 sw
rect 5582 1423 5591 1457
rect 5582 1413 5610 1423
rect 5467 1404 5551 1413
tri 5467 1385 5486 1404 ne
rect 5486 1385 5551 1404
rect 5368 1359 5428 1381
rect 5550 1381 5551 1385
rect 5568 1381 5610 1413
rect 5550 1359 5610 1381
rect 5456 1343 5473 1357
rect 5505 1343 5522 1357
tri 5293 1307 5315 1329 se
rect 5315 1322 5330 1343
tri 5315 1307 5330 1322 nw
rect 5649 1322 5664 1498
tri 5664 1491 5677 1504 nw
rect 5750 1423 5765 1651
tri 5287 1301 5293 1307 se
rect 5293 1301 5302 1307
rect 5287 1285 5302 1301
tri 5302 1294 5315 1307 nw
rect 5456 1299 5473 1313
rect 5505 1299 5522 1313
tri 5649 1307 5664 1322 ne
tri 5664 1307 5686 1329 sw
rect 5287 1249 5302 1257
rect 5368 1285 5428 1299
rect 5383 1275 5428 1285
rect 5383 1257 5411 1275
tri 5287 1234 5302 1249 ne
tri 5302 1234 5324 1256 sw
rect 5368 1247 5411 1257
rect 5426 1271 5428 1275
rect 5550 1285 5610 1299
tri 5664 1294 5677 1307 ne
rect 5677 1301 5686 1307
tri 5686 1301 5692 1307 sw
rect 5550 1275 5595 1285
rect 5426 1247 5500 1271
rect 5368 1243 5500 1247
tri 5500 1243 5528 1271 sw
rect 5550 1261 5552 1275
tri 5550 1259 5552 1261 ne
rect 5564 1257 5595 1275
rect 5564 1247 5610 1257
rect 5677 1286 5692 1301
tri 5302 1222 5314 1234 ne
rect 5314 1229 5324 1234
tri 5324 1229 5329 1234 sw
rect 5213 883 5228 1111
rect 5314 1121 5329 1229
rect 5368 1187 5396 1243
tri 5488 1225 5506 1243 ne
rect 5506 1223 5528 1243
tri 5528 1223 5548 1243 sw
tri 5564 1229 5582 1247 ne
rect 5387 1153 5396 1187
rect 5430 1214 5472 1215
rect 5430 1180 5435 1214
rect 5465 1180 5472 1214
rect 5430 1171 5472 1180
rect 5506 1214 5548 1223
rect 5506 1180 5513 1214
rect 5543 1180 5548 1214
rect 5506 1175 5548 1180
rect 5582 1187 5610 1247
tri 5655 1234 5677 1256 se
rect 5677 1249 5692 1257
tri 5677 1234 5692 1249 nw
tri 5649 1228 5655 1234 se
rect 5655 1228 5664 1234
rect 5368 1143 5396 1153
tri 5396 1143 5420 1167 sw
rect 5314 1073 5330 1121
rect 5368 1111 5410 1143
tri 5427 1135 5428 1136 sw
rect 5427 1111 5428 1135
tri 5430 1134 5467 1171 ne
rect 5467 1143 5472 1171
tri 5472 1143 5498 1169 sw
rect 5582 1153 5591 1187
rect 5582 1143 5610 1153
rect 5467 1134 5551 1143
tri 5467 1115 5486 1134 ne
rect 5486 1115 5551 1134
rect 5368 1089 5428 1111
rect 5550 1111 5551 1115
rect 5568 1111 5610 1143
rect 5550 1089 5610 1111
rect 5456 1073 5473 1087
rect 5505 1073 5522 1087
tri 5293 1037 5315 1059 se
rect 5315 1052 5330 1073
tri 5315 1037 5330 1052 nw
rect 5649 1052 5664 1228
tri 5664 1221 5677 1234 nw
rect 5750 1153 5765 1381
tri 5287 1031 5293 1037 se
rect 5293 1031 5302 1037
rect 5287 1015 5302 1031
tri 5302 1024 5315 1037 nw
rect 5456 1029 5473 1043
rect 5505 1029 5522 1043
tri 5649 1037 5664 1052 ne
tri 5664 1037 5686 1059 sw
rect 5287 979 5302 987
rect 5368 1015 5428 1029
rect 5383 1005 5428 1015
rect 5383 987 5411 1005
tri 5287 964 5302 979 ne
tri 5302 964 5324 986 sw
rect 5368 977 5411 987
rect 5426 1001 5428 1005
rect 5550 1015 5610 1029
tri 5664 1024 5677 1037 ne
rect 5677 1031 5686 1037
tri 5686 1031 5692 1037 sw
rect 5550 1005 5595 1015
rect 5426 977 5500 1001
rect 5368 973 5500 977
tri 5500 973 5528 1001 sw
rect 5550 991 5552 1005
tri 5550 989 5552 991 ne
rect 5564 987 5595 1005
rect 5564 977 5610 987
rect 5677 1016 5692 1031
tri 5302 952 5314 964 ne
rect 5314 959 5324 964
tri 5324 959 5329 964 sw
rect 5213 613 5228 841
rect 5314 803 5329 959
rect 5368 917 5396 973
tri 5488 955 5506 973 ne
rect 5506 953 5528 973
tri 5528 953 5548 973 sw
tri 5564 959 5582 977 ne
rect 5387 883 5396 917
rect 5430 944 5472 945
rect 5430 910 5435 944
rect 5465 910 5472 944
rect 5430 901 5472 910
rect 5506 944 5548 953
rect 5506 910 5513 944
rect 5543 910 5548 944
rect 5506 905 5548 910
rect 5582 917 5610 977
tri 5655 964 5677 986 se
rect 5677 979 5692 987
tri 5677 964 5692 979 nw
tri 5649 958 5655 964 se
rect 5655 958 5664 964
rect 5368 873 5396 883
tri 5396 873 5420 897 sw
rect 5368 841 5410 873
tri 5427 865 5428 866 sw
rect 5427 841 5428 865
tri 5430 864 5467 901 ne
rect 5467 873 5472 901
tri 5472 873 5498 899 sw
rect 5582 883 5591 917
rect 5582 873 5610 883
rect 5467 864 5551 873
tri 5467 845 5486 864 ne
rect 5486 845 5551 864
rect 5368 819 5428 841
rect 5550 841 5551 845
rect 5568 841 5610 873
rect 5550 819 5610 841
rect 5456 803 5473 817
rect 5505 803 5522 817
tri 5293 767 5315 789 se
rect 5315 782 5330 803
tri 5315 767 5330 782 nw
rect 5649 782 5664 958
tri 5664 951 5677 964 nw
rect 5750 883 5765 1111
tri 5287 761 5293 767 se
rect 5293 761 5302 767
rect 5287 745 5302 761
tri 5302 754 5315 767 nw
rect 5456 759 5473 773
rect 5505 759 5522 773
tri 5649 767 5664 782 ne
tri 5664 767 5686 789 sw
rect 5287 709 5302 717
rect 5368 745 5428 759
rect 5383 735 5428 745
rect 5383 717 5411 735
tri 5287 694 5302 709 ne
tri 5302 694 5324 716 sw
rect 5368 707 5411 717
rect 5426 731 5428 735
rect 5550 745 5610 759
tri 5664 754 5677 767 ne
rect 5677 761 5686 767
tri 5686 761 5692 767 sw
rect 5550 735 5595 745
rect 5426 707 5500 731
rect 5368 703 5500 707
tri 5500 703 5528 731 sw
rect 5550 721 5552 735
tri 5550 719 5552 721 ne
rect 5564 717 5595 735
rect 5564 707 5610 717
rect 5677 746 5692 761
tri 5302 682 5314 694 ne
rect 5314 689 5324 694
tri 5324 689 5329 694 sw
rect 5213 343 5228 571
rect 5314 581 5329 689
rect 5368 647 5396 703
tri 5488 685 5506 703 ne
rect 5506 683 5528 703
tri 5528 683 5548 703 sw
tri 5564 689 5582 707 ne
rect 5387 613 5396 647
rect 5430 674 5472 675
rect 5430 640 5435 674
rect 5465 640 5472 674
rect 5430 631 5472 640
rect 5506 674 5548 683
rect 5506 640 5513 674
rect 5543 640 5548 674
rect 5506 635 5548 640
rect 5582 647 5610 707
tri 5655 694 5677 716 se
rect 5677 709 5692 717
tri 5677 694 5692 709 nw
tri 5649 688 5655 694 se
rect 5655 688 5664 694
rect 5368 603 5396 613
tri 5396 603 5420 627 sw
rect 5314 533 5330 581
rect 5368 571 5410 603
tri 5427 595 5428 596 sw
rect 5427 571 5428 595
tri 5430 594 5467 631 ne
rect 5467 603 5472 631
tri 5472 603 5498 629 sw
rect 5582 613 5591 647
rect 5582 603 5610 613
rect 5467 594 5551 603
tri 5467 575 5486 594 ne
rect 5486 575 5551 594
rect 5368 549 5428 571
rect 5550 571 5551 575
rect 5568 571 5610 603
rect 5550 549 5610 571
rect 5456 533 5473 547
rect 5505 533 5522 547
tri 5293 497 5315 519 se
rect 5315 512 5330 533
tri 5315 497 5330 512 nw
rect 5649 512 5664 688
tri 5664 681 5677 694 nw
rect 5750 613 5765 841
tri 5287 491 5293 497 se
rect 5293 491 5302 497
rect 5287 475 5302 491
tri 5302 484 5315 497 nw
rect 5456 489 5473 503
rect 5505 489 5522 503
tri 5649 497 5664 512 ne
tri 5664 497 5686 519 sw
rect 5287 439 5302 447
rect 5368 475 5428 489
rect 5383 465 5428 475
rect 5383 447 5411 465
tri 5287 424 5302 439 ne
tri 5302 424 5324 446 sw
rect 5368 437 5411 447
rect 5426 461 5428 465
rect 5550 475 5610 489
tri 5664 484 5677 497 ne
rect 5677 491 5686 497
tri 5686 491 5692 497 sw
rect 5550 465 5595 475
rect 5426 437 5500 461
rect 5368 433 5500 437
tri 5500 433 5528 461 sw
rect 5550 451 5552 465
tri 5550 449 5552 451 ne
rect 5564 447 5595 465
rect 5564 437 5610 447
rect 5677 476 5692 491
tri 5302 412 5314 424 ne
rect 5314 419 5324 424
tri 5324 419 5329 424 sw
rect 5213 73 5228 301
rect 5314 263 5329 419
rect 5368 377 5396 433
tri 5488 415 5506 433 ne
rect 5506 413 5528 433
tri 5528 413 5548 433 sw
tri 5564 419 5582 437 ne
rect 5387 343 5396 377
rect 5430 404 5472 405
rect 5430 370 5435 404
rect 5465 370 5472 404
rect 5430 361 5472 370
rect 5506 404 5548 413
rect 5506 370 5513 404
rect 5543 370 5548 404
rect 5506 365 5548 370
rect 5582 377 5610 437
tri 5655 424 5677 446 se
rect 5677 439 5692 447
tri 5677 424 5692 439 nw
tri 5649 418 5655 424 se
rect 5655 418 5664 424
rect 5368 333 5396 343
tri 5396 333 5420 357 sw
rect 5368 301 5410 333
tri 5427 325 5428 326 sw
rect 5427 301 5428 325
tri 5430 324 5467 361 ne
rect 5467 333 5472 361
tri 5472 333 5498 359 sw
rect 5582 343 5591 377
rect 5582 333 5610 343
rect 5467 324 5551 333
tri 5467 305 5486 324 ne
rect 5486 305 5551 324
rect 5368 279 5428 301
rect 5550 301 5551 305
rect 5568 301 5610 333
rect 5550 279 5610 301
rect 5456 263 5473 277
rect 5505 263 5522 277
tri 5293 227 5315 249 se
rect 5315 242 5330 263
tri 5315 227 5330 242 nw
rect 5649 242 5664 418
tri 5664 411 5677 424 nw
rect 5750 343 5765 571
tri 5287 221 5293 227 se
rect 5293 221 5302 227
rect 5287 205 5302 221
tri 5302 214 5315 227 nw
rect 5456 219 5473 233
rect 5505 219 5522 233
tri 5649 227 5664 242 ne
tri 5664 227 5686 249 sw
rect 5287 169 5302 177
rect 5368 205 5428 219
rect 5383 195 5428 205
rect 5383 177 5411 195
tri 5287 154 5302 169 ne
tri 5302 154 5324 176 sw
rect 5368 167 5411 177
rect 5426 191 5428 195
rect 5550 205 5610 219
tri 5664 214 5677 227 ne
rect 5677 221 5686 227
tri 5686 221 5692 227 sw
rect 5550 195 5595 205
rect 5426 167 5500 191
rect 5368 163 5500 167
tri 5500 163 5528 191 sw
rect 5550 181 5552 195
tri 5550 179 5552 181 ne
rect 5564 177 5595 195
rect 5564 167 5610 177
rect 5677 206 5692 221
tri 5302 142 5314 154 ne
rect 5314 149 5324 154
tri 5324 149 5329 154 sw
rect 5213 -55 5228 31
rect 5314 -55 5329 149
rect 5368 107 5396 163
tri 5488 145 5506 163 ne
rect 5506 143 5528 163
tri 5528 143 5548 163 sw
tri 5564 149 5582 167 ne
rect 5387 73 5396 107
rect 5430 134 5472 135
rect 5430 100 5435 134
rect 5465 100 5472 134
rect 5430 91 5472 100
rect 5506 134 5548 143
rect 5506 100 5513 134
rect 5543 100 5548 134
rect 5506 95 5548 100
rect 5582 107 5610 167
tri 5655 154 5677 176 se
rect 5677 169 5692 177
tri 5677 154 5692 169 nw
tri 5649 148 5655 154 se
rect 5655 148 5664 154
rect 5368 63 5396 73
tri 5396 63 5420 87 sw
rect 5368 31 5410 63
tri 5427 55 5428 56 sw
rect 5427 31 5428 55
tri 5430 54 5467 91 ne
rect 5467 63 5472 91
tri 5472 63 5498 89 sw
rect 5582 73 5591 107
rect 5582 63 5610 73
rect 5467 54 5551 63
tri 5467 35 5486 54 ne
rect 5486 35 5551 54
rect 5368 9 5428 31
rect 5550 31 5551 35
rect 5568 31 5610 63
rect 5550 9 5610 31
rect 5456 -7 5473 7
rect 5505 -7 5522 7
rect 5649 -55 5664 148
tri 5664 141 5677 154 nw
rect 5750 73 5765 301
rect 5750 -55 5765 31
rect 5793 4123 5808 4361
tri 5873 4277 5895 4299 se
rect 5895 4292 5910 4361
tri 5895 4277 5910 4292 nw
rect 6229 4292 6244 4361
tri 5867 4271 5873 4277 se
rect 5873 4271 5882 4277
rect 5867 4255 5882 4271
tri 5882 4264 5895 4277 nw
rect 6036 4269 6053 4283
rect 6085 4269 6102 4283
tri 6229 4277 6244 4292 ne
tri 6244 4277 6266 4299 sw
rect 5867 4219 5882 4227
rect 5948 4255 6008 4269
rect 5963 4245 6008 4255
rect 5963 4227 5991 4245
tri 5867 4204 5882 4219 ne
tri 5882 4204 5904 4226 sw
rect 5948 4217 5991 4227
rect 6006 4241 6008 4245
rect 6130 4255 6190 4269
tri 6244 4264 6257 4277 ne
rect 6257 4271 6266 4277
tri 6266 4271 6272 4277 sw
rect 6130 4245 6175 4255
rect 6006 4217 6080 4241
rect 5948 4213 6080 4217
tri 6080 4213 6108 4241 sw
rect 6130 4231 6132 4245
tri 6130 4229 6132 4231 ne
rect 6144 4227 6175 4245
rect 6144 4217 6190 4227
rect 6257 4256 6272 4271
tri 5882 4192 5894 4204 ne
rect 5894 4199 5904 4204
tri 5904 4199 5909 4204 sw
rect 5793 3853 5808 4081
rect 5894 4043 5909 4199
rect 5948 4157 5976 4213
tri 6068 4195 6086 4213 ne
rect 6086 4193 6108 4213
tri 6108 4193 6128 4213 sw
tri 6144 4199 6162 4217 ne
rect 5967 4123 5976 4157
rect 6010 4184 6052 4185
rect 6010 4150 6015 4184
rect 6045 4150 6052 4184
rect 6010 4141 6052 4150
rect 6086 4184 6128 4193
rect 6086 4150 6093 4184
rect 6123 4150 6128 4184
rect 6086 4145 6128 4150
rect 6162 4157 6190 4217
tri 6235 4204 6257 4226 se
rect 6257 4219 6272 4227
tri 6257 4204 6272 4219 nw
tri 6229 4198 6235 4204 se
rect 6235 4198 6244 4204
rect 5948 4113 5976 4123
tri 5976 4113 6000 4137 sw
rect 5948 4081 5990 4113
tri 6007 4105 6008 4106 sw
rect 6007 4081 6008 4105
tri 6010 4104 6047 4141 ne
rect 6047 4113 6052 4141
tri 6052 4113 6078 4139 sw
rect 6162 4123 6171 4157
rect 6162 4113 6190 4123
rect 6047 4104 6131 4113
tri 6047 4085 6066 4104 ne
rect 6066 4085 6131 4104
rect 5948 4059 6008 4081
rect 6130 4081 6131 4085
rect 6148 4081 6190 4113
rect 6130 4059 6190 4081
rect 6036 4043 6053 4057
rect 6085 4043 6102 4057
tri 5873 4007 5895 4029 se
rect 5895 4022 5910 4043
tri 5895 4007 5910 4022 nw
rect 6229 4022 6244 4198
tri 6244 4191 6257 4204 nw
rect 6330 4123 6345 4361
tri 5867 4001 5873 4007 se
rect 5873 4001 5882 4007
rect 5867 3985 5882 4001
tri 5882 3994 5895 4007 nw
rect 6036 3999 6053 4013
rect 6085 3999 6102 4013
tri 6229 4007 6244 4022 ne
tri 6244 4007 6266 4029 sw
rect 5867 3949 5882 3957
rect 5948 3985 6008 3999
rect 5963 3975 6008 3985
rect 5963 3957 5991 3975
tri 5867 3934 5882 3949 ne
tri 5882 3934 5904 3956 sw
rect 5948 3947 5991 3957
rect 6006 3971 6008 3975
rect 6130 3985 6190 3999
tri 6244 3994 6257 4007 ne
rect 6257 4001 6266 4007
tri 6266 4001 6272 4007 sw
rect 6130 3975 6175 3985
rect 6006 3947 6080 3971
rect 5948 3943 6080 3947
tri 6080 3943 6108 3971 sw
rect 6130 3961 6132 3975
tri 6130 3959 6132 3961 ne
rect 6144 3957 6175 3975
rect 6144 3947 6190 3957
rect 6257 3986 6272 4001
tri 5882 3922 5894 3934 ne
rect 5894 3929 5904 3934
tri 5904 3929 5909 3934 sw
rect 5793 3583 5808 3811
rect 5894 3821 5909 3929
rect 5948 3887 5976 3943
tri 6068 3925 6086 3943 ne
rect 6086 3923 6108 3943
tri 6108 3923 6128 3943 sw
tri 6144 3929 6162 3947 ne
rect 5967 3853 5976 3887
rect 6010 3914 6052 3915
rect 6010 3880 6015 3914
rect 6045 3880 6052 3914
rect 6010 3871 6052 3880
rect 6086 3914 6128 3923
rect 6086 3880 6093 3914
rect 6123 3880 6128 3914
rect 6086 3875 6128 3880
rect 6162 3887 6190 3947
tri 6235 3934 6257 3956 se
rect 6257 3949 6272 3957
tri 6257 3934 6272 3949 nw
tri 6229 3928 6235 3934 se
rect 6235 3928 6244 3934
rect 5948 3843 5976 3853
tri 5976 3843 6000 3867 sw
rect 5894 3773 5910 3821
rect 5948 3811 5990 3843
tri 6007 3835 6008 3836 sw
rect 6007 3811 6008 3835
tri 6010 3834 6047 3871 ne
rect 6047 3843 6052 3871
tri 6052 3843 6078 3869 sw
rect 6162 3853 6171 3887
rect 6162 3843 6190 3853
rect 6047 3834 6131 3843
tri 6047 3815 6066 3834 ne
rect 6066 3815 6131 3834
rect 5948 3789 6008 3811
rect 6130 3811 6131 3815
rect 6148 3811 6190 3843
rect 6130 3789 6190 3811
rect 6036 3773 6053 3787
rect 6085 3773 6102 3787
tri 5873 3737 5895 3759 se
rect 5895 3752 5910 3773
tri 5895 3737 5910 3752 nw
rect 6229 3752 6244 3928
tri 6244 3921 6257 3934 nw
rect 6330 3853 6345 4081
tri 5867 3731 5873 3737 se
rect 5873 3731 5882 3737
rect 5867 3715 5882 3731
tri 5882 3724 5895 3737 nw
rect 6036 3729 6053 3743
rect 6085 3729 6102 3743
tri 6229 3737 6244 3752 ne
tri 6244 3737 6266 3759 sw
rect 5867 3679 5882 3687
rect 5948 3715 6008 3729
rect 5963 3705 6008 3715
rect 5963 3687 5991 3705
tri 5867 3664 5882 3679 ne
tri 5882 3664 5904 3686 sw
rect 5948 3677 5991 3687
rect 6006 3701 6008 3705
rect 6130 3715 6190 3729
tri 6244 3724 6257 3737 ne
rect 6257 3731 6266 3737
tri 6266 3731 6272 3737 sw
rect 6130 3705 6175 3715
rect 6006 3677 6080 3701
rect 5948 3673 6080 3677
tri 6080 3673 6108 3701 sw
rect 6130 3691 6132 3705
tri 6130 3689 6132 3691 ne
rect 6144 3687 6175 3705
rect 6144 3677 6190 3687
rect 6257 3716 6272 3731
tri 5882 3652 5894 3664 ne
rect 5894 3659 5904 3664
tri 5904 3659 5909 3664 sw
rect 5793 3313 5808 3541
rect 5894 3503 5909 3659
rect 5948 3617 5976 3673
tri 6068 3655 6086 3673 ne
rect 6086 3653 6108 3673
tri 6108 3653 6128 3673 sw
tri 6144 3659 6162 3677 ne
rect 5967 3583 5976 3617
rect 6010 3644 6052 3645
rect 6010 3610 6015 3644
rect 6045 3610 6052 3644
rect 6010 3601 6052 3610
rect 6086 3644 6128 3653
rect 6086 3610 6093 3644
rect 6123 3610 6128 3644
rect 6086 3605 6128 3610
rect 6162 3617 6190 3677
tri 6235 3664 6257 3686 se
rect 6257 3679 6272 3687
tri 6257 3664 6272 3679 nw
tri 6229 3658 6235 3664 se
rect 6235 3658 6244 3664
rect 5948 3573 5976 3583
tri 5976 3573 6000 3597 sw
rect 5948 3541 5990 3573
tri 6007 3565 6008 3566 sw
rect 6007 3541 6008 3565
tri 6010 3564 6047 3601 ne
rect 6047 3573 6052 3601
tri 6052 3573 6078 3599 sw
rect 6162 3583 6171 3617
rect 6162 3573 6190 3583
rect 6047 3564 6131 3573
tri 6047 3545 6066 3564 ne
rect 6066 3545 6131 3564
rect 5948 3519 6008 3541
rect 6130 3541 6131 3545
rect 6148 3541 6190 3573
rect 6130 3519 6190 3541
rect 6036 3503 6053 3517
rect 6085 3503 6102 3517
tri 5873 3467 5895 3489 se
rect 5895 3482 5910 3503
tri 5895 3467 5910 3482 nw
rect 6229 3482 6244 3658
tri 6244 3651 6257 3664 nw
rect 6330 3583 6345 3811
tri 5867 3461 5873 3467 se
rect 5873 3461 5882 3467
rect 5867 3445 5882 3461
tri 5882 3454 5895 3467 nw
rect 6036 3459 6053 3473
rect 6085 3459 6102 3473
tri 6229 3467 6244 3482 ne
tri 6244 3467 6266 3489 sw
rect 5867 3409 5882 3417
rect 5948 3445 6008 3459
rect 5963 3435 6008 3445
rect 5963 3417 5991 3435
tri 5867 3394 5882 3409 ne
tri 5882 3394 5904 3416 sw
rect 5948 3407 5991 3417
rect 6006 3431 6008 3435
rect 6130 3445 6190 3459
tri 6244 3454 6257 3467 ne
rect 6257 3461 6266 3467
tri 6266 3461 6272 3467 sw
rect 6130 3435 6175 3445
rect 6006 3407 6080 3431
rect 5948 3403 6080 3407
tri 6080 3403 6108 3431 sw
rect 6130 3421 6132 3435
tri 6130 3419 6132 3421 ne
rect 6144 3417 6175 3435
rect 6144 3407 6190 3417
rect 6257 3446 6272 3461
tri 5882 3382 5894 3394 ne
rect 5894 3389 5904 3394
tri 5904 3389 5909 3394 sw
rect 5793 3043 5808 3271
rect 5894 3281 5909 3389
rect 5948 3347 5976 3403
tri 6068 3385 6086 3403 ne
rect 6086 3383 6108 3403
tri 6108 3383 6128 3403 sw
tri 6144 3389 6162 3407 ne
rect 5967 3313 5976 3347
rect 6010 3374 6052 3375
rect 6010 3340 6015 3374
rect 6045 3340 6052 3374
rect 6010 3331 6052 3340
rect 6086 3374 6128 3383
rect 6086 3340 6093 3374
rect 6123 3340 6128 3374
rect 6086 3335 6128 3340
rect 6162 3347 6190 3407
tri 6235 3394 6257 3416 se
rect 6257 3409 6272 3417
tri 6257 3394 6272 3409 nw
tri 6229 3388 6235 3394 se
rect 6235 3388 6244 3394
rect 5948 3303 5976 3313
tri 5976 3303 6000 3327 sw
rect 5894 3233 5910 3281
rect 5948 3271 5990 3303
tri 6007 3295 6008 3296 sw
rect 6007 3271 6008 3295
tri 6010 3294 6047 3331 ne
rect 6047 3303 6052 3331
tri 6052 3303 6078 3329 sw
rect 6162 3313 6171 3347
rect 6162 3303 6190 3313
rect 6047 3294 6131 3303
tri 6047 3275 6066 3294 ne
rect 6066 3275 6131 3294
rect 5948 3249 6008 3271
rect 6130 3271 6131 3275
rect 6148 3271 6190 3303
rect 6130 3249 6190 3271
rect 6036 3233 6053 3247
rect 6085 3233 6102 3247
tri 5873 3197 5895 3219 se
rect 5895 3212 5910 3233
tri 5895 3197 5910 3212 nw
rect 6229 3212 6244 3388
tri 6244 3381 6257 3394 nw
rect 6330 3313 6345 3541
tri 5867 3191 5873 3197 se
rect 5873 3191 5882 3197
rect 5867 3175 5882 3191
tri 5882 3184 5895 3197 nw
rect 6036 3189 6053 3203
rect 6085 3189 6102 3203
tri 6229 3197 6244 3212 ne
tri 6244 3197 6266 3219 sw
rect 5867 3139 5882 3147
rect 5948 3175 6008 3189
rect 5963 3165 6008 3175
rect 5963 3147 5991 3165
tri 5867 3124 5882 3139 ne
tri 5882 3124 5904 3146 sw
rect 5948 3137 5991 3147
rect 6006 3161 6008 3165
rect 6130 3175 6190 3189
tri 6244 3184 6257 3197 ne
rect 6257 3191 6266 3197
tri 6266 3191 6272 3197 sw
rect 6130 3165 6175 3175
rect 6006 3137 6080 3161
rect 5948 3133 6080 3137
tri 6080 3133 6108 3161 sw
rect 6130 3151 6132 3165
tri 6130 3149 6132 3151 ne
rect 6144 3147 6175 3165
rect 6144 3137 6190 3147
rect 6257 3176 6272 3191
tri 5882 3112 5894 3124 ne
rect 5894 3119 5904 3124
tri 5904 3119 5909 3124 sw
rect 5793 2773 5808 3001
rect 5894 2963 5909 3119
rect 5948 3077 5976 3133
tri 6068 3115 6086 3133 ne
rect 6086 3113 6108 3133
tri 6108 3113 6128 3133 sw
tri 6144 3119 6162 3137 ne
rect 5967 3043 5976 3077
rect 6010 3104 6052 3105
rect 6010 3070 6015 3104
rect 6045 3070 6052 3104
rect 6010 3061 6052 3070
rect 6086 3104 6128 3113
rect 6086 3070 6093 3104
rect 6123 3070 6128 3104
rect 6086 3065 6128 3070
rect 6162 3077 6190 3137
tri 6235 3124 6257 3146 se
rect 6257 3139 6272 3147
tri 6257 3124 6272 3139 nw
tri 6229 3118 6235 3124 se
rect 6235 3118 6244 3124
rect 5948 3033 5976 3043
tri 5976 3033 6000 3057 sw
rect 5948 3001 5990 3033
tri 6007 3025 6008 3026 sw
rect 6007 3001 6008 3025
tri 6010 3024 6047 3061 ne
rect 6047 3033 6052 3061
tri 6052 3033 6078 3059 sw
rect 6162 3043 6171 3077
rect 6162 3033 6190 3043
rect 6047 3024 6131 3033
tri 6047 3005 6066 3024 ne
rect 6066 3005 6131 3024
rect 5948 2979 6008 3001
rect 6130 3001 6131 3005
rect 6148 3001 6190 3033
rect 6130 2979 6190 3001
rect 6036 2963 6053 2977
rect 6085 2963 6102 2977
tri 5873 2927 5895 2949 se
rect 5895 2942 5910 2963
tri 5895 2927 5910 2942 nw
rect 6229 2942 6244 3118
tri 6244 3111 6257 3124 nw
rect 6330 3043 6345 3271
tri 5867 2921 5873 2927 se
rect 5873 2921 5882 2927
rect 5867 2905 5882 2921
tri 5882 2914 5895 2927 nw
rect 6036 2919 6053 2933
rect 6085 2919 6102 2933
tri 6229 2927 6244 2942 ne
tri 6244 2927 6266 2949 sw
rect 5867 2869 5882 2877
rect 5948 2905 6008 2919
rect 5963 2895 6008 2905
rect 5963 2877 5991 2895
tri 5867 2854 5882 2869 ne
tri 5882 2854 5904 2876 sw
rect 5948 2867 5991 2877
rect 6006 2891 6008 2895
rect 6130 2905 6190 2919
tri 6244 2914 6257 2927 ne
rect 6257 2921 6266 2927
tri 6266 2921 6272 2927 sw
rect 6130 2895 6175 2905
rect 6006 2867 6080 2891
rect 5948 2863 6080 2867
tri 6080 2863 6108 2891 sw
rect 6130 2881 6132 2895
tri 6130 2879 6132 2881 ne
rect 6144 2877 6175 2895
rect 6144 2867 6190 2877
rect 6257 2906 6272 2921
tri 5882 2842 5894 2854 ne
rect 5894 2849 5904 2854
tri 5904 2849 5909 2854 sw
rect 5793 2503 5808 2731
rect 5894 2741 5909 2849
rect 5948 2807 5976 2863
tri 6068 2845 6086 2863 ne
rect 6086 2843 6108 2863
tri 6108 2843 6128 2863 sw
tri 6144 2849 6162 2867 ne
rect 5967 2773 5976 2807
rect 6010 2834 6052 2835
rect 6010 2800 6015 2834
rect 6045 2800 6052 2834
rect 6010 2791 6052 2800
rect 6086 2834 6128 2843
rect 6086 2800 6093 2834
rect 6123 2800 6128 2834
rect 6086 2795 6128 2800
rect 6162 2807 6190 2867
tri 6235 2854 6257 2876 se
rect 6257 2869 6272 2877
tri 6257 2854 6272 2869 nw
tri 6229 2848 6235 2854 se
rect 6235 2848 6244 2854
rect 5948 2763 5976 2773
tri 5976 2763 6000 2787 sw
rect 5894 2693 5910 2741
rect 5948 2731 5990 2763
tri 6007 2755 6008 2756 sw
rect 6007 2731 6008 2755
tri 6010 2754 6047 2791 ne
rect 6047 2763 6052 2791
tri 6052 2763 6078 2789 sw
rect 6162 2773 6171 2807
rect 6162 2763 6190 2773
rect 6047 2754 6131 2763
tri 6047 2735 6066 2754 ne
rect 6066 2735 6131 2754
rect 5948 2709 6008 2731
rect 6130 2731 6131 2735
rect 6148 2731 6190 2763
rect 6130 2709 6190 2731
rect 6036 2693 6053 2707
rect 6085 2693 6102 2707
tri 5873 2657 5895 2679 se
rect 5895 2672 5910 2693
tri 5895 2657 5910 2672 nw
rect 6229 2672 6244 2848
tri 6244 2841 6257 2854 nw
rect 6330 2773 6345 3001
tri 5867 2651 5873 2657 se
rect 5873 2651 5882 2657
rect 5867 2635 5882 2651
tri 5882 2644 5895 2657 nw
rect 6036 2649 6053 2663
rect 6085 2649 6102 2663
tri 6229 2657 6244 2672 ne
tri 6244 2657 6266 2679 sw
rect 5867 2599 5882 2607
rect 5948 2635 6008 2649
rect 5963 2625 6008 2635
rect 5963 2607 5991 2625
tri 5867 2584 5882 2599 ne
tri 5882 2584 5904 2606 sw
rect 5948 2597 5991 2607
rect 6006 2621 6008 2625
rect 6130 2635 6190 2649
tri 6244 2644 6257 2657 ne
rect 6257 2651 6266 2657
tri 6266 2651 6272 2657 sw
rect 6130 2625 6175 2635
rect 6006 2597 6080 2621
rect 5948 2593 6080 2597
tri 6080 2593 6108 2621 sw
rect 6130 2611 6132 2625
tri 6130 2609 6132 2611 ne
rect 6144 2607 6175 2625
rect 6144 2597 6190 2607
rect 6257 2636 6272 2651
tri 5882 2572 5894 2584 ne
rect 5894 2579 5904 2584
tri 5904 2579 5909 2584 sw
rect 5793 2233 5808 2461
rect 5894 2423 5909 2579
rect 5948 2537 5976 2593
tri 6068 2575 6086 2593 ne
rect 6086 2573 6108 2593
tri 6108 2573 6128 2593 sw
tri 6144 2579 6162 2597 ne
rect 5967 2503 5976 2537
rect 6010 2564 6052 2565
rect 6010 2530 6015 2564
rect 6045 2530 6052 2564
rect 6010 2521 6052 2530
rect 6086 2564 6128 2573
rect 6086 2530 6093 2564
rect 6123 2530 6128 2564
rect 6086 2525 6128 2530
rect 6162 2537 6190 2597
tri 6235 2584 6257 2606 se
rect 6257 2599 6272 2607
tri 6257 2584 6272 2599 nw
tri 6229 2578 6235 2584 se
rect 6235 2578 6244 2584
rect 5948 2493 5976 2503
tri 5976 2493 6000 2517 sw
rect 5948 2461 5990 2493
tri 6007 2485 6008 2486 sw
rect 6007 2461 6008 2485
tri 6010 2484 6047 2521 ne
rect 6047 2493 6052 2521
tri 6052 2493 6078 2519 sw
rect 6162 2503 6171 2537
rect 6162 2493 6190 2503
rect 6047 2484 6131 2493
tri 6047 2465 6066 2484 ne
rect 6066 2465 6131 2484
rect 5948 2439 6008 2461
rect 6130 2461 6131 2465
rect 6148 2461 6190 2493
rect 6130 2439 6190 2461
rect 6036 2423 6053 2437
rect 6085 2423 6102 2437
tri 5873 2387 5895 2409 se
rect 5895 2402 5910 2423
tri 5895 2387 5910 2402 nw
rect 6229 2402 6244 2578
tri 6244 2571 6257 2584 nw
rect 6330 2503 6345 2731
tri 5867 2381 5873 2387 se
rect 5873 2381 5882 2387
rect 5867 2365 5882 2381
tri 5882 2374 5895 2387 nw
rect 6036 2379 6053 2393
rect 6085 2379 6102 2393
tri 6229 2387 6244 2402 ne
tri 6244 2387 6266 2409 sw
rect 5867 2329 5882 2337
rect 5948 2365 6008 2379
rect 5963 2355 6008 2365
rect 5963 2337 5991 2355
tri 5867 2314 5882 2329 ne
tri 5882 2314 5904 2336 sw
rect 5948 2327 5991 2337
rect 6006 2351 6008 2355
rect 6130 2365 6190 2379
tri 6244 2374 6257 2387 ne
rect 6257 2381 6266 2387
tri 6266 2381 6272 2387 sw
rect 6130 2355 6175 2365
rect 6006 2327 6080 2351
rect 5948 2323 6080 2327
tri 6080 2323 6108 2351 sw
rect 6130 2341 6132 2355
tri 6130 2339 6132 2341 ne
rect 6144 2337 6175 2355
rect 6144 2327 6190 2337
rect 6257 2366 6272 2381
tri 5882 2302 5894 2314 ne
rect 5894 2309 5904 2314
tri 5904 2309 5909 2314 sw
rect 5793 1963 5808 2191
rect 5894 2201 5909 2309
rect 5948 2267 5976 2323
tri 6068 2305 6086 2323 ne
rect 6086 2303 6108 2323
tri 6108 2303 6128 2323 sw
tri 6144 2309 6162 2327 ne
rect 5967 2233 5976 2267
rect 6010 2294 6052 2295
rect 6010 2260 6015 2294
rect 6045 2260 6052 2294
rect 6010 2251 6052 2260
rect 6086 2294 6128 2303
rect 6086 2260 6093 2294
rect 6123 2260 6128 2294
rect 6086 2255 6128 2260
rect 6162 2267 6190 2327
tri 6235 2314 6257 2336 se
rect 6257 2329 6272 2337
tri 6257 2314 6272 2329 nw
tri 6229 2308 6235 2314 se
rect 6235 2308 6244 2314
rect 5948 2223 5976 2233
tri 5976 2223 6000 2247 sw
rect 5894 2153 5910 2201
rect 5948 2191 5990 2223
tri 6007 2215 6008 2216 sw
rect 6007 2191 6008 2215
tri 6010 2214 6047 2251 ne
rect 6047 2223 6052 2251
tri 6052 2223 6078 2249 sw
rect 6162 2233 6171 2267
rect 6162 2223 6190 2233
rect 6047 2214 6131 2223
tri 6047 2195 6066 2214 ne
rect 6066 2195 6131 2214
rect 5948 2169 6008 2191
rect 6130 2191 6131 2195
rect 6148 2191 6190 2223
rect 6130 2169 6190 2191
rect 6036 2153 6053 2167
rect 6085 2153 6102 2167
tri 5873 2117 5895 2139 se
rect 5895 2132 5910 2153
tri 5895 2117 5910 2132 nw
rect 6229 2132 6244 2308
tri 6244 2301 6257 2314 nw
rect 6330 2233 6345 2461
tri 5867 2111 5873 2117 se
rect 5873 2111 5882 2117
rect 5867 2095 5882 2111
tri 5882 2104 5895 2117 nw
rect 6036 2109 6053 2123
rect 6085 2109 6102 2123
tri 6229 2117 6244 2132 ne
tri 6244 2117 6266 2139 sw
rect 5867 2059 5882 2067
rect 5948 2095 6008 2109
rect 5963 2085 6008 2095
rect 5963 2067 5991 2085
tri 5867 2044 5882 2059 ne
tri 5882 2044 5904 2066 sw
rect 5948 2057 5991 2067
rect 6006 2081 6008 2085
rect 6130 2095 6190 2109
tri 6244 2104 6257 2117 ne
rect 6257 2111 6266 2117
tri 6266 2111 6272 2117 sw
rect 6130 2085 6175 2095
rect 6006 2057 6080 2081
rect 5948 2053 6080 2057
tri 6080 2053 6108 2081 sw
rect 6130 2071 6132 2085
tri 6130 2069 6132 2071 ne
rect 6144 2067 6175 2085
rect 6144 2057 6190 2067
rect 6257 2096 6272 2111
tri 5882 2032 5894 2044 ne
rect 5894 2039 5904 2044
tri 5904 2039 5909 2044 sw
rect 5793 1693 5808 1921
rect 5894 1883 5909 2039
rect 5948 1997 5976 2053
tri 6068 2035 6086 2053 ne
rect 6086 2033 6108 2053
tri 6108 2033 6128 2053 sw
tri 6144 2039 6162 2057 ne
rect 5967 1963 5976 1997
rect 6010 2024 6052 2025
rect 6010 1990 6015 2024
rect 6045 1990 6052 2024
rect 6010 1981 6052 1990
rect 6086 2024 6128 2033
rect 6086 1990 6093 2024
rect 6123 1990 6128 2024
rect 6086 1985 6128 1990
rect 6162 1997 6190 2057
tri 6235 2044 6257 2066 se
rect 6257 2059 6272 2067
tri 6257 2044 6272 2059 nw
tri 6229 2038 6235 2044 se
rect 6235 2038 6244 2044
rect 5948 1953 5976 1963
tri 5976 1953 6000 1977 sw
rect 5948 1921 5990 1953
tri 6007 1945 6008 1946 sw
rect 6007 1921 6008 1945
tri 6010 1944 6047 1981 ne
rect 6047 1953 6052 1981
tri 6052 1953 6078 1979 sw
rect 6162 1963 6171 1997
rect 6162 1953 6190 1963
rect 6047 1944 6131 1953
tri 6047 1925 6066 1944 ne
rect 6066 1925 6131 1944
rect 5948 1899 6008 1921
rect 6130 1921 6131 1925
rect 6148 1921 6190 1953
rect 6130 1899 6190 1921
rect 6036 1883 6053 1897
rect 6085 1883 6102 1897
tri 5873 1847 5895 1869 se
rect 5895 1862 5910 1883
tri 5895 1847 5910 1862 nw
rect 6229 1862 6244 2038
tri 6244 2031 6257 2044 nw
rect 6330 1963 6345 2191
tri 5867 1841 5873 1847 se
rect 5873 1841 5882 1847
rect 5867 1825 5882 1841
tri 5882 1834 5895 1847 nw
rect 6036 1839 6053 1853
rect 6085 1839 6102 1853
tri 6229 1847 6244 1862 ne
tri 6244 1847 6266 1869 sw
rect 5867 1789 5882 1797
rect 5948 1825 6008 1839
rect 5963 1815 6008 1825
rect 5963 1797 5991 1815
tri 5867 1774 5882 1789 ne
tri 5882 1774 5904 1796 sw
rect 5948 1787 5991 1797
rect 6006 1811 6008 1815
rect 6130 1825 6190 1839
tri 6244 1834 6257 1847 ne
rect 6257 1841 6266 1847
tri 6266 1841 6272 1847 sw
rect 6130 1815 6175 1825
rect 6006 1787 6080 1811
rect 5948 1783 6080 1787
tri 6080 1783 6108 1811 sw
rect 6130 1801 6132 1815
tri 6130 1799 6132 1801 ne
rect 6144 1797 6175 1815
rect 6144 1787 6190 1797
rect 6257 1826 6272 1841
tri 5882 1762 5894 1774 ne
rect 5894 1769 5904 1774
tri 5904 1769 5909 1774 sw
rect 5793 1423 5808 1651
rect 5894 1661 5909 1769
rect 5948 1727 5976 1783
tri 6068 1765 6086 1783 ne
rect 6086 1763 6108 1783
tri 6108 1763 6128 1783 sw
tri 6144 1769 6162 1787 ne
rect 5967 1693 5976 1727
rect 6010 1754 6052 1755
rect 6010 1720 6015 1754
rect 6045 1720 6052 1754
rect 6010 1711 6052 1720
rect 6086 1754 6128 1763
rect 6086 1720 6093 1754
rect 6123 1720 6128 1754
rect 6086 1715 6128 1720
rect 6162 1727 6190 1787
tri 6235 1774 6257 1796 se
rect 6257 1789 6272 1797
tri 6257 1774 6272 1789 nw
tri 6229 1768 6235 1774 se
rect 6235 1768 6244 1774
rect 5948 1683 5976 1693
tri 5976 1683 6000 1707 sw
rect 5894 1613 5910 1661
rect 5948 1651 5990 1683
tri 6007 1675 6008 1676 sw
rect 6007 1651 6008 1675
tri 6010 1674 6047 1711 ne
rect 6047 1683 6052 1711
tri 6052 1683 6078 1709 sw
rect 6162 1693 6171 1727
rect 6162 1683 6190 1693
rect 6047 1674 6131 1683
tri 6047 1655 6066 1674 ne
rect 6066 1655 6131 1674
rect 5948 1629 6008 1651
rect 6130 1651 6131 1655
rect 6148 1651 6190 1683
rect 6130 1629 6190 1651
rect 6036 1613 6053 1627
rect 6085 1613 6102 1627
tri 5873 1577 5895 1599 se
rect 5895 1592 5910 1613
tri 5895 1577 5910 1592 nw
rect 6229 1592 6244 1768
tri 6244 1761 6257 1774 nw
rect 6330 1693 6345 1921
tri 5867 1571 5873 1577 se
rect 5873 1571 5882 1577
rect 5867 1555 5882 1571
tri 5882 1564 5895 1577 nw
rect 6036 1569 6053 1583
rect 6085 1569 6102 1583
tri 6229 1577 6244 1592 ne
tri 6244 1577 6266 1599 sw
rect 5867 1519 5882 1527
rect 5948 1555 6008 1569
rect 5963 1545 6008 1555
rect 5963 1527 5991 1545
tri 5867 1504 5882 1519 ne
tri 5882 1504 5904 1526 sw
rect 5948 1517 5991 1527
rect 6006 1541 6008 1545
rect 6130 1555 6190 1569
tri 6244 1564 6257 1577 ne
rect 6257 1571 6266 1577
tri 6266 1571 6272 1577 sw
rect 6130 1545 6175 1555
rect 6006 1517 6080 1541
rect 5948 1513 6080 1517
tri 6080 1513 6108 1541 sw
rect 6130 1531 6132 1545
tri 6130 1529 6132 1531 ne
rect 6144 1527 6175 1545
rect 6144 1517 6190 1527
rect 6257 1556 6272 1571
tri 5882 1492 5894 1504 ne
rect 5894 1499 5904 1504
tri 5904 1499 5909 1504 sw
rect 5793 1153 5808 1381
rect 5894 1343 5909 1499
rect 5948 1457 5976 1513
tri 6068 1495 6086 1513 ne
rect 6086 1493 6108 1513
tri 6108 1493 6128 1513 sw
tri 6144 1499 6162 1517 ne
rect 5967 1423 5976 1457
rect 6010 1484 6052 1485
rect 6010 1450 6015 1484
rect 6045 1450 6052 1484
rect 6010 1441 6052 1450
rect 6086 1484 6128 1493
rect 6086 1450 6093 1484
rect 6123 1450 6128 1484
rect 6086 1445 6128 1450
rect 6162 1457 6190 1517
tri 6235 1504 6257 1526 se
rect 6257 1519 6272 1527
tri 6257 1504 6272 1519 nw
tri 6229 1498 6235 1504 se
rect 6235 1498 6244 1504
rect 5948 1413 5976 1423
tri 5976 1413 6000 1437 sw
rect 5948 1381 5990 1413
tri 6007 1405 6008 1406 sw
rect 6007 1381 6008 1405
tri 6010 1404 6047 1441 ne
rect 6047 1413 6052 1441
tri 6052 1413 6078 1439 sw
rect 6162 1423 6171 1457
rect 6162 1413 6190 1423
rect 6047 1404 6131 1413
tri 6047 1385 6066 1404 ne
rect 6066 1385 6131 1404
rect 5948 1359 6008 1381
rect 6130 1381 6131 1385
rect 6148 1381 6190 1413
rect 6130 1359 6190 1381
rect 6036 1343 6053 1357
rect 6085 1343 6102 1357
tri 5873 1307 5895 1329 se
rect 5895 1322 5910 1343
tri 5895 1307 5910 1322 nw
rect 6229 1322 6244 1498
tri 6244 1491 6257 1504 nw
rect 6330 1423 6345 1651
tri 5867 1301 5873 1307 se
rect 5873 1301 5882 1307
rect 5867 1285 5882 1301
tri 5882 1294 5895 1307 nw
rect 6036 1299 6053 1313
rect 6085 1299 6102 1313
tri 6229 1307 6244 1322 ne
tri 6244 1307 6266 1329 sw
rect 5867 1249 5882 1257
rect 5948 1285 6008 1299
rect 5963 1275 6008 1285
rect 5963 1257 5991 1275
tri 5867 1234 5882 1249 ne
tri 5882 1234 5904 1256 sw
rect 5948 1247 5991 1257
rect 6006 1271 6008 1275
rect 6130 1285 6190 1299
tri 6244 1294 6257 1307 ne
rect 6257 1301 6266 1307
tri 6266 1301 6272 1307 sw
rect 6130 1275 6175 1285
rect 6006 1247 6080 1271
rect 5948 1243 6080 1247
tri 6080 1243 6108 1271 sw
rect 6130 1261 6132 1275
tri 6130 1259 6132 1261 ne
rect 6144 1257 6175 1275
rect 6144 1247 6190 1257
rect 6257 1286 6272 1301
tri 5882 1222 5894 1234 ne
rect 5894 1229 5904 1234
tri 5904 1229 5909 1234 sw
rect 5793 883 5808 1111
rect 5894 1121 5909 1229
rect 5948 1187 5976 1243
tri 6068 1225 6086 1243 ne
rect 6086 1223 6108 1243
tri 6108 1223 6128 1243 sw
tri 6144 1229 6162 1247 ne
rect 5967 1153 5976 1187
rect 6010 1214 6052 1215
rect 6010 1180 6015 1214
rect 6045 1180 6052 1214
rect 6010 1171 6052 1180
rect 6086 1214 6128 1223
rect 6086 1180 6093 1214
rect 6123 1180 6128 1214
rect 6086 1175 6128 1180
rect 6162 1187 6190 1247
tri 6235 1234 6257 1256 se
rect 6257 1249 6272 1257
tri 6257 1234 6272 1249 nw
tri 6229 1228 6235 1234 se
rect 6235 1228 6244 1234
rect 5948 1143 5976 1153
tri 5976 1143 6000 1167 sw
rect 5894 1073 5910 1121
rect 5948 1111 5990 1143
tri 6007 1135 6008 1136 sw
rect 6007 1111 6008 1135
tri 6010 1134 6047 1171 ne
rect 6047 1143 6052 1171
tri 6052 1143 6078 1169 sw
rect 6162 1153 6171 1187
rect 6162 1143 6190 1153
rect 6047 1134 6131 1143
tri 6047 1115 6066 1134 ne
rect 6066 1115 6131 1134
rect 5948 1089 6008 1111
rect 6130 1111 6131 1115
rect 6148 1111 6190 1143
rect 6130 1089 6190 1111
rect 6036 1073 6053 1087
rect 6085 1073 6102 1087
tri 5873 1037 5895 1059 se
rect 5895 1052 5910 1073
tri 5895 1037 5910 1052 nw
rect 6229 1052 6244 1228
tri 6244 1221 6257 1234 nw
rect 6330 1153 6345 1381
tri 5867 1031 5873 1037 se
rect 5873 1031 5882 1037
rect 5867 1015 5882 1031
tri 5882 1024 5895 1037 nw
rect 6036 1029 6053 1043
rect 6085 1029 6102 1043
tri 6229 1037 6244 1052 ne
tri 6244 1037 6266 1059 sw
rect 5867 979 5882 987
rect 5948 1015 6008 1029
rect 5963 1005 6008 1015
rect 5963 987 5991 1005
tri 5867 964 5882 979 ne
tri 5882 964 5904 986 sw
rect 5948 977 5991 987
rect 6006 1001 6008 1005
rect 6130 1015 6190 1029
tri 6244 1024 6257 1037 ne
rect 6257 1031 6266 1037
tri 6266 1031 6272 1037 sw
rect 6130 1005 6175 1015
rect 6006 977 6080 1001
rect 5948 973 6080 977
tri 6080 973 6108 1001 sw
rect 6130 991 6132 1005
tri 6130 989 6132 991 ne
rect 6144 987 6175 1005
rect 6144 977 6190 987
rect 6257 1016 6272 1031
tri 5882 952 5894 964 ne
rect 5894 959 5904 964
tri 5904 959 5909 964 sw
rect 5793 613 5808 841
rect 5894 803 5909 959
rect 5948 917 5976 973
tri 6068 955 6086 973 ne
rect 6086 953 6108 973
tri 6108 953 6128 973 sw
tri 6144 959 6162 977 ne
rect 5967 883 5976 917
rect 6010 944 6052 945
rect 6010 910 6015 944
rect 6045 910 6052 944
rect 6010 901 6052 910
rect 6086 944 6128 953
rect 6086 910 6093 944
rect 6123 910 6128 944
rect 6086 905 6128 910
rect 6162 917 6190 977
tri 6235 964 6257 986 se
rect 6257 979 6272 987
tri 6257 964 6272 979 nw
tri 6229 958 6235 964 se
rect 6235 958 6244 964
rect 5948 873 5976 883
tri 5976 873 6000 897 sw
rect 5948 841 5990 873
tri 6007 865 6008 866 sw
rect 6007 841 6008 865
tri 6010 864 6047 901 ne
rect 6047 873 6052 901
tri 6052 873 6078 899 sw
rect 6162 883 6171 917
rect 6162 873 6190 883
rect 6047 864 6131 873
tri 6047 845 6066 864 ne
rect 6066 845 6131 864
rect 5948 819 6008 841
rect 6130 841 6131 845
rect 6148 841 6190 873
rect 6130 819 6190 841
rect 6036 803 6053 817
rect 6085 803 6102 817
tri 5873 767 5895 789 se
rect 5895 782 5910 803
tri 5895 767 5910 782 nw
rect 6229 782 6244 958
tri 6244 951 6257 964 nw
rect 6330 883 6345 1111
tri 5867 761 5873 767 se
rect 5873 761 5882 767
rect 5867 745 5882 761
tri 5882 754 5895 767 nw
rect 6036 759 6053 773
rect 6085 759 6102 773
tri 6229 767 6244 782 ne
tri 6244 767 6266 789 sw
rect 5867 709 5882 717
rect 5948 745 6008 759
rect 5963 735 6008 745
rect 5963 717 5991 735
tri 5867 694 5882 709 ne
tri 5882 694 5904 716 sw
rect 5948 707 5991 717
rect 6006 731 6008 735
rect 6130 745 6190 759
tri 6244 754 6257 767 ne
rect 6257 761 6266 767
tri 6266 761 6272 767 sw
rect 6130 735 6175 745
rect 6006 707 6080 731
rect 5948 703 6080 707
tri 6080 703 6108 731 sw
rect 6130 721 6132 735
tri 6130 719 6132 721 ne
rect 6144 717 6175 735
rect 6144 707 6190 717
rect 6257 746 6272 761
tri 5882 682 5894 694 ne
rect 5894 689 5904 694
tri 5904 689 5909 694 sw
rect 5793 343 5808 571
rect 5894 581 5909 689
rect 5948 647 5976 703
tri 6068 685 6086 703 ne
rect 6086 683 6108 703
tri 6108 683 6128 703 sw
tri 6144 689 6162 707 ne
rect 5967 613 5976 647
rect 6010 674 6052 675
rect 6010 640 6015 674
rect 6045 640 6052 674
rect 6010 631 6052 640
rect 6086 674 6128 683
rect 6086 640 6093 674
rect 6123 640 6128 674
rect 6086 635 6128 640
rect 6162 647 6190 707
tri 6235 694 6257 716 se
rect 6257 709 6272 717
tri 6257 694 6272 709 nw
tri 6229 688 6235 694 se
rect 6235 688 6244 694
rect 5948 603 5976 613
tri 5976 603 6000 627 sw
rect 5894 533 5910 581
rect 5948 571 5990 603
tri 6007 595 6008 596 sw
rect 6007 571 6008 595
tri 6010 594 6047 631 ne
rect 6047 603 6052 631
tri 6052 603 6078 629 sw
rect 6162 613 6171 647
rect 6162 603 6190 613
rect 6047 594 6131 603
tri 6047 575 6066 594 ne
rect 6066 575 6131 594
rect 5948 549 6008 571
rect 6130 571 6131 575
rect 6148 571 6190 603
rect 6130 549 6190 571
rect 6036 533 6053 547
rect 6085 533 6102 547
tri 5873 497 5895 519 se
rect 5895 512 5910 533
tri 5895 497 5910 512 nw
rect 6229 512 6244 688
tri 6244 681 6257 694 nw
rect 6330 613 6345 841
tri 5867 491 5873 497 se
rect 5873 491 5882 497
rect 5867 475 5882 491
tri 5882 484 5895 497 nw
rect 6036 489 6053 503
rect 6085 489 6102 503
tri 6229 497 6244 512 ne
tri 6244 497 6266 519 sw
rect 5867 439 5882 447
rect 5948 475 6008 489
rect 5963 465 6008 475
rect 5963 447 5991 465
tri 5867 424 5882 439 ne
tri 5882 424 5904 446 sw
rect 5948 437 5991 447
rect 6006 461 6008 465
rect 6130 475 6190 489
tri 6244 484 6257 497 ne
rect 6257 491 6266 497
tri 6266 491 6272 497 sw
rect 6130 465 6175 475
rect 6006 437 6080 461
rect 5948 433 6080 437
tri 6080 433 6108 461 sw
rect 6130 451 6132 465
tri 6130 449 6132 451 ne
rect 6144 447 6175 465
rect 6144 437 6190 447
rect 6257 476 6272 491
tri 5882 412 5894 424 ne
rect 5894 419 5904 424
tri 5904 419 5909 424 sw
rect 5793 73 5808 301
rect 5894 263 5909 419
rect 5948 377 5976 433
tri 6068 415 6086 433 ne
rect 6086 413 6108 433
tri 6108 413 6128 433 sw
tri 6144 419 6162 437 ne
rect 5967 343 5976 377
rect 6010 404 6052 405
rect 6010 370 6015 404
rect 6045 370 6052 404
rect 6010 361 6052 370
rect 6086 404 6128 413
rect 6086 370 6093 404
rect 6123 370 6128 404
rect 6086 365 6128 370
rect 6162 377 6190 437
tri 6235 424 6257 446 se
rect 6257 439 6272 447
tri 6257 424 6272 439 nw
tri 6229 418 6235 424 se
rect 6235 418 6244 424
rect 5948 333 5976 343
tri 5976 333 6000 357 sw
rect 5948 301 5990 333
tri 6007 325 6008 326 sw
rect 6007 301 6008 325
tri 6010 324 6047 361 ne
rect 6047 333 6052 361
tri 6052 333 6078 359 sw
rect 6162 343 6171 377
rect 6162 333 6190 343
rect 6047 324 6131 333
tri 6047 305 6066 324 ne
rect 6066 305 6131 324
rect 5948 279 6008 301
rect 6130 301 6131 305
rect 6148 301 6190 333
rect 6130 279 6190 301
rect 6036 263 6053 277
rect 6085 263 6102 277
tri 5873 227 5895 249 se
rect 5895 242 5910 263
tri 5895 227 5910 242 nw
rect 6229 242 6244 418
tri 6244 411 6257 424 nw
rect 6330 343 6345 571
tri 5867 221 5873 227 se
rect 5873 221 5882 227
rect 5867 205 5882 221
tri 5882 214 5895 227 nw
rect 6036 219 6053 233
rect 6085 219 6102 233
tri 6229 227 6244 242 ne
tri 6244 227 6266 249 sw
rect 5867 169 5882 177
rect 5948 205 6008 219
rect 5963 195 6008 205
rect 5963 177 5991 195
tri 5867 154 5882 169 ne
tri 5882 154 5904 176 sw
rect 5948 167 5991 177
rect 6006 191 6008 195
rect 6130 205 6190 219
tri 6244 214 6257 227 ne
rect 6257 221 6266 227
tri 6266 221 6272 227 sw
rect 6130 195 6175 205
rect 6006 167 6080 191
rect 5948 163 6080 167
tri 6080 163 6108 191 sw
rect 6130 181 6132 195
tri 6130 179 6132 181 ne
rect 6144 177 6175 195
rect 6144 167 6190 177
rect 6257 206 6272 221
tri 5882 142 5894 154 ne
rect 5894 149 5904 154
tri 5904 149 5909 154 sw
rect 5793 -55 5808 31
rect 5894 -55 5909 149
rect 5948 107 5976 163
tri 6068 145 6086 163 ne
rect 6086 143 6108 163
tri 6108 143 6128 163 sw
tri 6144 149 6162 167 ne
rect 5967 73 5976 107
rect 6010 134 6052 135
rect 6010 100 6015 134
rect 6045 100 6052 134
rect 6010 91 6052 100
rect 6086 134 6128 143
rect 6086 100 6093 134
rect 6123 100 6128 134
rect 6086 95 6128 100
rect 6162 107 6190 167
tri 6235 154 6257 176 se
rect 6257 169 6272 177
tri 6257 154 6272 169 nw
tri 6229 148 6235 154 se
rect 6235 148 6244 154
rect 5948 63 5976 73
tri 5976 63 6000 87 sw
rect 5948 31 5990 63
tri 6007 55 6008 56 sw
rect 6007 31 6008 55
tri 6010 54 6047 91 ne
rect 6047 63 6052 91
tri 6052 63 6078 89 sw
rect 6162 73 6171 107
rect 6162 63 6190 73
rect 6047 54 6131 63
tri 6047 35 6066 54 ne
rect 6066 35 6131 54
rect 5948 9 6008 31
rect 6130 31 6131 35
rect 6148 31 6190 63
rect 6130 9 6190 31
rect 6036 -7 6053 7
rect 6085 -7 6102 7
rect 6229 -55 6244 148
tri 6244 141 6257 154 nw
rect 6330 73 6345 301
rect 6330 -55 6345 31
rect 6373 4123 6388 4361
tri 6453 4277 6475 4299 se
rect 6475 4292 6490 4361
tri 6475 4277 6490 4292 nw
rect 6809 4292 6824 4361
tri 6447 4271 6453 4277 se
rect 6453 4271 6462 4277
rect 6447 4255 6462 4271
tri 6462 4264 6475 4277 nw
rect 6616 4269 6633 4283
rect 6665 4269 6682 4283
tri 6809 4277 6824 4292 ne
tri 6824 4277 6846 4299 sw
rect 6447 4219 6462 4227
rect 6528 4255 6588 4269
rect 6543 4245 6588 4255
rect 6543 4227 6571 4245
tri 6447 4204 6462 4219 ne
tri 6462 4204 6484 4226 sw
rect 6528 4217 6571 4227
rect 6586 4241 6588 4245
rect 6710 4255 6770 4269
tri 6824 4264 6837 4277 ne
rect 6837 4271 6846 4277
tri 6846 4271 6852 4277 sw
rect 6710 4245 6755 4255
rect 6586 4217 6660 4241
rect 6528 4213 6660 4217
tri 6660 4213 6688 4241 sw
rect 6710 4231 6712 4245
tri 6710 4229 6712 4231 ne
rect 6724 4227 6755 4245
rect 6724 4217 6770 4227
rect 6837 4256 6852 4271
tri 6462 4192 6474 4204 ne
rect 6474 4199 6484 4204
tri 6484 4199 6489 4204 sw
rect 6373 3853 6388 4081
rect 6474 4043 6489 4199
rect 6528 4157 6556 4213
tri 6648 4195 6666 4213 ne
rect 6666 4193 6688 4213
tri 6688 4193 6708 4213 sw
tri 6724 4199 6742 4217 ne
rect 6547 4123 6556 4157
rect 6590 4184 6632 4185
rect 6590 4150 6595 4184
rect 6625 4150 6632 4184
rect 6590 4141 6632 4150
rect 6666 4184 6708 4193
rect 6666 4150 6673 4184
rect 6703 4150 6708 4184
rect 6666 4145 6708 4150
rect 6742 4157 6770 4217
tri 6815 4204 6837 4226 se
rect 6837 4219 6852 4227
tri 6837 4204 6852 4219 nw
tri 6809 4198 6815 4204 se
rect 6815 4198 6824 4204
rect 6528 4113 6556 4123
tri 6556 4113 6580 4137 sw
rect 6528 4081 6570 4113
tri 6587 4105 6588 4106 sw
rect 6587 4081 6588 4105
tri 6590 4104 6627 4141 ne
rect 6627 4113 6632 4141
tri 6632 4113 6658 4139 sw
rect 6742 4123 6751 4157
rect 6742 4113 6770 4123
rect 6627 4104 6711 4113
tri 6627 4085 6646 4104 ne
rect 6646 4085 6711 4104
rect 6528 4059 6588 4081
rect 6710 4081 6711 4085
rect 6728 4081 6770 4113
rect 6710 4059 6770 4081
rect 6616 4043 6633 4057
rect 6665 4043 6682 4057
tri 6453 4007 6475 4029 se
rect 6475 4022 6490 4043
tri 6475 4007 6490 4022 nw
rect 6809 4022 6824 4198
tri 6824 4191 6837 4204 nw
rect 6910 4123 6925 4361
tri 6447 4001 6453 4007 se
rect 6453 4001 6462 4007
rect 6447 3985 6462 4001
tri 6462 3994 6475 4007 nw
rect 6616 3999 6633 4013
rect 6665 3999 6682 4013
tri 6809 4007 6824 4022 ne
tri 6824 4007 6846 4029 sw
rect 6447 3949 6462 3957
rect 6528 3985 6588 3999
rect 6543 3975 6588 3985
rect 6543 3957 6571 3975
tri 6447 3934 6462 3949 ne
tri 6462 3934 6484 3956 sw
rect 6528 3947 6571 3957
rect 6586 3971 6588 3975
rect 6710 3985 6770 3999
tri 6824 3994 6837 4007 ne
rect 6837 4001 6846 4007
tri 6846 4001 6852 4007 sw
rect 6710 3975 6755 3985
rect 6586 3947 6660 3971
rect 6528 3943 6660 3947
tri 6660 3943 6688 3971 sw
rect 6710 3961 6712 3975
tri 6710 3959 6712 3961 ne
rect 6724 3957 6755 3975
rect 6724 3947 6770 3957
rect 6837 3986 6852 4001
tri 6462 3922 6474 3934 ne
rect 6474 3929 6484 3934
tri 6484 3929 6489 3934 sw
rect 6373 3583 6388 3811
rect 6474 3821 6489 3929
rect 6528 3887 6556 3943
tri 6648 3925 6666 3943 ne
rect 6666 3923 6688 3943
tri 6688 3923 6708 3943 sw
tri 6724 3929 6742 3947 ne
rect 6547 3853 6556 3887
rect 6590 3914 6632 3915
rect 6590 3880 6595 3914
rect 6625 3880 6632 3914
rect 6590 3871 6632 3880
rect 6666 3914 6708 3923
rect 6666 3880 6673 3914
rect 6703 3880 6708 3914
rect 6666 3875 6708 3880
rect 6742 3887 6770 3947
tri 6815 3934 6837 3956 se
rect 6837 3949 6852 3957
tri 6837 3934 6852 3949 nw
tri 6809 3928 6815 3934 se
rect 6815 3928 6824 3934
rect 6528 3843 6556 3853
tri 6556 3843 6580 3867 sw
rect 6474 3773 6490 3821
rect 6528 3811 6570 3843
tri 6587 3835 6588 3836 sw
rect 6587 3811 6588 3835
tri 6590 3834 6627 3871 ne
rect 6627 3843 6632 3871
tri 6632 3843 6658 3869 sw
rect 6742 3853 6751 3887
rect 6742 3843 6770 3853
rect 6627 3834 6711 3843
tri 6627 3815 6646 3834 ne
rect 6646 3815 6711 3834
rect 6528 3789 6588 3811
rect 6710 3811 6711 3815
rect 6728 3811 6770 3843
rect 6710 3789 6770 3811
rect 6616 3773 6633 3787
rect 6665 3773 6682 3787
tri 6453 3737 6475 3759 se
rect 6475 3752 6490 3773
tri 6475 3737 6490 3752 nw
rect 6809 3752 6824 3928
tri 6824 3921 6837 3934 nw
rect 6910 3853 6925 4081
tri 6447 3731 6453 3737 se
rect 6453 3731 6462 3737
rect 6447 3715 6462 3731
tri 6462 3724 6475 3737 nw
rect 6616 3729 6633 3743
rect 6665 3729 6682 3743
tri 6809 3737 6824 3752 ne
tri 6824 3737 6846 3759 sw
rect 6447 3679 6462 3687
rect 6528 3715 6588 3729
rect 6543 3705 6588 3715
rect 6543 3687 6571 3705
tri 6447 3664 6462 3679 ne
tri 6462 3664 6484 3686 sw
rect 6528 3677 6571 3687
rect 6586 3701 6588 3705
rect 6710 3715 6770 3729
tri 6824 3724 6837 3737 ne
rect 6837 3731 6846 3737
tri 6846 3731 6852 3737 sw
rect 6710 3705 6755 3715
rect 6586 3677 6660 3701
rect 6528 3673 6660 3677
tri 6660 3673 6688 3701 sw
rect 6710 3691 6712 3705
tri 6710 3689 6712 3691 ne
rect 6724 3687 6755 3705
rect 6724 3677 6770 3687
rect 6837 3716 6852 3731
tri 6462 3652 6474 3664 ne
rect 6474 3659 6484 3664
tri 6484 3659 6489 3664 sw
rect 6373 3313 6388 3541
rect 6474 3503 6489 3659
rect 6528 3617 6556 3673
tri 6648 3655 6666 3673 ne
rect 6666 3653 6688 3673
tri 6688 3653 6708 3673 sw
tri 6724 3659 6742 3677 ne
rect 6547 3583 6556 3617
rect 6590 3644 6632 3645
rect 6590 3610 6595 3644
rect 6625 3610 6632 3644
rect 6590 3601 6632 3610
rect 6666 3644 6708 3653
rect 6666 3610 6673 3644
rect 6703 3610 6708 3644
rect 6666 3605 6708 3610
rect 6742 3617 6770 3677
tri 6815 3664 6837 3686 se
rect 6837 3679 6852 3687
tri 6837 3664 6852 3679 nw
tri 6809 3658 6815 3664 se
rect 6815 3658 6824 3664
rect 6528 3573 6556 3583
tri 6556 3573 6580 3597 sw
rect 6528 3541 6570 3573
tri 6587 3565 6588 3566 sw
rect 6587 3541 6588 3565
tri 6590 3564 6627 3601 ne
rect 6627 3573 6632 3601
tri 6632 3573 6658 3599 sw
rect 6742 3583 6751 3617
rect 6742 3573 6770 3583
rect 6627 3564 6711 3573
tri 6627 3545 6646 3564 ne
rect 6646 3545 6711 3564
rect 6528 3519 6588 3541
rect 6710 3541 6711 3545
rect 6728 3541 6770 3573
rect 6710 3519 6770 3541
rect 6616 3503 6633 3517
rect 6665 3503 6682 3517
tri 6453 3467 6475 3489 se
rect 6475 3482 6490 3503
tri 6475 3467 6490 3482 nw
rect 6809 3482 6824 3658
tri 6824 3651 6837 3664 nw
rect 6910 3583 6925 3811
tri 6447 3461 6453 3467 se
rect 6453 3461 6462 3467
rect 6447 3445 6462 3461
tri 6462 3454 6475 3467 nw
rect 6616 3459 6633 3473
rect 6665 3459 6682 3473
tri 6809 3467 6824 3482 ne
tri 6824 3467 6846 3489 sw
rect 6447 3409 6462 3417
rect 6528 3445 6588 3459
rect 6543 3435 6588 3445
rect 6543 3417 6571 3435
tri 6447 3394 6462 3409 ne
tri 6462 3394 6484 3416 sw
rect 6528 3407 6571 3417
rect 6586 3431 6588 3435
rect 6710 3445 6770 3459
tri 6824 3454 6837 3467 ne
rect 6837 3461 6846 3467
tri 6846 3461 6852 3467 sw
rect 6710 3435 6755 3445
rect 6586 3407 6660 3431
rect 6528 3403 6660 3407
tri 6660 3403 6688 3431 sw
rect 6710 3421 6712 3435
tri 6710 3419 6712 3421 ne
rect 6724 3417 6755 3435
rect 6724 3407 6770 3417
rect 6837 3446 6852 3461
tri 6462 3382 6474 3394 ne
rect 6474 3389 6484 3394
tri 6484 3389 6489 3394 sw
rect 6373 3043 6388 3271
rect 6474 3281 6489 3389
rect 6528 3347 6556 3403
tri 6648 3385 6666 3403 ne
rect 6666 3383 6688 3403
tri 6688 3383 6708 3403 sw
tri 6724 3389 6742 3407 ne
rect 6547 3313 6556 3347
rect 6590 3374 6632 3375
rect 6590 3340 6595 3374
rect 6625 3340 6632 3374
rect 6590 3331 6632 3340
rect 6666 3374 6708 3383
rect 6666 3340 6673 3374
rect 6703 3340 6708 3374
rect 6666 3335 6708 3340
rect 6742 3347 6770 3407
tri 6815 3394 6837 3416 se
rect 6837 3409 6852 3417
tri 6837 3394 6852 3409 nw
tri 6809 3388 6815 3394 se
rect 6815 3388 6824 3394
rect 6528 3303 6556 3313
tri 6556 3303 6580 3327 sw
rect 6474 3233 6490 3281
rect 6528 3271 6570 3303
tri 6587 3295 6588 3296 sw
rect 6587 3271 6588 3295
tri 6590 3294 6627 3331 ne
rect 6627 3303 6632 3331
tri 6632 3303 6658 3329 sw
rect 6742 3313 6751 3347
rect 6742 3303 6770 3313
rect 6627 3294 6711 3303
tri 6627 3275 6646 3294 ne
rect 6646 3275 6711 3294
rect 6528 3249 6588 3271
rect 6710 3271 6711 3275
rect 6728 3271 6770 3303
rect 6710 3249 6770 3271
rect 6616 3233 6633 3247
rect 6665 3233 6682 3247
tri 6453 3197 6475 3219 se
rect 6475 3212 6490 3233
tri 6475 3197 6490 3212 nw
rect 6809 3212 6824 3388
tri 6824 3381 6837 3394 nw
rect 6910 3313 6925 3541
tri 6447 3191 6453 3197 se
rect 6453 3191 6462 3197
rect 6447 3175 6462 3191
tri 6462 3184 6475 3197 nw
rect 6616 3189 6633 3203
rect 6665 3189 6682 3203
tri 6809 3197 6824 3212 ne
tri 6824 3197 6846 3219 sw
rect 6447 3139 6462 3147
rect 6528 3175 6588 3189
rect 6543 3165 6588 3175
rect 6543 3147 6571 3165
tri 6447 3124 6462 3139 ne
tri 6462 3124 6484 3146 sw
rect 6528 3137 6571 3147
rect 6586 3161 6588 3165
rect 6710 3175 6770 3189
tri 6824 3184 6837 3197 ne
rect 6837 3191 6846 3197
tri 6846 3191 6852 3197 sw
rect 6710 3165 6755 3175
rect 6586 3137 6660 3161
rect 6528 3133 6660 3137
tri 6660 3133 6688 3161 sw
rect 6710 3151 6712 3165
tri 6710 3149 6712 3151 ne
rect 6724 3147 6755 3165
rect 6724 3137 6770 3147
rect 6837 3176 6852 3191
tri 6462 3112 6474 3124 ne
rect 6474 3119 6484 3124
tri 6484 3119 6489 3124 sw
rect 6373 2773 6388 3001
rect 6474 2963 6489 3119
rect 6528 3077 6556 3133
tri 6648 3115 6666 3133 ne
rect 6666 3113 6688 3133
tri 6688 3113 6708 3133 sw
tri 6724 3119 6742 3137 ne
rect 6547 3043 6556 3077
rect 6590 3104 6632 3105
rect 6590 3070 6595 3104
rect 6625 3070 6632 3104
rect 6590 3061 6632 3070
rect 6666 3104 6708 3113
rect 6666 3070 6673 3104
rect 6703 3070 6708 3104
rect 6666 3065 6708 3070
rect 6742 3077 6770 3137
tri 6815 3124 6837 3146 se
rect 6837 3139 6852 3147
tri 6837 3124 6852 3139 nw
tri 6809 3118 6815 3124 se
rect 6815 3118 6824 3124
rect 6528 3033 6556 3043
tri 6556 3033 6580 3057 sw
rect 6528 3001 6570 3033
tri 6587 3025 6588 3026 sw
rect 6587 3001 6588 3025
tri 6590 3024 6627 3061 ne
rect 6627 3033 6632 3061
tri 6632 3033 6658 3059 sw
rect 6742 3043 6751 3077
rect 6742 3033 6770 3043
rect 6627 3024 6711 3033
tri 6627 3005 6646 3024 ne
rect 6646 3005 6711 3024
rect 6528 2979 6588 3001
rect 6710 3001 6711 3005
rect 6728 3001 6770 3033
rect 6710 2979 6770 3001
rect 6616 2963 6633 2977
rect 6665 2963 6682 2977
tri 6453 2927 6475 2949 se
rect 6475 2942 6490 2963
tri 6475 2927 6490 2942 nw
rect 6809 2942 6824 3118
tri 6824 3111 6837 3124 nw
rect 6910 3043 6925 3271
tri 6447 2921 6453 2927 se
rect 6453 2921 6462 2927
rect 6447 2905 6462 2921
tri 6462 2914 6475 2927 nw
rect 6616 2919 6633 2933
rect 6665 2919 6682 2933
tri 6809 2927 6824 2942 ne
tri 6824 2927 6846 2949 sw
rect 6447 2869 6462 2877
rect 6528 2905 6588 2919
rect 6543 2895 6588 2905
rect 6543 2877 6571 2895
tri 6447 2854 6462 2869 ne
tri 6462 2854 6484 2876 sw
rect 6528 2867 6571 2877
rect 6586 2891 6588 2895
rect 6710 2905 6770 2919
tri 6824 2914 6837 2927 ne
rect 6837 2921 6846 2927
tri 6846 2921 6852 2927 sw
rect 6710 2895 6755 2905
rect 6586 2867 6660 2891
rect 6528 2863 6660 2867
tri 6660 2863 6688 2891 sw
rect 6710 2881 6712 2895
tri 6710 2879 6712 2881 ne
rect 6724 2877 6755 2895
rect 6724 2867 6770 2877
rect 6837 2906 6852 2921
tri 6462 2842 6474 2854 ne
rect 6474 2849 6484 2854
tri 6484 2849 6489 2854 sw
rect 6373 2503 6388 2731
rect 6474 2741 6489 2849
rect 6528 2807 6556 2863
tri 6648 2845 6666 2863 ne
rect 6666 2843 6688 2863
tri 6688 2843 6708 2863 sw
tri 6724 2849 6742 2867 ne
rect 6547 2773 6556 2807
rect 6590 2834 6632 2835
rect 6590 2800 6595 2834
rect 6625 2800 6632 2834
rect 6590 2791 6632 2800
rect 6666 2834 6708 2843
rect 6666 2800 6673 2834
rect 6703 2800 6708 2834
rect 6666 2795 6708 2800
rect 6742 2807 6770 2867
tri 6815 2854 6837 2876 se
rect 6837 2869 6852 2877
tri 6837 2854 6852 2869 nw
tri 6809 2848 6815 2854 se
rect 6815 2848 6824 2854
rect 6528 2763 6556 2773
tri 6556 2763 6580 2787 sw
rect 6474 2693 6490 2741
rect 6528 2731 6570 2763
tri 6587 2755 6588 2756 sw
rect 6587 2731 6588 2755
tri 6590 2754 6627 2791 ne
rect 6627 2763 6632 2791
tri 6632 2763 6658 2789 sw
rect 6742 2773 6751 2807
rect 6742 2763 6770 2773
rect 6627 2754 6711 2763
tri 6627 2735 6646 2754 ne
rect 6646 2735 6711 2754
rect 6528 2709 6588 2731
rect 6710 2731 6711 2735
rect 6728 2731 6770 2763
rect 6710 2709 6770 2731
rect 6616 2693 6633 2707
rect 6665 2693 6682 2707
tri 6453 2657 6475 2679 se
rect 6475 2672 6490 2693
tri 6475 2657 6490 2672 nw
rect 6809 2672 6824 2848
tri 6824 2841 6837 2854 nw
rect 6910 2773 6925 3001
tri 6447 2651 6453 2657 se
rect 6453 2651 6462 2657
rect 6447 2635 6462 2651
tri 6462 2644 6475 2657 nw
rect 6616 2649 6633 2663
rect 6665 2649 6682 2663
tri 6809 2657 6824 2672 ne
tri 6824 2657 6846 2679 sw
rect 6447 2599 6462 2607
rect 6528 2635 6588 2649
rect 6543 2625 6588 2635
rect 6543 2607 6571 2625
tri 6447 2584 6462 2599 ne
tri 6462 2584 6484 2606 sw
rect 6528 2597 6571 2607
rect 6586 2621 6588 2625
rect 6710 2635 6770 2649
tri 6824 2644 6837 2657 ne
rect 6837 2651 6846 2657
tri 6846 2651 6852 2657 sw
rect 6710 2625 6755 2635
rect 6586 2597 6660 2621
rect 6528 2593 6660 2597
tri 6660 2593 6688 2621 sw
rect 6710 2611 6712 2625
tri 6710 2609 6712 2611 ne
rect 6724 2607 6755 2625
rect 6724 2597 6770 2607
rect 6837 2636 6852 2651
tri 6462 2572 6474 2584 ne
rect 6474 2579 6484 2584
tri 6484 2579 6489 2584 sw
rect 6373 2233 6388 2461
rect 6474 2423 6489 2579
rect 6528 2537 6556 2593
tri 6648 2575 6666 2593 ne
rect 6666 2573 6688 2593
tri 6688 2573 6708 2593 sw
tri 6724 2579 6742 2597 ne
rect 6547 2503 6556 2537
rect 6590 2564 6632 2565
rect 6590 2530 6595 2564
rect 6625 2530 6632 2564
rect 6590 2521 6632 2530
rect 6666 2564 6708 2573
rect 6666 2530 6673 2564
rect 6703 2530 6708 2564
rect 6666 2525 6708 2530
rect 6742 2537 6770 2597
tri 6815 2584 6837 2606 se
rect 6837 2599 6852 2607
tri 6837 2584 6852 2599 nw
tri 6809 2578 6815 2584 se
rect 6815 2578 6824 2584
rect 6528 2493 6556 2503
tri 6556 2493 6580 2517 sw
rect 6528 2461 6570 2493
tri 6587 2485 6588 2486 sw
rect 6587 2461 6588 2485
tri 6590 2484 6627 2521 ne
rect 6627 2493 6632 2521
tri 6632 2493 6658 2519 sw
rect 6742 2503 6751 2537
rect 6742 2493 6770 2503
rect 6627 2484 6711 2493
tri 6627 2465 6646 2484 ne
rect 6646 2465 6711 2484
rect 6528 2439 6588 2461
rect 6710 2461 6711 2465
rect 6728 2461 6770 2493
rect 6710 2439 6770 2461
rect 6616 2423 6633 2437
rect 6665 2423 6682 2437
tri 6453 2387 6475 2409 se
rect 6475 2402 6490 2423
tri 6475 2387 6490 2402 nw
rect 6809 2402 6824 2578
tri 6824 2571 6837 2584 nw
rect 6910 2503 6925 2731
tri 6447 2381 6453 2387 se
rect 6453 2381 6462 2387
rect 6447 2365 6462 2381
tri 6462 2374 6475 2387 nw
rect 6616 2379 6633 2393
rect 6665 2379 6682 2393
tri 6809 2387 6824 2402 ne
tri 6824 2387 6846 2409 sw
rect 6447 2329 6462 2337
rect 6528 2365 6588 2379
rect 6543 2355 6588 2365
rect 6543 2337 6571 2355
tri 6447 2314 6462 2329 ne
tri 6462 2314 6484 2336 sw
rect 6528 2327 6571 2337
rect 6586 2351 6588 2355
rect 6710 2365 6770 2379
tri 6824 2374 6837 2387 ne
rect 6837 2381 6846 2387
tri 6846 2381 6852 2387 sw
rect 6710 2355 6755 2365
rect 6586 2327 6660 2351
rect 6528 2323 6660 2327
tri 6660 2323 6688 2351 sw
rect 6710 2341 6712 2355
tri 6710 2339 6712 2341 ne
rect 6724 2337 6755 2355
rect 6724 2327 6770 2337
rect 6837 2366 6852 2381
tri 6462 2302 6474 2314 ne
rect 6474 2309 6484 2314
tri 6484 2309 6489 2314 sw
rect 6373 1963 6388 2191
rect 6474 2201 6489 2309
rect 6528 2267 6556 2323
tri 6648 2305 6666 2323 ne
rect 6666 2303 6688 2323
tri 6688 2303 6708 2323 sw
tri 6724 2309 6742 2327 ne
rect 6547 2233 6556 2267
rect 6590 2294 6632 2295
rect 6590 2260 6595 2294
rect 6625 2260 6632 2294
rect 6590 2251 6632 2260
rect 6666 2294 6708 2303
rect 6666 2260 6673 2294
rect 6703 2260 6708 2294
rect 6666 2255 6708 2260
rect 6742 2267 6770 2327
tri 6815 2314 6837 2336 se
rect 6837 2329 6852 2337
tri 6837 2314 6852 2329 nw
tri 6809 2308 6815 2314 se
rect 6815 2308 6824 2314
rect 6528 2223 6556 2233
tri 6556 2223 6580 2247 sw
rect 6474 2153 6490 2201
rect 6528 2191 6570 2223
tri 6587 2215 6588 2216 sw
rect 6587 2191 6588 2215
tri 6590 2214 6627 2251 ne
rect 6627 2223 6632 2251
tri 6632 2223 6658 2249 sw
rect 6742 2233 6751 2267
rect 6742 2223 6770 2233
rect 6627 2214 6711 2223
tri 6627 2195 6646 2214 ne
rect 6646 2195 6711 2214
rect 6528 2169 6588 2191
rect 6710 2191 6711 2195
rect 6728 2191 6770 2223
rect 6710 2169 6770 2191
rect 6616 2153 6633 2167
rect 6665 2153 6682 2167
tri 6453 2117 6475 2139 se
rect 6475 2132 6490 2153
tri 6475 2117 6490 2132 nw
rect 6809 2132 6824 2308
tri 6824 2301 6837 2314 nw
rect 6910 2233 6925 2461
tri 6447 2111 6453 2117 se
rect 6453 2111 6462 2117
rect 6447 2095 6462 2111
tri 6462 2104 6475 2117 nw
rect 6616 2109 6633 2123
rect 6665 2109 6682 2123
tri 6809 2117 6824 2132 ne
tri 6824 2117 6846 2139 sw
rect 6447 2059 6462 2067
rect 6528 2095 6588 2109
rect 6543 2085 6588 2095
rect 6543 2067 6571 2085
tri 6447 2044 6462 2059 ne
tri 6462 2044 6484 2066 sw
rect 6528 2057 6571 2067
rect 6586 2081 6588 2085
rect 6710 2095 6770 2109
tri 6824 2104 6837 2117 ne
rect 6837 2111 6846 2117
tri 6846 2111 6852 2117 sw
rect 6710 2085 6755 2095
rect 6586 2057 6660 2081
rect 6528 2053 6660 2057
tri 6660 2053 6688 2081 sw
rect 6710 2071 6712 2085
tri 6710 2069 6712 2071 ne
rect 6724 2067 6755 2085
rect 6724 2057 6770 2067
rect 6837 2096 6852 2111
tri 6462 2032 6474 2044 ne
rect 6474 2039 6484 2044
tri 6484 2039 6489 2044 sw
rect 6373 1693 6388 1921
rect 6474 1883 6489 2039
rect 6528 1997 6556 2053
tri 6648 2035 6666 2053 ne
rect 6666 2033 6688 2053
tri 6688 2033 6708 2053 sw
tri 6724 2039 6742 2057 ne
rect 6547 1963 6556 1997
rect 6590 2024 6632 2025
rect 6590 1990 6595 2024
rect 6625 1990 6632 2024
rect 6590 1981 6632 1990
rect 6666 2024 6708 2033
rect 6666 1990 6673 2024
rect 6703 1990 6708 2024
rect 6666 1985 6708 1990
rect 6742 1997 6770 2057
tri 6815 2044 6837 2066 se
rect 6837 2059 6852 2067
tri 6837 2044 6852 2059 nw
tri 6809 2038 6815 2044 se
rect 6815 2038 6824 2044
rect 6528 1953 6556 1963
tri 6556 1953 6580 1977 sw
rect 6528 1921 6570 1953
tri 6587 1945 6588 1946 sw
rect 6587 1921 6588 1945
tri 6590 1944 6627 1981 ne
rect 6627 1953 6632 1981
tri 6632 1953 6658 1979 sw
rect 6742 1963 6751 1997
rect 6742 1953 6770 1963
rect 6627 1944 6711 1953
tri 6627 1925 6646 1944 ne
rect 6646 1925 6711 1944
rect 6528 1899 6588 1921
rect 6710 1921 6711 1925
rect 6728 1921 6770 1953
rect 6710 1899 6770 1921
rect 6616 1883 6633 1897
rect 6665 1883 6682 1897
tri 6453 1847 6475 1869 se
rect 6475 1862 6490 1883
tri 6475 1847 6490 1862 nw
rect 6809 1862 6824 2038
tri 6824 2031 6837 2044 nw
rect 6910 1963 6925 2191
tri 6447 1841 6453 1847 se
rect 6453 1841 6462 1847
rect 6447 1825 6462 1841
tri 6462 1834 6475 1847 nw
rect 6616 1839 6633 1853
rect 6665 1839 6682 1853
tri 6809 1847 6824 1862 ne
tri 6824 1847 6846 1869 sw
rect 6447 1789 6462 1797
rect 6528 1825 6588 1839
rect 6543 1815 6588 1825
rect 6543 1797 6571 1815
tri 6447 1774 6462 1789 ne
tri 6462 1774 6484 1796 sw
rect 6528 1787 6571 1797
rect 6586 1811 6588 1815
rect 6710 1825 6770 1839
tri 6824 1834 6837 1847 ne
rect 6837 1841 6846 1847
tri 6846 1841 6852 1847 sw
rect 6710 1815 6755 1825
rect 6586 1787 6660 1811
rect 6528 1783 6660 1787
tri 6660 1783 6688 1811 sw
rect 6710 1801 6712 1815
tri 6710 1799 6712 1801 ne
rect 6724 1797 6755 1815
rect 6724 1787 6770 1797
rect 6837 1826 6852 1841
tri 6462 1762 6474 1774 ne
rect 6474 1769 6484 1774
tri 6484 1769 6489 1774 sw
rect 6373 1423 6388 1651
rect 6474 1661 6489 1769
rect 6528 1727 6556 1783
tri 6648 1765 6666 1783 ne
rect 6666 1763 6688 1783
tri 6688 1763 6708 1783 sw
tri 6724 1769 6742 1787 ne
rect 6547 1693 6556 1727
rect 6590 1754 6632 1755
rect 6590 1720 6595 1754
rect 6625 1720 6632 1754
rect 6590 1711 6632 1720
rect 6666 1754 6708 1763
rect 6666 1720 6673 1754
rect 6703 1720 6708 1754
rect 6666 1715 6708 1720
rect 6742 1727 6770 1787
tri 6815 1774 6837 1796 se
rect 6837 1789 6852 1797
tri 6837 1774 6852 1789 nw
tri 6809 1768 6815 1774 se
rect 6815 1768 6824 1774
rect 6528 1683 6556 1693
tri 6556 1683 6580 1707 sw
rect 6474 1613 6490 1661
rect 6528 1651 6570 1683
tri 6587 1675 6588 1676 sw
rect 6587 1651 6588 1675
tri 6590 1674 6627 1711 ne
rect 6627 1683 6632 1711
tri 6632 1683 6658 1709 sw
rect 6742 1693 6751 1727
rect 6742 1683 6770 1693
rect 6627 1674 6711 1683
tri 6627 1655 6646 1674 ne
rect 6646 1655 6711 1674
rect 6528 1629 6588 1651
rect 6710 1651 6711 1655
rect 6728 1651 6770 1683
rect 6710 1629 6770 1651
rect 6616 1613 6633 1627
rect 6665 1613 6682 1627
tri 6453 1577 6475 1599 se
rect 6475 1592 6490 1613
tri 6475 1577 6490 1592 nw
rect 6809 1592 6824 1768
tri 6824 1761 6837 1774 nw
rect 6910 1693 6925 1921
tri 6447 1571 6453 1577 se
rect 6453 1571 6462 1577
rect 6447 1555 6462 1571
tri 6462 1564 6475 1577 nw
rect 6616 1569 6633 1583
rect 6665 1569 6682 1583
tri 6809 1577 6824 1592 ne
tri 6824 1577 6846 1599 sw
rect 6447 1519 6462 1527
rect 6528 1555 6588 1569
rect 6543 1545 6588 1555
rect 6543 1527 6571 1545
tri 6447 1504 6462 1519 ne
tri 6462 1504 6484 1526 sw
rect 6528 1517 6571 1527
rect 6586 1541 6588 1545
rect 6710 1555 6770 1569
tri 6824 1564 6837 1577 ne
rect 6837 1571 6846 1577
tri 6846 1571 6852 1577 sw
rect 6710 1545 6755 1555
rect 6586 1517 6660 1541
rect 6528 1513 6660 1517
tri 6660 1513 6688 1541 sw
rect 6710 1531 6712 1545
tri 6710 1529 6712 1531 ne
rect 6724 1527 6755 1545
rect 6724 1517 6770 1527
rect 6837 1556 6852 1571
tri 6462 1492 6474 1504 ne
rect 6474 1499 6484 1504
tri 6484 1499 6489 1504 sw
rect 6373 1153 6388 1381
rect 6474 1343 6489 1499
rect 6528 1457 6556 1513
tri 6648 1495 6666 1513 ne
rect 6666 1493 6688 1513
tri 6688 1493 6708 1513 sw
tri 6724 1499 6742 1517 ne
rect 6547 1423 6556 1457
rect 6590 1484 6632 1485
rect 6590 1450 6595 1484
rect 6625 1450 6632 1484
rect 6590 1441 6632 1450
rect 6666 1484 6708 1493
rect 6666 1450 6673 1484
rect 6703 1450 6708 1484
rect 6666 1445 6708 1450
rect 6742 1457 6770 1517
tri 6815 1504 6837 1526 se
rect 6837 1519 6852 1527
tri 6837 1504 6852 1519 nw
tri 6809 1498 6815 1504 se
rect 6815 1498 6824 1504
rect 6528 1413 6556 1423
tri 6556 1413 6580 1437 sw
rect 6528 1381 6570 1413
tri 6587 1405 6588 1406 sw
rect 6587 1381 6588 1405
tri 6590 1404 6627 1441 ne
rect 6627 1413 6632 1441
tri 6632 1413 6658 1439 sw
rect 6742 1423 6751 1457
rect 6742 1413 6770 1423
rect 6627 1404 6711 1413
tri 6627 1385 6646 1404 ne
rect 6646 1385 6711 1404
rect 6528 1359 6588 1381
rect 6710 1381 6711 1385
rect 6728 1381 6770 1413
rect 6710 1359 6770 1381
rect 6616 1343 6633 1357
rect 6665 1343 6682 1357
tri 6453 1307 6475 1329 se
rect 6475 1322 6490 1343
tri 6475 1307 6490 1322 nw
rect 6809 1322 6824 1498
tri 6824 1491 6837 1504 nw
rect 6910 1423 6925 1651
tri 6447 1301 6453 1307 se
rect 6453 1301 6462 1307
rect 6447 1285 6462 1301
tri 6462 1294 6475 1307 nw
rect 6616 1299 6633 1313
rect 6665 1299 6682 1313
tri 6809 1307 6824 1322 ne
tri 6824 1307 6846 1329 sw
rect 6447 1249 6462 1257
rect 6528 1285 6588 1299
rect 6543 1275 6588 1285
rect 6543 1257 6571 1275
tri 6447 1234 6462 1249 ne
tri 6462 1234 6484 1256 sw
rect 6528 1247 6571 1257
rect 6586 1271 6588 1275
rect 6710 1285 6770 1299
tri 6824 1294 6837 1307 ne
rect 6837 1301 6846 1307
tri 6846 1301 6852 1307 sw
rect 6710 1275 6755 1285
rect 6586 1247 6660 1271
rect 6528 1243 6660 1247
tri 6660 1243 6688 1271 sw
rect 6710 1261 6712 1275
tri 6710 1259 6712 1261 ne
rect 6724 1257 6755 1275
rect 6724 1247 6770 1257
rect 6837 1286 6852 1301
tri 6462 1222 6474 1234 ne
rect 6474 1229 6484 1234
tri 6484 1229 6489 1234 sw
rect 6373 883 6388 1111
rect 6474 1121 6489 1229
rect 6528 1187 6556 1243
tri 6648 1225 6666 1243 ne
rect 6666 1223 6688 1243
tri 6688 1223 6708 1243 sw
tri 6724 1229 6742 1247 ne
rect 6547 1153 6556 1187
rect 6590 1214 6632 1215
rect 6590 1180 6595 1214
rect 6625 1180 6632 1214
rect 6590 1171 6632 1180
rect 6666 1214 6708 1223
rect 6666 1180 6673 1214
rect 6703 1180 6708 1214
rect 6666 1175 6708 1180
rect 6742 1187 6770 1247
tri 6815 1234 6837 1256 se
rect 6837 1249 6852 1257
tri 6837 1234 6852 1249 nw
tri 6809 1228 6815 1234 se
rect 6815 1228 6824 1234
rect 6528 1143 6556 1153
tri 6556 1143 6580 1167 sw
rect 6474 1073 6490 1121
rect 6528 1111 6570 1143
tri 6587 1135 6588 1136 sw
rect 6587 1111 6588 1135
tri 6590 1134 6627 1171 ne
rect 6627 1143 6632 1171
tri 6632 1143 6658 1169 sw
rect 6742 1153 6751 1187
rect 6742 1143 6770 1153
rect 6627 1134 6711 1143
tri 6627 1115 6646 1134 ne
rect 6646 1115 6711 1134
rect 6528 1089 6588 1111
rect 6710 1111 6711 1115
rect 6728 1111 6770 1143
rect 6710 1089 6770 1111
rect 6616 1073 6633 1087
rect 6665 1073 6682 1087
tri 6453 1037 6475 1059 se
rect 6475 1052 6490 1073
tri 6475 1037 6490 1052 nw
rect 6809 1052 6824 1228
tri 6824 1221 6837 1234 nw
rect 6910 1153 6925 1381
tri 6447 1031 6453 1037 se
rect 6453 1031 6462 1037
rect 6447 1015 6462 1031
tri 6462 1024 6475 1037 nw
rect 6616 1029 6633 1043
rect 6665 1029 6682 1043
tri 6809 1037 6824 1052 ne
tri 6824 1037 6846 1059 sw
rect 6447 979 6462 987
rect 6528 1015 6588 1029
rect 6543 1005 6588 1015
rect 6543 987 6571 1005
tri 6447 964 6462 979 ne
tri 6462 964 6484 986 sw
rect 6528 977 6571 987
rect 6586 1001 6588 1005
rect 6710 1015 6770 1029
tri 6824 1024 6837 1037 ne
rect 6837 1031 6846 1037
tri 6846 1031 6852 1037 sw
rect 6710 1005 6755 1015
rect 6586 977 6660 1001
rect 6528 973 6660 977
tri 6660 973 6688 1001 sw
rect 6710 991 6712 1005
tri 6710 989 6712 991 ne
rect 6724 987 6755 1005
rect 6724 977 6770 987
rect 6837 1016 6852 1031
tri 6462 952 6474 964 ne
rect 6474 959 6484 964
tri 6484 959 6489 964 sw
rect 6373 613 6388 841
rect 6474 803 6489 959
rect 6528 917 6556 973
tri 6648 955 6666 973 ne
rect 6666 953 6688 973
tri 6688 953 6708 973 sw
tri 6724 959 6742 977 ne
rect 6547 883 6556 917
rect 6590 944 6632 945
rect 6590 910 6595 944
rect 6625 910 6632 944
rect 6590 901 6632 910
rect 6666 944 6708 953
rect 6666 910 6673 944
rect 6703 910 6708 944
rect 6666 905 6708 910
rect 6742 917 6770 977
tri 6815 964 6837 986 se
rect 6837 979 6852 987
tri 6837 964 6852 979 nw
tri 6809 958 6815 964 se
rect 6815 958 6824 964
rect 6528 873 6556 883
tri 6556 873 6580 897 sw
rect 6528 841 6570 873
tri 6587 865 6588 866 sw
rect 6587 841 6588 865
tri 6590 864 6627 901 ne
rect 6627 873 6632 901
tri 6632 873 6658 899 sw
rect 6742 883 6751 917
rect 6742 873 6770 883
rect 6627 864 6711 873
tri 6627 845 6646 864 ne
rect 6646 845 6711 864
rect 6528 819 6588 841
rect 6710 841 6711 845
rect 6728 841 6770 873
rect 6710 819 6770 841
rect 6616 803 6633 817
rect 6665 803 6682 817
tri 6453 767 6475 789 se
rect 6475 782 6490 803
tri 6475 767 6490 782 nw
rect 6809 782 6824 958
tri 6824 951 6837 964 nw
rect 6910 883 6925 1111
tri 6447 761 6453 767 se
rect 6453 761 6462 767
rect 6447 745 6462 761
tri 6462 754 6475 767 nw
rect 6616 759 6633 773
rect 6665 759 6682 773
tri 6809 767 6824 782 ne
tri 6824 767 6846 789 sw
rect 6447 709 6462 717
rect 6528 745 6588 759
rect 6543 735 6588 745
rect 6543 717 6571 735
tri 6447 694 6462 709 ne
tri 6462 694 6484 716 sw
rect 6528 707 6571 717
rect 6586 731 6588 735
rect 6710 745 6770 759
tri 6824 754 6837 767 ne
rect 6837 761 6846 767
tri 6846 761 6852 767 sw
rect 6710 735 6755 745
rect 6586 707 6660 731
rect 6528 703 6660 707
tri 6660 703 6688 731 sw
rect 6710 721 6712 735
tri 6710 719 6712 721 ne
rect 6724 717 6755 735
rect 6724 707 6770 717
rect 6837 746 6852 761
tri 6462 682 6474 694 ne
rect 6474 689 6484 694
tri 6484 689 6489 694 sw
rect 6373 343 6388 571
rect 6474 581 6489 689
rect 6528 647 6556 703
tri 6648 685 6666 703 ne
rect 6666 683 6688 703
tri 6688 683 6708 703 sw
tri 6724 689 6742 707 ne
rect 6547 613 6556 647
rect 6590 674 6632 675
rect 6590 640 6595 674
rect 6625 640 6632 674
rect 6590 631 6632 640
rect 6666 674 6708 683
rect 6666 640 6673 674
rect 6703 640 6708 674
rect 6666 635 6708 640
rect 6742 647 6770 707
tri 6815 694 6837 716 se
rect 6837 709 6852 717
tri 6837 694 6852 709 nw
tri 6809 688 6815 694 se
rect 6815 688 6824 694
rect 6528 603 6556 613
tri 6556 603 6580 627 sw
rect 6474 533 6490 581
rect 6528 571 6570 603
tri 6587 595 6588 596 sw
rect 6587 571 6588 595
tri 6590 594 6627 631 ne
rect 6627 603 6632 631
tri 6632 603 6658 629 sw
rect 6742 613 6751 647
rect 6742 603 6770 613
rect 6627 594 6711 603
tri 6627 575 6646 594 ne
rect 6646 575 6711 594
rect 6528 549 6588 571
rect 6710 571 6711 575
rect 6728 571 6770 603
rect 6710 549 6770 571
rect 6616 533 6633 547
rect 6665 533 6682 547
tri 6453 497 6475 519 se
rect 6475 512 6490 533
tri 6475 497 6490 512 nw
rect 6809 512 6824 688
tri 6824 681 6837 694 nw
rect 6910 613 6925 841
tri 6447 491 6453 497 se
rect 6453 491 6462 497
rect 6447 475 6462 491
tri 6462 484 6475 497 nw
rect 6616 489 6633 503
rect 6665 489 6682 503
tri 6809 497 6824 512 ne
tri 6824 497 6846 519 sw
rect 6447 439 6462 447
rect 6528 475 6588 489
rect 6543 465 6588 475
rect 6543 447 6571 465
tri 6447 424 6462 439 ne
tri 6462 424 6484 446 sw
rect 6528 437 6571 447
rect 6586 461 6588 465
rect 6710 475 6770 489
tri 6824 484 6837 497 ne
rect 6837 491 6846 497
tri 6846 491 6852 497 sw
rect 6710 465 6755 475
rect 6586 437 6660 461
rect 6528 433 6660 437
tri 6660 433 6688 461 sw
rect 6710 451 6712 465
tri 6710 449 6712 451 ne
rect 6724 447 6755 465
rect 6724 437 6770 447
rect 6837 476 6852 491
tri 6462 412 6474 424 ne
rect 6474 419 6484 424
tri 6484 419 6489 424 sw
rect 6373 73 6388 301
rect 6474 263 6489 419
rect 6528 377 6556 433
tri 6648 415 6666 433 ne
rect 6666 413 6688 433
tri 6688 413 6708 433 sw
tri 6724 419 6742 437 ne
rect 6547 343 6556 377
rect 6590 404 6632 405
rect 6590 370 6595 404
rect 6625 370 6632 404
rect 6590 361 6632 370
rect 6666 404 6708 413
rect 6666 370 6673 404
rect 6703 370 6708 404
rect 6666 365 6708 370
rect 6742 377 6770 437
tri 6815 424 6837 446 se
rect 6837 439 6852 447
tri 6837 424 6852 439 nw
tri 6809 418 6815 424 se
rect 6815 418 6824 424
rect 6528 333 6556 343
tri 6556 333 6580 357 sw
rect 6528 301 6570 333
tri 6587 325 6588 326 sw
rect 6587 301 6588 325
tri 6590 324 6627 361 ne
rect 6627 333 6632 361
tri 6632 333 6658 359 sw
rect 6742 343 6751 377
rect 6742 333 6770 343
rect 6627 324 6711 333
tri 6627 305 6646 324 ne
rect 6646 305 6711 324
rect 6528 279 6588 301
rect 6710 301 6711 305
rect 6728 301 6770 333
rect 6710 279 6770 301
rect 6616 263 6633 277
rect 6665 263 6682 277
tri 6453 227 6475 249 se
rect 6475 242 6490 263
tri 6475 227 6490 242 nw
rect 6809 242 6824 418
tri 6824 411 6837 424 nw
rect 6910 343 6925 571
tri 6447 221 6453 227 se
rect 6453 221 6462 227
rect 6447 205 6462 221
tri 6462 214 6475 227 nw
rect 6616 219 6633 233
rect 6665 219 6682 233
tri 6809 227 6824 242 ne
tri 6824 227 6846 249 sw
rect 6447 169 6462 177
rect 6528 205 6588 219
rect 6543 195 6588 205
rect 6543 177 6571 195
tri 6447 154 6462 169 ne
tri 6462 154 6484 176 sw
rect 6528 167 6571 177
rect 6586 191 6588 195
rect 6710 205 6770 219
tri 6824 214 6837 227 ne
rect 6837 221 6846 227
tri 6846 221 6852 227 sw
rect 6710 195 6755 205
rect 6586 167 6660 191
rect 6528 163 6660 167
tri 6660 163 6688 191 sw
rect 6710 181 6712 195
tri 6710 179 6712 181 ne
rect 6724 177 6755 195
rect 6724 167 6770 177
rect 6837 206 6852 221
tri 6462 142 6474 154 ne
rect 6474 149 6484 154
tri 6484 149 6489 154 sw
rect 6373 -55 6388 31
rect 6474 -55 6489 149
rect 6528 107 6556 163
tri 6648 145 6666 163 ne
rect 6666 143 6688 163
tri 6688 143 6708 163 sw
tri 6724 149 6742 167 ne
rect 6547 73 6556 107
rect 6590 134 6632 135
rect 6590 100 6595 134
rect 6625 100 6632 134
rect 6590 91 6632 100
rect 6666 134 6708 143
rect 6666 100 6673 134
rect 6703 100 6708 134
rect 6666 95 6708 100
rect 6742 107 6770 167
tri 6815 154 6837 176 se
rect 6837 169 6852 177
tri 6837 154 6852 169 nw
tri 6809 148 6815 154 se
rect 6815 148 6824 154
rect 6528 63 6556 73
tri 6556 63 6580 87 sw
rect 6528 31 6570 63
tri 6587 55 6588 56 sw
rect 6587 31 6588 55
tri 6590 54 6627 91 ne
rect 6627 63 6632 91
tri 6632 63 6658 89 sw
rect 6742 73 6751 107
rect 6742 63 6770 73
rect 6627 54 6711 63
tri 6627 35 6646 54 ne
rect 6646 35 6711 54
rect 6528 9 6588 31
rect 6710 31 6711 35
rect 6728 31 6770 63
rect 6710 9 6770 31
rect 6616 -7 6633 7
rect 6665 -7 6682 7
rect 6809 -55 6824 148
tri 6824 141 6837 154 nw
rect 6910 73 6925 301
rect 6910 -55 6925 31
<< viali >>
rect 253 4269 285 4283
rect 36 4145 66 4179
rect 253 4043 285 4057
rect 472 4145 502 4179
rect 253 3999 285 4013
rect 36 3875 66 3909
rect 253 3773 285 3787
rect 472 3876 502 3909
rect 253 3729 285 3743
rect 36 3605 66 3639
rect 253 3503 285 3517
rect 472 3606 502 3639
rect 253 3459 285 3473
rect 36 3335 66 3369
rect 253 3233 285 3247
rect 472 3336 502 3369
rect 253 3189 285 3203
rect 36 3065 66 3099
rect 253 2963 285 2977
rect 472 3066 502 3099
rect 253 2919 285 2933
rect 36 2795 66 2829
rect 253 2693 285 2707
rect 472 2796 502 2829
rect 253 2649 285 2663
rect 36 2525 66 2559
rect 253 2423 285 2437
rect 472 2526 502 2559
rect 253 2379 285 2393
rect 36 2255 66 2289
rect 253 2153 285 2167
rect 472 2256 502 2289
rect 253 2109 285 2123
rect 36 1985 66 2019
rect 253 1883 285 1897
rect 472 1986 502 2019
rect 253 1839 285 1853
rect 36 1715 66 1749
rect 253 1613 285 1627
rect 472 1716 502 1749
rect 253 1569 285 1583
rect 36 1445 66 1479
rect 253 1343 285 1357
rect 472 1446 502 1479
rect 253 1299 285 1313
rect 36 1175 66 1209
rect 253 1073 285 1087
rect 472 1176 502 1209
rect 253 1029 285 1043
rect 36 905 66 939
rect 253 803 285 817
rect 472 906 502 939
rect 253 759 285 773
rect 36 635 66 669
rect 253 533 285 547
rect 472 636 502 669
rect 253 489 285 503
rect 36 365 66 399
rect 253 263 285 277
rect 472 366 502 399
rect 253 219 285 233
rect 36 95 66 129
rect 253 -7 285 7
rect 472 96 502 129
rect 833 4269 865 4283
rect 616 4145 646 4179
rect 833 4043 865 4057
rect 1052 4145 1082 4179
rect 833 3999 865 4013
rect 616 3875 646 3909
rect 833 3773 865 3787
rect 1052 3875 1082 3909
rect 833 3729 865 3743
rect 616 3605 646 3639
rect 833 3503 865 3517
rect 1052 3605 1082 3639
rect 833 3459 865 3473
rect 616 3335 646 3369
rect 833 3233 865 3247
rect 1052 3335 1082 3369
rect 833 3189 865 3203
rect 616 3065 646 3099
rect 833 2963 865 2977
rect 1052 3065 1082 3099
rect 833 2919 865 2933
rect 616 2795 646 2829
rect 833 2693 865 2707
rect 1052 2795 1082 2829
rect 833 2649 865 2663
rect 616 2525 646 2559
rect 833 2423 865 2437
rect 1052 2525 1082 2559
rect 833 2379 865 2393
rect 616 2255 646 2289
rect 833 2153 865 2167
rect 1052 2255 1082 2289
rect 833 2109 865 2123
rect 616 1985 646 2019
rect 833 1883 865 1897
rect 1052 1985 1082 2019
rect 833 1839 865 1853
rect 616 1715 646 1749
rect 833 1613 865 1627
rect 1052 1715 1082 1749
rect 833 1569 865 1583
rect 616 1445 646 1479
rect 833 1343 865 1357
rect 1052 1445 1082 1479
rect 833 1299 865 1313
rect 616 1175 646 1209
rect 833 1073 865 1087
rect 1052 1175 1082 1209
rect 833 1029 865 1043
rect 616 905 646 939
rect 833 803 865 817
rect 1052 905 1082 939
rect 833 759 865 773
rect 616 635 646 669
rect 833 533 865 547
rect 1052 635 1082 669
rect 833 489 865 503
rect 616 365 646 399
rect 833 263 865 277
rect 1052 365 1082 399
rect 833 219 865 233
rect 616 95 646 129
rect 833 -7 865 7
rect 1052 95 1082 129
rect 1413 4269 1445 4283
rect 1196 4145 1226 4179
rect 1413 4043 1445 4057
rect 1632 4146 1662 4179
rect 1413 3999 1445 4013
rect 1196 3875 1226 3909
rect 1413 3773 1445 3787
rect 1632 3876 1662 3909
rect 1413 3729 1445 3743
rect 1196 3605 1226 3639
rect 1413 3503 1445 3517
rect 1632 3606 1662 3639
rect 1413 3459 1445 3473
rect 1196 3335 1226 3369
rect 1413 3233 1445 3247
rect 1632 3336 1662 3369
rect 1413 3189 1445 3203
rect 1196 3065 1226 3099
rect 1413 2963 1445 2977
rect 1632 3066 1662 3099
rect 1413 2919 1445 2933
rect 1196 2795 1226 2829
rect 1413 2693 1445 2707
rect 1632 2796 1662 2829
rect 1413 2649 1445 2663
rect 1196 2525 1226 2559
rect 1413 2423 1445 2437
rect 1632 2526 1662 2559
rect 1413 2379 1445 2393
rect 1196 2255 1226 2289
rect 1413 2153 1445 2167
rect 1632 2256 1662 2289
rect 1413 2109 1445 2123
rect 1196 1985 1226 2019
rect 1413 1883 1445 1897
rect 1632 1986 1662 2019
rect 1413 1839 1445 1853
rect 1196 1715 1226 1749
rect 1413 1613 1445 1627
rect 1632 1716 1662 1749
rect 1413 1569 1445 1583
rect 1196 1445 1226 1479
rect 1413 1343 1445 1357
rect 1632 1446 1662 1479
rect 1413 1299 1445 1313
rect 1196 1175 1226 1209
rect 1413 1073 1445 1087
rect 1632 1176 1662 1209
rect 1413 1029 1445 1043
rect 1196 905 1226 939
rect 1413 803 1445 817
rect 1632 906 1662 939
rect 1413 759 1445 773
rect 1196 635 1226 669
rect 1413 533 1445 547
rect 1632 636 1662 669
rect 1413 489 1445 503
rect 1196 365 1226 399
rect 1413 263 1445 277
rect 1632 366 1662 399
rect 1413 219 1445 233
rect 1196 95 1226 129
rect 1413 -7 1445 7
rect 1632 96 1662 129
rect 1993 4269 2025 4283
rect 1776 4145 1806 4179
rect 1993 4043 2025 4057
rect 2212 4145 2242 4179
rect 1993 3999 2025 4013
rect 1776 3875 1806 3909
rect 1993 3773 2025 3787
rect 2212 3875 2242 3909
rect 1993 3729 2025 3743
rect 1776 3605 1806 3639
rect 1993 3503 2025 3517
rect 2212 3605 2242 3639
rect 1993 3459 2025 3473
rect 1776 3335 1806 3369
rect 1993 3233 2025 3247
rect 2212 3335 2242 3369
rect 1993 3189 2025 3203
rect 1776 3065 1806 3099
rect 1993 2963 2025 2977
rect 2212 3065 2242 3099
rect 1993 2919 2025 2933
rect 1776 2795 1806 2829
rect 1993 2693 2025 2707
rect 2212 2795 2242 2829
rect 1993 2649 2025 2663
rect 1776 2525 1806 2559
rect 1993 2423 2025 2437
rect 2212 2525 2242 2559
rect 1993 2379 2025 2393
rect 1776 2255 1806 2289
rect 1993 2153 2025 2167
rect 2212 2255 2242 2289
rect 1993 2109 2025 2123
rect 1776 1985 1806 2019
rect 1993 1883 2025 1897
rect 2212 1985 2242 2019
rect 1993 1839 2025 1853
rect 1776 1715 1806 1749
rect 1993 1613 2025 1627
rect 2212 1715 2242 1749
rect 1993 1569 2025 1583
rect 1776 1445 1806 1479
rect 1993 1343 2025 1357
rect 2212 1445 2242 1479
rect 1993 1299 2025 1313
rect 1776 1175 1806 1209
rect 1993 1073 2025 1087
rect 2212 1175 2242 1209
rect 1993 1029 2025 1043
rect 1776 905 1806 939
rect 1993 803 2025 817
rect 2212 905 2242 939
rect 1993 759 2025 773
rect 1776 635 1806 669
rect 1993 533 2025 547
rect 2212 635 2242 669
rect 1993 489 2025 503
rect 1776 365 1806 399
rect 1993 263 2025 277
rect 2212 365 2242 399
rect 1993 219 2025 233
rect 1776 95 1806 129
rect 1993 -7 2025 7
rect 2212 95 2242 129
rect 2573 4269 2605 4283
rect 2356 4145 2386 4179
rect 2573 4043 2605 4057
rect 2792 4146 2822 4179
rect 2573 3999 2605 4013
rect 2356 3875 2386 3909
rect 2573 3773 2605 3787
rect 2792 3876 2822 3909
rect 2573 3729 2605 3743
rect 2356 3605 2386 3639
rect 2573 3503 2605 3517
rect 2792 3606 2822 3639
rect 2573 3459 2605 3473
rect 2356 3335 2386 3369
rect 2573 3233 2605 3247
rect 2792 3336 2822 3369
rect 2573 3189 2605 3203
rect 2356 3065 2386 3099
rect 2573 2963 2605 2977
rect 2792 3066 2822 3099
rect 2573 2919 2605 2933
rect 2356 2795 2386 2829
rect 2573 2693 2605 2707
rect 2792 2796 2822 2829
rect 2573 2649 2605 2663
rect 2356 2525 2386 2559
rect 2573 2423 2605 2437
rect 2792 2526 2822 2559
rect 2573 2379 2605 2393
rect 2356 2255 2386 2289
rect 2573 2153 2605 2167
rect 2792 2256 2822 2289
rect 2573 2109 2605 2123
rect 2356 1985 2386 2019
rect 2573 1883 2605 1897
rect 2792 1986 2822 2019
rect 2573 1839 2605 1853
rect 2356 1715 2386 1749
rect 2573 1613 2605 1627
rect 2792 1716 2822 1749
rect 2573 1569 2605 1583
rect 2356 1445 2386 1479
rect 2573 1343 2605 1357
rect 2792 1446 2822 1479
rect 2573 1299 2605 1313
rect 2356 1175 2386 1209
rect 2573 1073 2605 1087
rect 2792 1176 2822 1209
rect 2573 1029 2605 1043
rect 2356 905 2386 939
rect 2573 803 2605 817
rect 2792 906 2822 939
rect 2573 759 2605 773
rect 2356 635 2386 669
rect 2573 533 2605 547
rect 2792 636 2822 669
rect 2573 489 2605 503
rect 2356 365 2386 399
rect 2573 263 2605 277
rect 2792 366 2822 399
rect 2573 219 2605 233
rect 2356 95 2386 129
rect 2573 -7 2605 7
rect 2792 96 2822 129
rect 3153 4269 3185 4283
rect 2936 4145 2966 4179
rect 3153 4043 3185 4057
rect 3372 4145 3402 4179
rect 3153 3999 3185 4013
rect 2936 3875 2966 3909
rect 3153 3773 3185 3787
rect 3372 3875 3402 3909
rect 3153 3729 3185 3743
rect 2936 3605 2966 3639
rect 3153 3503 3185 3517
rect 3372 3605 3402 3639
rect 3153 3459 3185 3473
rect 2936 3335 2966 3369
rect 3153 3233 3185 3247
rect 3372 3335 3402 3369
rect 3153 3189 3185 3203
rect 2936 3065 2966 3099
rect 3153 2963 3185 2977
rect 3372 3065 3402 3099
rect 3153 2919 3185 2933
rect 2936 2795 2966 2829
rect 3153 2693 3185 2707
rect 3372 2795 3402 2829
rect 3153 2649 3185 2663
rect 2936 2525 2966 2559
rect 3153 2423 3185 2437
rect 3372 2525 3402 2559
rect 3153 2379 3185 2393
rect 2936 2255 2966 2289
rect 3153 2153 3185 2167
rect 3372 2255 3402 2289
rect 3153 2109 3185 2123
rect 2936 1985 2966 2019
rect 3153 1883 3185 1897
rect 3372 1985 3402 2019
rect 3153 1839 3185 1853
rect 2936 1715 2966 1749
rect 3153 1613 3185 1627
rect 3372 1715 3402 1749
rect 3153 1569 3185 1583
rect 2936 1445 2966 1479
rect 3153 1343 3185 1357
rect 3372 1445 3402 1479
rect 3153 1299 3185 1313
rect 2936 1175 2966 1209
rect 3153 1073 3185 1087
rect 3372 1175 3402 1209
rect 3153 1029 3185 1043
rect 2936 905 2966 939
rect 3153 803 3185 817
rect 3372 905 3402 939
rect 3153 759 3185 773
rect 2936 635 2966 669
rect 3153 533 3185 547
rect 3372 635 3402 669
rect 3153 489 3185 503
rect 2936 365 2966 399
rect 3153 263 3185 277
rect 3372 365 3402 399
rect 3153 219 3185 233
rect 2936 95 2966 129
rect 3153 -7 3185 7
rect 3372 95 3402 129
rect 3733 4269 3765 4283
rect 3516 4145 3546 4179
rect 3733 4043 3765 4057
rect 3952 4146 3982 4179
rect 3733 3999 3765 4013
rect 3516 3875 3546 3909
rect 3733 3773 3765 3787
rect 3952 3876 3982 3909
rect 3733 3729 3765 3743
rect 3516 3605 3546 3639
rect 3733 3503 3765 3517
rect 3952 3606 3982 3639
rect 3733 3459 3765 3473
rect 3516 3335 3546 3369
rect 3733 3233 3765 3247
rect 3952 3336 3982 3369
rect 3733 3189 3765 3203
rect 3516 3065 3546 3099
rect 3733 2963 3765 2977
rect 3952 3066 3982 3099
rect 3733 2919 3765 2933
rect 3516 2795 3546 2829
rect 3733 2693 3765 2707
rect 3952 2796 3982 2829
rect 3733 2649 3765 2663
rect 3516 2525 3546 2559
rect 3733 2423 3765 2437
rect 3952 2526 3982 2559
rect 3733 2379 3765 2393
rect 3516 2255 3546 2289
rect 3733 2153 3765 2167
rect 3952 2256 3982 2289
rect 3733 2109 3765 2123
rect 3516 1985 3546 2019
rect 3733 1883 3765 1897
rect 3952 1986 3982 2019
rect 3733 1839 3765 1853
rect 3516 1715 3546 1749
rect 3733 1613 3765 1627
rect 3952 1716 3982 1749
rect 3733 1569 3765 1583
rect 3516 1445 3546 1479
rect 3733 1343 3765 1357
rect 3952 1446 3982 1479
rect 3733 1299 3765 1313
rect 3516 1175 3546 1209
rect 3733 1073 3765 1087
rect 3952 1176 3982 1209
rect 3733 1029 3765 1043
rect 3516 905 3546 939
rect 3733 803 3765 817
rect 3952 906 3982 939
rect 3733 759 3765 773
rect 3516 635 3546 669
rect 3733 533 3765 547
rect 3952 636 3982 669
rect 3733 489 3765 503
rect 3516 365 3546 399
rect 3733 263 3765 277
rect 3952 366 3982 399
rect 3733 219 3765 233
rect 3516 95 3546 129
rect 3733 -7 3765 7
rect 3952 96 3982 129
rect 4313 4269 4345 4283
rect 4096 4145 4126 4179
rect 4313 4043 4345 4057
rect 4532 4145 4562 4179
rect 4313 3999 4345 4013
rect 4096 3875 4126 3909
rect 4313 3773 4345 3787
rect 4532 3875 4562 3909
rect 4313 3729 4345 3743
rect 4096 3605 4126 3639
rect 4313 3503 4345 3517
rect 4532 3605 4562 3639
rect 4313 3459 4345 3473
rect 4096 3335 4126 3369
rect 4313 3233 4345 3247
rect 4532 3335 4562 3369
rect 4313 3189 4345 3203
rect 4096 3065 4126 3099
rect 4313 2963 4345 2977
rect 4532 3065 4562 3099
rect 4313 2919 4345 2933
rect 4096 2795 4126 2829
rect 4313 2693 4345 2707
rect 4532 2795 4562 2829
rect 4313 2649 4345 2663
rect 4096 2525 4126 2559
rect 4313 2423 4345 2437
rect 4532 2525 4562 2559
rect 4313 2379 4345 2393
rect 4096 2255 4126 2289
rect 4313 2153 4345 2167
rect 4532 2255 4562 2289
rect 4313 2109 4345 2123
rect 4096 1985 4126 2019
rect 4313 1883 4345 1897
rect 4532 1985 4562 2019
rect 4313 1839 4345 1853
rect 4096 1715 4126 1749
rect 4313 1613 4345 1627
rect 4532 1715 4562 1749
rect 4313 1569 4345 1583
rect 4096 1445 4126 1479
rect 4313 1343 4345 1357
rect 4532 1445 4562 1479
rect 4313 1299 4345 1313
rect 4096 1175 4126 1209
rect 4313 1073 4345 1087
rect 4532 1175 4562 1209
rect 4313 1029 4345 1043
rect 4096 905 4126 939
rect 4313 803 4345 817
rect 4532 905 4562 939
rect 4313 759 4345 773
rect 4096 635 4126 669
rect 4313 533 4345 547
rect 4532 635 4562 669
rect 4313 489 4345 503
rect 4096 365 4126 399
rect 4313 263 4345 277
rect 4532 365 4562 399
rect 4313 219 4345 233
rect 4096 95 4126 129
rect 4313 -7 4345 7
rect 4532 95 4562 129
rect 4893 4269 4925 4283
rect 4676 4145 4706 4179
rect 4893 4043 4925 4057
rect 5112 4146 5142 4179
rect 4893 3999 4925 4013
rect 4676 3875 4706 3909
rect 4893 3773 4925 3787
rect 5112 3876 5142 3909
rect 4893 3729 4925 3743
rect 4676 3605 4706 3639
rect 4893 3503 4925 3517
rect 5112 3606 5142 3639
rect 4893 3459 4925 3473
rect 4676 3335 4706 3369
rect 4893 3233 4925 3247
rect 5112 3336 5142 3369
rect 4893 3189 4925 3203
rect 4676 3065 4706 3099
rect 4893 2963 4925 2977
rect 5112 3066 5142 3099
rect 4893 2919 4925 2933
rect 4676 2795 4706 2829
rect 4893 2693 4925 2707
rect 5112 2796 5142 2829
rect 4893 2649 4925 2663
rect 4676 2525 4706 2559
rect 4893 2423 4925 2437
rect 5112 2526 5142 2559
rect 4893 2379 4925 2393
rect 4676 2255 4706 2289
rect 4893 2153 4925 2167
rect 5112 2256 5142 2289
rect 4893 2109 4925 2123
rect 4676 1985 4706 2019
rect 4893 1883 4925 1897
rect 5112 1986 5142 2019
rect 4893 1839 4925 1853
rect 4676 1715 4706 1749
rect 4893 1613 4925 1627
rect 5112 1716 5142 1749
rect 4893 1569 4925 1583
rect 4676 1445 4706 1479
rect 4893 1343 4925 1357
rect 5112 1446 5142 1479
rect 4893 1299 4925 1313
rect 4676 1175 4706 1209
rect 4893 1073 4925 1087
rect 5112 1176 5142 1209
rect 4893 1029 4925 1043
rect 4676 905 4706 939
rect 4893 803 4925 817
rect 5112 906 5142 939
rect 4893 759 4925 773
rect 4676 635 4706 669
rect 4893 533 4925 547
rect 5112 636 5142 669
rect 4893 489 4925 503
rect 4676 365 4706 399
rect 4893 263 4925 277
rect 5112 366 5142 399
rect 4893 219 4925 233
rect 4676 95 4706 129
rect 4893 -7 4925 7
rect 5112 96 5142 129
rect 5473 4269 5505 4283
rect 5256 4145 5286 4179
rect 5473 4043 5505 4057
rect 5692 4145 5722 4179
rect 5473 3999 5505 4013
rect 5256 3875 5286 3909
rect 5473 3773 5505 3787
rect 5692 3875 5722 3909
rect 5473 3729 5505 3743
rect 5256 3605 5286 3639
rect 5473 3503 5505 3517
rect 5692 3605 5722 3639
rect 5473 3459 5505 3473
rect 5256 3335 5286 3369
rect 5473 3233 5505 3247
rect 5692 3335 5722 3369
rect 5473 3189 5505 3203
rect 5256 3065 5286 3099
rect 5473 2963 5505 2977
rect 5692 3065 5722 3099
rect 5473 2919 5505 2933
rect 5256 2795 5286 2829
rect 5473 2693 5505 2707
rect 5692 2795 5722 2829
rect 5473 2649 5505 2663
rect 5256 2525 5286 2559
rect 5473 2423 5505 2437
rect 5692 2525 5722 2559
rect 5473 2379 5505 2393
rect 5256 2255 5286 2289
rect 5473 2153 5505 2167
rect 5692 2255 5722 2289
rect 5473 2109 5505 2123
rect 5256 1985 5286 2019
rect 5473 1883 5505 1897
rect 5692 1985 5722 2019
rect 5473 1839 5505 1853
rect 5256 1715 5286 1749
rect 5473 1613 5505 1627
rect 5692 1715 5722 1749
rect 5473 1569 5505 1583
rect 5256 1445 5286 1479
rect 5473 1343 5505 1357
rect 5692 1445 5722 1479
rect 5473 1299 5505 1313
rect 5256 1175 5286 1209
rect 5473 1073 5505 1087
rect 5692 1175 5722 1209
rect 5473 1029 5505 1043
rect 5256 905 5286 939
rect 5473 803 5505 817
rect 5692 905 5722 939
rect 5473 759 5505 773
rect 5256 635 5286 669
rect 5473 533 5505 547
rect 5692 635 5722 669
rect 5473 489 5505 503
rect 5256 365 5286 399
rect 5473 263 5505 277
rect 5692 365 5722 399
rect 5473 219 5505 233
rect 5256 95 5286 129
rect 5473 -7 5505 7
rect 5692 95 5722 129
rect 6053 4269 6085 4283
rect 5836 4145 5866 4179
rect 6053 4043 6085 4057
rect 6272 4146 6302 4179
rect 6053 3999 6085 4013
rect 5836 3875 5866 3909
rect 6053 3773 6085 3787
rect 6272 3876 6302 3909
rect 6053 3729 6085 3743
rect 5836 3605 5866 3639
rect 6053 3503 6085 3517
rect 6272 3606 6302 3639
rect 6053 3459 6085 3473
rect 5836 3335 5866 3369
rect 6053 3233 6085 3247
rect 6272 3336 6302 3369
rect 6053 3189 6085 3203
rect 5836 3065 5866 3099
rect 6053 2963 6085 2977
rect 6272 3066 6302 3099
rect 6053 2919 6085 2933
rect 5836 2795 5866 2829
rect 6053 2693 6085 2707
rect 6272 2796 6302 2829
rect 6053 2649 6085 2663
rect 5836 2525 5866 2559
rect 6053 2423 6085 2437
rect 6272 2526 6302 2559
rect 6053 2379 6085 2393
rect 5836 2255 5866 2289
rect 6053 2153 6085 2167
rect 6272 2256 6302 2289
rect 6053 2109 6085 2123
rect 5836 1985 5866 2019
rect 6053 1883 6085 1897
rect 6272 1986 6302 2019
rect 6053 1839 6085 1853
rect 5836 1715 5866 1749
rect 6053 1613 6085 1627
rect 6272 1716 6302 1749
rect 6053 1569 6085 1583
rect 5836 1445 5866 1479
rect 6053 1343 6085 1357
rect 6272 1446 6302 1479
rect 6053 1299 6085 1313
rect 5836 1175 5866 1209
rect 6053 1073 6085 1087
rect 6272 1176 6302 1209
rect 6053 1029 6085 1043
rect 5836 905 5866 939
rect 6053 803 6085 817
rect 6272 906 6302 939
rect 6053 759 6085 773
rect 5836 635 5866 669
rect 6053 533 6085 547
rect 6272 636 6302 669
rect 6053 489 6085 503
rect 5836 365 5866 399
rect 6053 263 6085 277
rect 6272 366 6302 399
rect 6053 219 6085 233
rect 5836 95 5866 129
rect 6053 -7 6085 7
rect 6272 96 6302 129
rect 6633 4269 6665 4283
rect 6416 4145 6446 4179
rect 6633 4043 6665 4057
rect 6852 4145 6882 4179
rect 6633 3999 6665 4013
rect 6416 3875 6446 3909
rect 6633 3773 6665 3787
rect 6852 3875 6882 3909
rect 6633 3729 6665 3743
rect 6416 3605 6446 3639
rect 6633 3503 6665 3517
rect 6852 3605 6882 3639
rect 6633 3459 6665 3473
rect 6416 3335 6446 3369
rect 6633 3233 6665 3247
rect 6852 3335 6882 3369
rect 6633 3189 6665 3203
rect 6416 3065 6446 3099
rect 6633 2963 6665 2977
rect 6852 3065 6882 3099
rect 6633 2919 6665 2933
rect 6416 2795 6446 2829
rect 6633 2693 6665 2707
rect 6852 2795 6882 2829
rect 6633 2649 6665 2663
rect 6416 2525 6446 2559
rect 6633 2423 6665 2437
rect 6852 2525 6882 2559
rect 6633 2379 6665 2393
rect 6416 2255 6446 2289
rect 6633 2153 6665 2167
rect 6852 2255 6882 2289
rect 6633 2109 6665 2123
rect 6416 1985 6446 2019
rect 6633 1883 6665 1897
rect 6852 1985 6882 2019
rect 6633 1839 6665 1853
rect 6416 1715 6446 1749
rect 6633 1613 6665 1627
rect 6852 1715 6882 1749
rect 6633 1569 6665 1583
rect 6416 1445 6446 1479
rect 6633 1343 6665 1357
rect 6852 1445 6882 1479
rect 6633 1299 6665 1313
rect 6416 1175 6446 1209
rect 6633 1073 6665 1087
rect 6852 1175 6882 1209
rect 6633 1029 6665 1043
rect 6416 905 6446 939
rect 6633 803 6665 817
rect 6852 905 6882 939
rect 6633 759 6665 773
rect 6416 635 6446 669
rect 6633 533 6665 547
rect 6852 635 6882 669
rect 6633 489 6665 503
rect 6416 365 6446 399
rect 6633 263 6665 277
rect 6852 365 6882 399
rect 6633 219 6665 233
rect 6416 95 6446 129
rect 6633 -7 6665 7
rect 6852 95 6882 129
<< metal1 >>
rect -91 4269 253 4283
rect 285 4269 833 4283
rect 865 4269 1413 4283
rect 1445 4269 1993 4283
rect 2025 4269 2573 4283
rect 2605 4269 3153 4283
rect 3185 4269 3733 4283
rect 3765 4269 4313 4283
rect 4345 4269 4893 4283
rect 4925 4269 5473 4283
rect 5505 4269 6053 4283
rect 6085 4269 6633 4283
rect 6665 4269 6925 4283
tri 428 4205 462 4239 se
rect 462 4205 512 4239
tri 512 4205 546 4239 sw
tri 1008 4205 1042 4239 se
rect 1042 4205 1092 4239
tri 1092 4205 1126 4239 sw
tri 1588 4205 1622 4239 se
rect 1622 4205 1672 4239
tri 1672 4205 1706 4239 sw
tri 2168 4205 2202 4239 se
rect 2202 4205 2252 4239
tri 2252 4205 2286 4239 sw
tri 2748 4205 2782 4239 se
rect 2782 4205 2832 4239
tri 2832 4205 2866 4239 sw
tri 3328 4205 3362 4239 se
rect 3362 4205 3412 4239
tri 3412 4205 3446 4239 sw
tri 3908 4205 3942 4239 se
rect 3942 4205 3992 4239
tri 3992 4205 4026 4239 sw
tri 4488 4205 4522 4239 se
rect 4522 4205 4572 4239
tri 4572 4205 4606 4239 sw
tri 5068 4205 5102 4239 se
rect 5102 4205 5152 4239
tri 5152 4205 5186 4239 sw
tri 5648 4205 5682 4239 se
rect 5682 4205 5732 4239
tri 5732 4205 5766 4239 sw
tri 6228 4205 6262 4239 se
rect 6262 4205 6312 4239
tri 6312 4205 6346 4239 sw
tri 6808 4205 6842 4239 se
rect 6842 4205 6892 4239
tri 6892 4205 6926 4239 sw
tri 402 4179 428 4205 se
rect 428 4179 446 4205
tri 446 4179 472 4205 nw
tri 502 4179 528 4205 ne
rect 528 4179 546 4205
tri 546 4179 572 4205 sw
tri 982 4179 1008 4205 se
rect 1008 4179 1026 4205
tri 1026 4179 1052 4205 nw
tri 1082 4179 1108 4205 ne
rect 1108 4179 1126 4205
tri 1126 4179 1152 4205 sw
tri 1562 4179 1588 4205 se
rect 1588 4179 1606 4205
tri 1606 4179 1632 4205 nw
tri 1662 4179 1688 4205 ne
rect 1688 4179 1706 4205
tri 1706 4179 1732 4205 sw
tri 2142 4179 2168 4205 se
rect 2168 4179 2186 4205
tri 2186 4179 2212 4205 nw
tri 2242 4179 2268 4205 ne
rect 2268 4179 2286 4205
tri 2286 4179 2312 4205 sw
tri 2722 4179 2748 4205 se
rect 2748 4179 2766 4205
tri 2766 4179 2792 4205 nw
tri 2822 4179 2848 4205 ne
rect 2848 4179 2866 4205
tri 2866 4179 2892 4205 sw
tri 3302 4179 3328 4205 se
rect 3328 4179 3346 4205
tri 3346 4179 3372 4205 nw
tri 3402 4179 3428 4205 ne
rect 3428 4179 3446 4205
tri 3446 4179 3472 4205 sw
tri 3882 4179 3908 4205 se
rect 3908 4179 3926 4205
tri 3926 4179 3952 4205 nw
tri 3982 4179 4008 4205 ne
rect 4008 4179 4026 4205
tri 4026 4179 4052 4205 sw
tri 4462 4179 4488 4205 se
rect 4488 4179 4506 4205
tri 4506 4179 4532 4205 nw
tri 4562 4179 4588 4205 ne
rect 4588 4179 4606 4205
tri 4606 4179 4632 4205 sw
tri 5042 4179 5068 4205 se
rect 5068 4179 5086 4205
tri 5086 4179 5112 4205 nw
tri 5142 4179 5168 4205 ne
rect 5168 4179 5186 4205
tri 5186 4179 5212 4205 sw
tri 5622 4179 5648 4205 se
rect 5648 4179 5666 4205
tri 5666 4179 5692 4205 nw
tri 5722 4179 5748 4205 ne
rect 5748 4179 5766 4205
tri 5766 4179 5792 4205 sw
tri 6202 4179 6228 4205 se
rect 6228 4179 6246 4205
tri 6246 4179 6272 4205 nw
tri 6302 4179 6328 4205 ne
rect 6328 4179 6346 4205
tri 6346 4179 6372 4205 sw
tri 6782 4179 6808 4205 se
rect 6808 4179 6826 4205
tri 6826 4179 6852 4205 nw
tri 6882 4179 6908 4205 ne
rect 6908 4179 6926 4205
tri 6926 4179 6952 4205 sw
rect -91 4145 36 4179
rect 66 4145 412 4179
tri 412 4145 446 4179 nw
tri 528 4145 562 4179 ne
rect 562 4145 616 4179
rect 646 4145 992 4179
tri 992 4145 1026 4179 nw
rect 1105 4145 1196 4179
rect 1226 4145 1572 4179
tri 1572 4145 1606 4179 nw
tri 1688 4145 1722 4179 ne
rect 1722 4145 1776 4179
rect 1806 4145 2152 4179
tri 2152 4145 2186 4179 nw
rect 2265 4145 2356 4179
rect 2386 4145 2732 4179
tri 2732 4145 2766 4179 nw
tri 2848 4145 2882 4179 ne
rect 2882 4145 2936 4179
rect 2966 4145 3312 4179
tri 3312 4145 3346 4179 nw
rect 3425 4145 3516 4179
rect 3546 4145 3892 4179
tri 3892 4145 3926 4179 nw
tri 4008 4145 4042 4179 ne
rect 4042 4145 4096 4179
rect 4126 4145 4472 4179
tri 4472 4145 4506 4179 nw
rect 4585 4145 4676 4179
rect 4706 4145 5052 4179
tri 5052 4145 5086 4179 nw
tri 5168 4145 5202 4179 ne
rect 5202 4145 5256 4179
rect 5286 4145 5632 4179
tri 5632 4145 5666 4179 nw
rect 5745 4145 5836 4179
rect 5866 4145 6212 4179
tri 6212 4145 6246 4179 nw
tri 6328 4145 6362 4179 ne
rect 6362 4145 6416 4179
rect 6446 4145 6792 4179
tri 6792 4145 6826 4179 nw
tri 6908 4145 6942 4179 ne
rect 6942 4145 6952 4179
rect -91 4043 253 4057
rect 285 4043 833 4057
rect 865 4043 1413 4057
rect 1445 4043 1993 4057
rect 2025 4043 2573 4057
rect 2605 4043 3153 4057
rect 3185 4043 3733 4057
rect 3765 4043 4313 4057
rect 4345 4043 4893 4057
rect 4925 4043 5473 4057
rect 5505 4043 6053 4057
rect 6085 4043 6633 4057
rect 6665 4043 6925 4057
rect -91 3999 253 4013
rect 285 3999 833 4013
rect 865 3999 1413 4013
rect 1445 3999 1993 4013
rect 2025 3999 2573 4013
rect 2605 3999 3153 4013
rect 3185 3999 3733 4013
rect 3765 3999 4313 4013
rect 4345 3999 4893 4013
rect 4925 3999 5473 4013
rect 5505 3999 6053 4013
rect 6085 3999 6633 4013
rect 6665 3999 6925 4013
tri 428 3935 462 3969 se
rect 462 3935 512 3969
tri 512 3935 546 3969 sw
tri 1008 3935 1042 3969 se
rect 1042 3935 1092 3969
tri 1092 3935 1126 3969 sw
tri 1588 3935 1622 3969 se
rect 1622 3935 1672 3969
tri 1672 3935 1706 3969 sw
tri 2168 3935 2202 3969 se
rect 2202 3935 2252 3969
tri 2252 3935 2286 3969 sw
tri 2748 3935 2782 3969 se
rect 2782 3935 2832 3969
tri 2832 3935 2866 3969 sw
tri 3328 3935 3362 3969 se
rect 3362 3935 3412 3969
tri 3412 3935 3446 3969 sw
tri 3908 3935 3942 3969 se
rect 3942 3935 3992 3969
tri 3992 3935 4026 3969 sw
tri 4488 3935 4522 3969 se
rect 4522 3935 4572 3969
tri 4572 3935 4606 3969 sw
tri 5068 3935 5102 3969 se
rect 5102 3935 5152 3969
tri 5152 3935 5186 3969 sw
tri 5648 3935 5682 3969 se
rect 5682 3935 5732 3969
tri 5732 3935 5766 3969 sw
tri 6228 3935 6262 3969 se
rect 6262 3935 6312 3969
tri 6312 3935 6346 3969 sw
tri 6808 3935 6842 3969 se
rect 6842 3935 6892 3969
tri 6892 3935 6926 3969 sw
tri 402 3909 428 3935 se
rect 428 3909 446 3935
tri 446 3909 472 3935 nw
tri 502 3909 528 3935 ne
rect 528 3909 546 3935
tri 546 3909 572 3935 sw
tri 982 3909 1008 3935 se
rect 1008 3909 1026 3935
tri 1026 3909 1052 3935 nw
tri 1082 3909 1108 3935 ne
rect 1108 3909 1126 3935
tri 1126 3909 1152 3935 sw
tri 1562 3909 1588 3935 se
rect 1588 3909 1606 3935
tri 1606 3909 1632 3935 nw
tri 1662 3909 1688 3935 ne
rect 1688 3909 1706 3935
tri 1706 3909 1732 3935 sw
tri 2142 3909 2168 3935 se
rect 2168 3909 2186 3935
tri 2186 3909 2212 3935 nw
tri 2242 3909 2268 3935 ne
rect 2268 3909 2286 3935
tri 2286 3909 2312 3935 sw
tri 2722 3909 2748 3935 se
rect 2748 3909 2766 3935
tri 2766 3909 2792 3935 nw
tri 2822 3909 2848 3935 ne
rect 2848 3909 2866 3935
tri 2866 3909 2892 3935 sw
tri 3302 3909 3328 3935 se
rect 3328 3909 3346 3935
tri 3346 3909 3372 3935 nw
tri 3402 3909 3428 3935 ne
rect 3428 3909 3446 3935
tri 3446 3909 3472 3935 sw
tri 3882 3909 3908 3935 se
rect 3908 3909 3926 3935
tri 3926 3909 3952 3935 nw
tri 3982 3909 4008 3935 ne
rect 4008 3909 4026 3935
tri 4026 3909 4052 3935 sw
tri 4462 3909 4488 3935 se
rect 4488 3909 4506 3935
tri 4506 3909 4532 3935 nw
tri 4562 3909 4588 3935 ne
rect 4588 3909 4606 3935
tri 4606 3909 4632 3935 sw
tri 5042 3909 5068 3935 se
rect 5068 3909 5086 3935
tri 5086 3909 5112 3935 nw
tri 5142 3909 5168 3935 ne
rect 5168 3909 5186 3935
tri 5186 3909 5212 3935 sw
tri 5622 3909 5648 3935 se
rect 5648 3909 5666 3935
tri 5666 3909 5692 3935 nw
tri 5722 3909 5748 3935 ne
rect 5748 3909 5766 3935
tri 5766 3909 5792 3935 sw
tri 6202 3909 6228 3935 se
rect 6228 3909 6246 3935
tri 6246 3909 6272 3935 nw
tri 6302 3909 6328 3935 ne
rect 6328 3909 6346 3935
tri 6346 3909 6372 3935 sw
tri 6782 3909 6808 3935 se
rect 6808 3909 6826 3935
tri 6826 3909 6852 3935 nw
tri 6882 3909 6908 3935 ne
rect 6908 3909 6926 3935
tri 6926 3909 6952 3935 sw
rect -91 3875 36 3909
rect 66 3875 412 3909
tri 412 3875 446 3909 nw
tri 528 3875 562 3909 ne
rect 562 3875 616 3909
rect 646 3875 992 3909
tri 992 3875 1026 3909 nw
rect 1105 3875 1196 3909
rect 1226 3875 1572 3909
tri 1572 3875 1606 3909 nw
tri 1688 3875 1722 3909 ne
rect 1722 3875 1776 3909
rect 1806 3875 2152 3909
tri 2152 3875 2186 3909 nw
rect 2265 3875 2356 3909
rect 2386 3875 2732 3909
tri 2732 3875 2766 3909 nw
tri 2848 3875 2882 3909 ne
rect 2882 3875 2936 3909
rect 2966 3875 3312 3909
tri 3312 3875 3346 3909 nw
rect 3425 3875 3516 3909
rect 3546 3875 3892 3909
tri 3892 3875 3926 3909 nw
tri 4008 3875 4042 3909 ne
rect 4042 3875 4096 3909
rect 4126 3875 4472 3909
tri 4472 3875 4506 3909 nw
rect 4585 3875 4676 3909
rect 4706 3875 5052 3909
tri 5052 3875 5086 3909 nw
tri 5168 3875 5202 3909 ne
rect 5202 3875 5256 3909
rect 5286 3875 5632 3909
tri 5632 3875 5666 3909 nw
rect 5745 3875 5836 3909
rect 5866 3875 6212 3909
tri 6212 3875 6246 3909 nw
tri 6328 3875 6362 3909 ne
rect 6362 3875 6416 3909
rect 6446 3875 6792 3909
tri 6792 3875 6826 3909 nw
tri 6908 3875 6942 3909 ne
rect 6942 3875 6952 3909
rect -91 3773 253 3787
rect 285 3773 833 3787
rect 865 3773 1413 3787
rect 1445 3773 1993 3787
rect 2025 3773 2573 3787
rect 2605 3773 3153 3787
rect 3185 3773 3733 3787
rect 3765 3773 4313 3787
rect 4345 3773 4893 3787
rect 4925 3773 5473 3787
rect 5505 3773 6053 3787
rect 6085 3773 6633 3787
rect 6665 3773 6925 3787
rect -91 3729 253 3743
rect 285 3729 833 3743
rect 865 3729 1413 3743
rect 1445 3729 1993 3743
rect 2025 3729 2573 3743
rect 2605 3729 3153 3743
rect 3185 3729 3733 3743
rect 3765 3729 4313 3743
rect 4345 3729 4893 3743
rect 4925 3729 5473 3743
rect 5505 3729 6053 3743
rect 6085 3729 6633 3743
rect 6665 3729 6925 3743
tri 428 3665 462 3699 se
rect 462 3665 512 3699
tri 512 3665 546 3699 sw
tri 1008 3665 1042 3699 se
rect 1042 3665 1092 3699
tri 1092 3665 1126 3699 sw
tri 1588 3665 1622 3699 se
rect 1622 3665 1672 3699
tri 1672 3665 1706 3699 sw
tri 2168 3665 2202 3699 se
rect 2202 3665 2252 3699
tri 2252 3665 2286 3699 sw
tri 2748 3665 2782 3699 se
rect 2782 3665 2832 3699
tri 2832 3665 2866 3699 sw
tri 3328 3665 3362 3699 se
rect 3362 3665 3412 3699
tri 3412 3665 3446 3699 sw
tri 3908 3665 3942 3699 se
rect 3942 3665 3992 3699
tri 3992 3665 4026 3699 sw
tri 4488 3665 4522 3699 se
rect 4522 3665 4572 3699
tri 4572 3665 4606 3699 sw
tri 5068 3665 5102 3699 se
rect 5102 3665 5152 3699
tri 5152 3665 5186 3699 sw
tri 5648 3665 5682 3699 se
rect 5682 3665 5732 3699
tri 5732 3665 5766 3699 sw
tri 6228 3665 6262 3699 se
rect 6262 3665 6312 3699
tri 6312 3665 6346 3699 sw
tri 6808 3665 6842 3699 se
rect 6842 3665 6892 3699
tri 6892 3665 6926 3699 sw
tri 402 3639 428 3665 se
rect 428 3639 446 3665
tri 446 3639 472 3665 nw
tri 502 3639 528 3665 ne
rect 528 3639 546 3665
tri 546 3639 572 3665 sw
tri 982 3639 1008 3665 se
rect 1008 3639 1026 3665
tri 1026 3639 1052 3665 nw
tri 1082 3639 1108 3665 ne
rect 1108 3639 1126 3665
tri 1126 3639 1152 3665 sw
tri 1562 3639 1588 3665 se
rect 1588 3639 1606 3665
tri 1606 3639 1632 3665 nw
tri 1662 3639 1688 3665 ne
rect 1688 3639 1706 3665
tri 1706 3639 1732 3665 sw
tri 2142 3639 2168 3665 se
rect 2168 3639 2186 3665
tri 2186 3639 2212 3665 nw
tri 2242 3639 2268 3665 ne
rect 2268 3639 2286 3665
tri 2286 3639 2312 3665 sw
tri 2722 3639 2748 3665 se
rect 2748 3639 2766 3665
tri 2766 3639 2792 3665 nw
tri 2822 3639 2848 3665 ne
rect 2848 3639 2866 3665
tri 2866 3639 2892 3665 sw
tri 3302 3639 3328 3665 se
rect 3328 3639 3346 3665
tri 3346 3639 3372 3665 nw
tri 3402 3639 3428 3665 ne
rect 3428 3639 3446 3665
tri 3446 3639 3472 3665 sw
tri 3882 3639 3908 3665 se
rect 3908 3639 3926 3665
tri 3926 3639 3952 3665 nw
tri 3982 3639 4008 3665 ne
rect 4008 3639 4026 3665
tri 4026 3639 4052 3665 sw
tri 4462 3639 4488 3665 se
rect 4488 3639 4506 3665
tri 4506 3639 4532 3665 nw
tri 4562 3639 4588 3665 ne
rect 4588 3639 4606 3665
tri 4606 3639 4632 3665 sw
tri 5042 3639 5068 3665 se
rect 5068 3639 5086 3665
tri 5086 3639 5112 3665 nw
tri 5142 3639 5168 3665 ne
rect 5168 3639 5186 3665
tri 5186 3639 5212 3665 sw
tri 5622 3639 5648 3665 se
rect 5648 3639 5666 3665
tri 5666 3639 5692 3665 nw
tri 5722 3639 5748 3665 ne
rect 5748 3639 5766 3665
tri 5766 3639 5792 3665 sw
tri 6202 3639 6228 3665 se
rect 6228 3639 6246 3665
tri 6246 3639 6272 3665 nw
tri 6302 3639 6328 3665 ne
rect 6328 3639 6346 3665
tri 6346 3639 6372 3665 sw
tri 6782 3639 6808 3665 se
rect 6808 3639 6826 3665
tri 6826 3639 6852 3665 nw
tri 6882 3639 6908 3665 ne
rect 6908 3639 6926 3665
tri 6926 3639 6952 3665 sw
rect -91 3605 36 3639
rect 66 3605 412 3639
tri 412 3605 446 3639 nw
tri 528 3605 562 3639 ne
rect 562 3605 616 3639
rect 646 3605 992 3639
tri 992 3605 1026 3639 nw
rect 1105 3605 1196 3639
rect 1226 3605 1572 3639
tri 1572 3605 1606 3639 nw
tri 1688 3605 1722 3639 ne
rect 1722 3605 1776 3639
rect 1806 3605 2152 3639
tri 2152 3605 2186 3639 nw
rect 2265 3605 2356 3639
rect 2386 3605 2732 3639
tri 2732 3605 2766 3639 nw
tri 2848 3605 2882 3639 ne
rect 2882 3605 2936 3639
rect 2966 3605 3312 3639
tri 3312 3605 3346 3639 nw
rect 3425 3605 3516 3639
rect 3546 3605 3892 3639
tri 3892 3605 3926 3639 nw
tri 4008 3605 4042 3639 ne
rect 4042 3605 4096 3639
rect 4126 3605 4472 3639
tri 4472 3605 4506 3639 nw
rect 4585 3605 4676 3639
rect 4706 3605 5052 3639
tri 5052 3605 5086 3639 nw
tri 5168 3605 5202 3639 ne
rect 5202 3605 5256 3639
rect 5286 3605 5632 3639
tri 5632 3605 5666 3639 nw
rect 5745 3605 5836 3639
rect 5866 3605 6212 3639
tri 6212 3605 6246 3639 nw
tri 6328 3605 6362 3639 ne
rect 6362 3605 6416 3639
rect 6446 3605 6792 3639
tri 6792 3605 6826 3639 nw
tri 6908 3605 6942 3639 ne
rect 6942 3605 6952 3639
rect -91 3503 253 3517
rect 285 3503 833 3517
rect 865 3503 1413 3517
rect 1445 3503 1993 3517
rect 2025 3503 2573 3517
rect 2605 3503 3153 3517
rect 3185 3503 3733 3517
rect 3765 3503 4313 3517
rect 4345 3503 4893 3517
rect 4925 3503 5473 3517
rect 5505 3503 6053 3517
rect 6085 3503 6633 3517
rect 6665 3503 6925 3517
rect -91 3459 253 3473
rect 285 3459 833 3473
rect 865 3459 1413 3473
rect 1445 3459 1993 3473
rect 2025 3459 2573 3473
rect 2605 3459 3153 3473
rect 3185 3459 3733 3473
rect 3765 3459 4313 3473
rect 4345 3459 4893 3473
rect 4925 3459 5473 3473
rect 5505 3459 6053 3473
rect 6085 3459 6633 3473
rect 6665 3459 6925 3473
tri 428 3395 462 3429 se
rect 462 3395 512 3429
tri 512 3395 546 3429 sw
tri 1008 3395 1042 3429 se
rect 1042 3395 1092 3429
tri 1092 3395 1126 3429 sw
tri 1588 3395 1622 3429 se
rect 1622 3395 1672 3429
tri 1672 3395 1706 3429 sw
tri 2168 3395 2202 3429 se
rect 2202 3395 2252 3429
tri 2252 3395 2286 3429 sw
tri 2748 3395 2782 3429 se
rect 2782 3395 2832 3429
tri 2832 3395 2866 3429 sw
tri 3328 3395 3362 3429 se
rect 3362 3395 3412 3429
tri 3412 3395 3446 3429 sw
tri 3908 3395 3942 3429 se
rect 3942 3395 3992 3429
tri 3992 3395 4026 3429 sw
tri 4488 3395 4522 3429 se
rect 4522 3395 4572 3429
tri 4572 3395 4606 3429 sw
tri 5068 3395 5102 3429 se
rect 5102 3395 5152 3429
tri 5152 3395 5186 3429 sw
tri 5648 3395 5682 3429 se
rect 5682 3395 5732 3429
tri 5732 3395 5766 3429 sw
tri 6228 3395 6262 3429 se
rect 6262 3395 6312 3429
tri 6312 3395 6346 3429 sw
tri 6808 3395 6842 3429 se
rect 6842 3395 6892 3429
tri 6892 3395 6926 3429 sw
tri 402 3369 428 3395 se
rect 428 3369 446 3395
tri 446 3369 472 3395 nw
tri 502 3369 528 3395 ne
rect 528 3369 546 3395
tri 546 3369 572 3395 sw
tri 982 3369 1008 3395 se
rect 1008 3369 1026 3395
tri 1026 3369 1052 3395 nw
tri 1082 3369 1108 3395 ne
rect 1108 3369 1126 3395
tri 1126 3369 1152 3395 sw
tri 1562 3369 1588 3395 se
rect 1588 3369 1606 3395
tri 1606 3369 1632 3395 nw
tri 1662 3369 1688 3395 ne
rect 1688 3369 1706 3395
tri 1706 3369 1732 3395 sw
tri 2142 3369 2168 3395 se
rect 2168 3369 2186 3395
tri 2186 3369 2212 3395 nw
tri 2242 3369 2268 3395 ne
rect 2268 3369 2286 3395
tri 2286 3369 2312 3395 sw
tri 2722 3369 2748 3395 se
rect 2748 3369 2766 3395
tri 2766 3369 2792 3395 nw
tri 2822 3369 2848 3395 ne
rect 2848 3369 2866 3395
tri 2866 3369 2892 3395 sw
tri 3302 3369 3328 3395 se
rect 3328 3369 3346 3395
tri 3346 3369 3372 3395 nw
tri 3402 3369 3428 3395 ne
rect 3428 3369 3446 3395
tri 3446 3369 3472 3395 sw
tri 3882 3369 3908 3395 se
rect 3908 3369 3926 3395
tri 3926 3369 3952 3395 nw
tri 3982 3369 4008 3395 ne
rect 4008 3369 4026 3395
tri 4026 3369 4052 3395 sw
tri 4462 3369 4488 3395 se
rect 4488 3369 4506 3395
tri 4506 3369 4532 3395 nw
tri 4562 3369 4588 3395 ne
rect 4588 3369 4606 3395
tri 4606 3369 4632 3395 sw
tri 5042 3369 5068 3395 se
rect 5068 3369 5086 3395
tri 5086 3369 5112 3395 nw
tri 5142 3369 5168 3395 ne
rect 5168 3369 5186 3395
tri 5186 3369 5212 3395 sw
tri 5622 3369 5648 3395 se
rect 5648 3369 5666 3395
tri 5666 3369 5692 3395 nw
tri 5722 3369 5748 3395 ne
rect 5748 3369 5766 3395
tri 5766 3369 5792 3395 sw
tri 6202 3369 6228 3395 se
rect 6228 3369 6246 3395
tri 6246 3369 6272 3395 nw
tri 6302 3369 6328 3395 ne
rect 6328 3369 6346 3395
tri 6346 3369 6372 3395 sw
tri 6782 3369 6808 3395 se
rect 6808 3369 6826 3395
tri 6826 3369 6852 3395 nw
tri 6882 3369 6908 3395 ne
rect 6908 3369 6926 3395
tri 6926 3369 6952 3395 sw
rect -91 3335 36 3369
rect 66 3335 412 3369
tri 412 3335 446 3369 nw
tri 528 3335 562 3369 ne
rect 562 3335 616 3369
rect 646 3335 992 3369
tri 992 3335 1026 3369 nw
rect 1105 3335 1196 3369
rect 1226 3335 1572 3369
tri 1572 3335 1606 3369 nw
tri 1688 3335 1722 3369 ne
rect 1722 3335 1776 3369
rect 1806 3335 2152 3369
tri 2152 3335 2186 3369 nw
rect 2265 3335 2356 3369
rect 2386 3335 2732 3369
tri 2732 3335 2766 3369 nw
tri 2848 3335 2882 3369 ne
rect 2882 3335 2936 3369
rect 2966 3335 3312 3369
tri 3312 3335 3346 3369 nw
rect 3425 3335 3516 3369
rect 3546 3335 3892 3369
tri 3892 3335 3926 3369 nw
tri 4008 3335 4042 3369 ne
rect 4042 3335 4096 3369
rect 4126 3335 4472 3369
tri 4472 3335 4506 3369 nw
rect 4585 3335 4676 3369
rect 4706 3335 5052 3369
tri 5052 3335 5086 3369 nw
tri 5168 3335 5202 3369 ne
rect 5202 3335 5256 3369
rect 5286 3335 5632 3369
tri 5632 3335 5666 3369 nw
rect 5745 3335 5836 3369
rect 5866 3335 6212 3369
tri 6212 3335 6246 3369 nw
tri 6328 3335 6362 3369 ne
rect 6362 3335 6416 3369
rect 6446 3335 6792 3369
tri 6792 3335 6826 3369 nw
tri 6908 3335 6942 3369 ne
rect 6942 3335 6952 3369
rect -91 3233 253 3247
rect 285 3233 833 3247
rect 865 3233 1413 3247
rect 1445 3233 1993 3247
rect 2025 3233 2573 3247
rect 2605 3233 3153 3247
rect 3185 3233 3733 3247
rect 3765 3233 4313 3247
rect 4345 3233 4893 3247
rect 4925 3233 5473 3247
rect 5505 3233 6053 3247
rect 6085 3233 6633 3247
rect 6665 3233 6925 3247
rect -91 3189 253 3203
rect 285 3189 833 3203
rect 865 3189 1413 3203
rect 1445 3189 1993 3203
rect 2025 3189 2573 3203
rect 2605 3189 3153 3203
rect 3185 3189 3733 3203
rect 3765 3189 4313 3203
rect 4345 3189 4893 3203
rect 4925 3189 5473 3203
rect 5505 3189 6053 3203
rect 6085 3189 6633 3203
rect 6665 3189 6925 3203
tri 428 3125 462 3159 se
rect 462 3125 512 3159
tri 512 3125 546 3159 sw
tri 1008 3125 1042 3159 se
rect 1042 3125 1092 3159
tri 1092 3125 1126 3159 sw
tri 1588 3125 1622 3159 se
rect 1622 3125 1672 3159
tri 1672 3125 1706 3159 sw
tri 2168 3125 2202 3159 se
rect 2202 3125 2252 3159
tri 2252 3125 2286 3159 sw
tri 2748 3125 2782 3159 se
rect 2782 3125 2832 3159
tri 2832 3125 2866 3159 sw
tri 3328 3125 3362 3159 se
rect 3362 3125 3412 3159
tri 3412 3125 3446 3159 sw
tri 3908 3125 3942 3159 se
rect 3942 3125 3992 3159
tri 3992 3125 4026 3159 sw
tri 4488 3125 4522 3159 se
rect 4522 3125 4572 3159
tri 4572 3125 4606 3159 sw
tri 5068 3125 5102 3159 se
rect 5102 3125 5152 3159
tri 5152 3125 5186 3159 sw
tri 5648 3125 5682 3159 se
rect 5682 3125 5732 3159
tri 5732 3125 5766 3159 sw
tri 6228 3125 6262 3159 se
rect 6262 3125 6312 3159
tri 6312 3125 6346 3159 sw
tri 6808 3125 6842 3159 se
rect 6842 3125 6892 3159
tri 6892 3125 6926 3159 sw
tri 402 3099 428 3125 se
rect 428 3099 446 3125
tri 446 3099 472 3125 nw
tri 502 3099 528 3125 ne
rect 528 3099 546 3125
tri 546 3099 572 3125 sw
tri 982 3099 1008 3125 se
rect 1008 3099 1026 3125
tri 1026 3099 1052 3125 nw
tri 1082 3099 1108 3125 ne
rect 1108 3099 1126 3125
tri 1126 3099 1152 3125 sw
tri 1562 3099 1588 3125 se
rect 1588 3099 1606 3125
tri 1606 3099 1632 3125 nw
tri 1662 3099 1688 3125 ne
rect 1688 3099 1706 3125
tri 1706 3099 1732 3125 sw
tri 2142 3099 2168 3125 se
rect 2168 3099 2186 3125
tri 2186 3099 2212 3125 nw
tri 2242 3099 2268 3125 ne
rect 2268 3099 2286 3125
tri 2286 3099 2312 3125 sw
tri 2722 3099 2748 3125 se
rect 2748 3099 2766 3125
tri 2766 3099 2792 3125 nw
tri 2822 3099 2848 3125 ne
rect 2848 3099 2866 3125
tri 2866 3099 2892 3125 sw
tri 3302 3099 3328 3125 se
rect 3328 3099 3346 3125
tri 3346 3099 3372 3125 nw
tri 3402 3099 3428 3125 ne
rect 3428 3099 3446 3125
tri 3446 3099 3472 3125 sw
tri 3882 3099 3908 3125 se
rect 3908 3099 3926 3125
tri 3926 3099 3952 3125 nw
tri 3982 3099 4008 3125 ne
rect 4008 3099 4026 3125
tri 4026 3099 4052 3125 sw
tri 4462 3099 4488 3125 se
rect 4488 3099 4506 3125
tri 4506 3099 4532 3125 nw
tri 4562 3099 4588 3125 ne
rect 4588 3099 4606 3125
tri 4606 3099 4632 3125 sw
tri 5042 3099 5068 3125 se
rect 5068 3099 5086 3125
tri 5086 3099 5112 3125 nw
tri 5142 3099 5168 3125 ne
rect 5168 3099 5186 3125
tri 5186 3099 5212 3125 sw
tri 5622 3099 5648 3125 se
rect 5648 3099 5666 3125
tri 5666 3099 5692 3125 nw
tri 5722 3099 5748 3125 ne
rect 5748 3099 5766 3125
tri 5766 3099 5792 3125 sw
tri 6202 3099 6228 3125 se
rect 6228 3099 6246 3125
tri 6246 3099 6272 3125 nw
tri 6302 3099 6328 3125 ne
rect 6328 3099 6346 3125
tri 6346 3099 6372 3125 sw
tri 6782 3099 6808 3125 se
rect 6808 3099 6826 3125
tri 6826 3099 6852 3125 nw
tri 6882 3099 6908 3125 ne
rect 6908 3099 6926 3125
tri 6926 3099 6952 3125 sw
rect -91 3065 36 3099
rect 66 3065 412 3099
tri 412 3065 446 3099 nw
tri 528 3065 562 3099 ne
rect 562 3065 616 3099
rect 646 3065 992 3099
tri 992 3065 1026 3099 nw
rect 1105 3065 1196 3099
rect 1226 3065 1572 3099
tri 1572 3065 1606 3099 nw
tri 1688 3065 1722 3099 ne
rect 1722 3065 1776 3099
rect 1806 3065 2152 3099
tri 2152 3065 2186 3099 nw
rect 2265 3065 2356 3099
rect 2386 3065 2732 3099
tri 2732 3065 2766 3099 nw
tri 2848 3065 2882 3099 ne
rect 2882 3065 2936 3099
rect 2966 3065 3312 3099
tri 3312 3065 3346 3099 nw
rect 3425 3065 3516 3099
rect 3546 3065 3892 3099
tri 3892 3065 3926 3099 nw
tri 4008 3065 4042 3099 ne
rect 4042 3065 4096 3099
rect 4126 3065 4472 3099
tri 4472 3065 4506 3099 nw
rect 4585 3065 4676 3099
rect 4706 3065 5052 3099
tri 5052 3065 5086 3099 nw
tri 5168 3065 5202 3099 ne
rect 5202 3065 5256 3099
rect 5286 3065 5632 3099
tri 5632 3065 5666 3099 nw
rect 5745 3065 5836 3099
rect 5866 3065 6212 3099
tri 6212 3065 6246 3099 nw
tri 6328 3065 6362 3099 ne
rect 6362 3065 6416 3099
rect 6446 3065 6792 3099
tri 6792 3065 6826 3099 nw
tri 6908 3065 6942 3099 ne
rect 6942 3065 6952 3099
rect -91 2963 253 2977
rect 285 2963 833 2977
rect 865 2963 1413 2977
rect 1445 2963 1993 2977
rect 2025 2963 2573 2977
rect 2605 2963 3153 2977
rect 3185 2963 3733 2977
rect 3765 2963 4313 2977
rect 4345 2963 4893 2977
rect 4925 2963 5473 2977
rect 5505 2963 6053 2977
rect 6085 2963 6633 2977
rect 6665 2963 6925 2977
rect -91 2919 253 2933
rect 285 2919 833 2933
rect 865 2919 1413 2933
rect 1445 2919 1993 2933
rect 2025 2919 2573 2933
rect 2605 2919 3153 2933
rect 3185 2919 3733 2933
rect 3765 2919 4313 2933
rect 4345 2919 4893 2933
rect 4925 2919 5473 2933
rect 5505 2919 6053 2933
rect 6085 2919 6633 2933
rect 6665 2919 6925 2933
tri 428 2855 462 2889 se
rect 462 2855 512 2889
tri 512 2855 546 2889 sw
tri 1008 2855 1042 2889 se
rect 1042 2855 1092 2889
tri 1092 2855 1126 2889 sw
tri 1588 2855 1622 2889 se
rect 1622 2855 1672 2889
tri 1672 2855 1706 2889 sw
tri 2168 2855 2202 2889 se
rect 2202 2855 2252 2889
tri 2252 2855 2286 2889 sw
tri 2748 2855 2782 2889 se
rect 2782 2855 2832 2889
tri 2832 2855 2866 2889 sw
tri 3328 2855 3362 2889 se
rect 3362 2855 3412 2889
tri 3412 2855 3446 2889 sw
tri 3908 2855 3942 2889 se
rect 3942 2855 3992 2889
tri 3992 2855 4026 2889 sw
tri 4488 2855 4522 2889 se
rect 4522 2855 4572 2889
tri 4572 2855 4606 2889 sw
tri 5068 2855 5102 2889 se
rect 5102 2855 5152 2889
tri 5152 2855 5186 2889 sw
tri 5648 2855 5682 2889 se
rect 5682 2855 5732 2889
tri 5732 2855 5766 2889 sw
tri 6228 2855 6262 2889 se
rect 6262 2855 6312 2889
tri 6312 2855 6346 2889 sw
tri 6808 2855 6842 2889 se
rect 6842 2855 6892 2889
tri 6892 2855 6926 2889 sw
tri 402 2829 428 2855 se
rect 428 2829 446 2855
tri 446 2829 472 2855 nw
tri 502 2829 528 2855 ne
rect 528 2829 546 2855
tri 546 2829 572 2855 sw
tri 982 2829 1008 2855 se
rect 1008 2829 1026 2855
tri 1026 2829 1052 2855 nw
tri 1082 2829 1108 2855 ne
rect 1108 2829 1126 2855
tri 1126 2829 1152 2855 sw
tri 1562 2829 1588 2855 se
rect 1588 2829 1606 2855
tri 1606 2829 1632 2855 nw
tri 1662 2829 1688 2855 ne
rect 1688 2829 1706 2855
tri 1706 2829 1732 2855 sw
tri 2142 2829 2168 2855 se
rect 2168 2829 2186 2855
tri 2186 2829 2212 2855 nw
tri 2242 2829 2268 2855 ne
rect 2268 2829 2286 2855
tri 2286 2829 2312 2855 sw
tri 2722 2829 2748 2855 se
rect 2748 2829 2766 2855
tri 2766 2829 2792 2855 nw
tri 2822 2829 2848 2855 ne
rect 2848 2829 2866 2855
tri 2866 2829 2892 2855 sw
tri 3302 2829 3328 2855 se
rect 3328 2829 3346 2855
tri 3346 2829 3372 2855 nw
tri 3402 2829 3428 2855 ne
rect 3428 2829 3446 2855
tri 3446 2829 3472 2855 sw
tri 3882 2829 3908 2855 se
rect 3908 2829 3926 2855
tri 3926 2829 3952 2855 nw
tri 3982 2829 4008 2855 ne
rect 4008 2829 4026 2855
tri 4026 2829 4052 2855 sw
tri 4462 2829 4488 2855 se
rect 4488 2829 4506 2855
tri 4506 2829 4532 2855 nw
tri 4562 2829 4588 2855 ne
rect 4588 2829 4606 2855
tri 4606 2829 4632 2855 sw
tri 5042 2829 5068 2855 se
rect 5068 2829 5086 2855
tri 5086 2829 5112 2855 nw
tri 5142 2829 5168 2855 ne
rect 5168 2829 5186 2855
tri 5186 2829 5212 2855 sw
tri 5622 2829 5648 2855 se
rect 5648 2829 5666 2855
tri 5666 2829 5692 2855 nw
tri 5722 2829 5748 2855 ne
rect 5748 2829 5766 2855
tri 5766 2829 5792 2855 sw
tri 6202 2829 6228 2855 se
rect 6228 2829 6246 2855
tri 6246 2829 6272 2855 nw
tri 6302 2829 6328 2855 ne
rect 6328 2829 6346 2855
tri 6346 2829 6372 2855 sw
tri 6782 2829 6808 2855 se
rect 6808 2829 6826 2855
tri 6826 2829 6852 2855 nw
tri 6882 2829 6908 2855 ne
rect 6908 2829 6926 2855
tri 6926 2829 6952 2855 sw
rect -91 2795 36 2829
rect 66 2795 412 2829
tri 412 2795 446 2829 nw
tri 528 2795 562 2829 ne
rect 562 2795 616 2829
rect 646 2795 992 2829
tri 992 2795 1026 2829 nw
rect 1105 2795 1196 2829
rect 1226 2795 1572 2829
tri 1572 2795 1606 2829 nw
tri 1688 2795 1722 2829 ne
rect 1722 2795 1776 2829
rect 1806 2795 2152 2829
tri 2152 2795 2186 2829 nw
rect 2265 2795 2356 2829
rect 2386 2795 2732 2829
tri 2732 2795 2766 2829 nw
tri 2848 2795 2882 2829 ne
rect 2882 2795 2936 2829
rect 2966 2795 3312 2829
tri 3312 2795 3346 2829 nw
rect 3425 2795 3516 2829
rect 3546 2795 3892 2829
tri 3892 2795 3926 2829 nw
tri 4008 2795 4042 2829 ne
rect 4042 2795 4096 2829
rect 4126 2795 4472 2829
tri 4472 2795 4506 2829 nw
rect 4585 2795 4676 2829
rect 4706 2795 5052 2829
tri 5052 2795 5086 2829 nw
tri 5168 2795 5202 2829 ne
rect 5202 2795 5256 2829
rect 5286 2795 5632 2829
tri 5632 2795 5666 2829 nw
rect 5745 2795 5836 2829
rect 5866 2795 6212 2829
tri 6212 2795 6246 2829 nw
tri 6328 2795 6362 2829 ne
rect 6362 2795 6416 2829
rect 6446 2795 6792 2829
tri 6792 2795 6826 2829 nw
tri 6908 2795 6942 2829 ne
rect 6942 2795 6952 2829
rect -91 2693 253 2707
rect 285 2693 833 2707
rect 865 2693 1413 2707
rect 1445 2693 1993 2707
rect 2025 2693 2573 2707
rect 2605 2693 3153 2707
rect 3185 2693 3733 2707
rect 3765 2693 4313 2707
rect 4345 2693 4893 2707
rect 4925 2693 5473 2707
rect 5505 2693 6053 2707
rect 6085 2693 6633 2707
rect 6665 2693 6925 2707
rect -91 2649 253 2663
rect 285 2649 833 2663
rect 865 2649 1413 2663
rect 1445 2649 1993 2663
rect 2025 2649 2573 2663
rect 2605 2649 3153 2663
rect 3185 2649 3733 2663
rect 3765 2649 4313 2663
rect 4345 2649 4893 2663
rect 4925 2649 5473 2663
rect 5505 2649 6053 2663
rect 6085 2649 6633 2663
rect 6665 2649 6925 2663
tri 428 2585 462 2619 se
rect 462 2585 512 2619
tri 512 2585 546 2619 sw
tri 1008 2585 1042 2619 se
rect 1042 2585 1092 2619
tri 1092 2585 1126 2619 sw
tri 1588 2585 1622 2619 se
rect 1622 2585 1672 2619
tri 1672 2585 1706 2619 sw
tri 2168 2585 2202 2619 se
rect 2202 2585 2252 2619
tri 2252 2585 2286 2619 sw
tri 2748 2585 2782 2619 se
rect 2782 2585 2832 2619
tri 2832 2585 2866 2619 sw
tri 3328 2585 3362 2619 se
rect 3362 2585 3412 2619
tri 3412 2585 3446 2619 sw
tri 3908 2585 3942 2619 se
rect 3942 2585 3992 2619
tri 3992 2585 4026 2619 sw
tri 4488 2585 4522 2619 se
rect 4522 2585 4572 2619
tri 4572 2585 4606 2619 sw
tri 5068 2585 5102 2619 se
rect 5102 2585 5152 2619
tri 5152 2585 5186 2619 sw
tri 5648 2585 5682 2619 se
rect 5682 2585 5732 2619
tri 5732 2585 5766 2619 sw
tri 6228 2585 6262 2619 se
rect 6262 2585 6312 2619
tri 6312 2585 6346 2619 sw
tri 6808 2585 6842 2619 se
rect 6842 2585 6892 2619
tri 6892 2585 6926 2619 sw
tri 402 2559 428 2585 se
rect 428 2559 446 2585
tri 446 2559 472 2585 nw
tri 502 2559 528 2585 ne
rect 528 2559 546 2585
tri 546 2559 572 2585 sw
tri 982 2559 1008 2585 se
rect 1008 2559 1026 2585
tri 1026 2559 1052 2585 nw
tri 1082 2559 1108 2585 ne
rect 1108 2559 1126 2585
tri 1126 2559 1152 2585 sw
tri 1562 2559 1588 2585 se
rect 1588 2559 1606 2585
tri 1606 2559 1632 2585 nw
tri 1662 2559 1688 2585 ne
rect 1688 2559 1706 2585
tri 1706 2559 1732 2585 sw
tri 2142 2559 2168 2585 se
rect 2168 2559 2186 2585
tri 2186 2559 2212 2585 nw
tri 2242 2559 2268 2585 ne
rect 2268 2559 2286 2585
tri 2286 2559 2312 2585 sw
tri 2722 2559 2748 2585 se
rect 2748 2559 2766 2585
tri 2766 2559 2792 2585 nw
tri 2822 2559 2848 2585 ne
rect 2848 2559 2866 2585
tri 2866 2559 2892 2585 sw
tri 3302 2559 3328 2585 se
rect 3328 2559 3346 2585
tri 3346 2559 3372 2585 nw
tri 3402 2559 3428 2585 ne
rect 3428 2559 3446 2585
tri 3446 2559 3472 2585 sw
tri 3882 2559 3908 2585 se
rect 3908 2559 3926 2585
tri 3926 2559 3952 2585 nw
tri 3982 2559 4008 2585 ne
rect 4008 2559 4026 2585
tri 4026 2559 4052 2585 sw
tri 4462 2559 4488 2585 se
rect 4488 2559 4506 2585
tri 4506 2559 4532 2585 nw
tri 4562 2559 4588 2585 ne
rect 4588 2559 4606 2585
tri 4606 2559 4632 2585 sw
tri 5042 2559 5068 2585 se
rect 5068 2559 5086 2585
tri 5086 2559 5112 2585 nw
tri 5142 2559 5168 2585 ne
rect 5168 2559 5186 2585
tri 5186 2559 5212 2585 sw
tri 5622 2559 5648 2585 se
rect 5648 2559 5666 2585
tri 5666 2559 5692 2585 nw
tri 5722 2559 5748 2585 ne
rect 5748 2559 5766 2585
tri 5766 2559 5792 2585 sw
tri 6202 2559 6228 2585 se
rect 6228 2559 6246 2585
tri 6246 2559 6272 2585 nw
tri 6302 2559 6328 2585 ne
rect 6328 2559 6346 2585
tri 6346 2559 6372 2585 sw
tri 6782 2559 6808 2585 se
rect 6808 2559 6826 2585
tri 6826 2559 6852 2585 nw
tri 6882 2559 6908 2585 ne
rect 6908 2559 6926 2585
tri 6926 2559 6952 2585 sw
rect -91 2525 36 2559
rect 66 2525 412 2559
tri 412 2525 446 2559 nw
tri 528 2525 562 2559 ne
rect 562 2525 616 2559
rect 646 2525 992 2559
tri 992 2525 1026 2559 nw
rect 1105 2525 1196 2559
rect 1226 2525 1572 2559
tri 1572 2525 1606 2559 nw
tri 1688 2525 1722 2559 ne
rect 1722 2525 1776 2559
rect 1806 2525 2152 2559
tri 2152 2525 2186 2559 nw
rect 2265 2525 2356 2559
rect 2386 2525 2732 2559
tri 2732 2525 2766 2559 nw
tri 2848 2525 2882 2559 ne
rect 2882 2525 2936 2559
rect 2966 2525 3312 2559
tri 3312 2525 3346 2559 nw
rect 3425 2525 3516 2559
rect 3546 2525 3892 2559
tri 3892 2525 3926 2559 nw
tri 4008 2525 4042 2559 ne
rect 4042 2525 4096 2559
rect 4126 2525 4472 2559
tri 4472 2525 4506 2559 nw
rect 4585 2525 4676 2559
rect 4706 2525 5052 2559
tri 5052 2525 5086 2559 nw
tri 5168 2525 5202 2559 ne
rect 5202 2525 5256 2559
rect 5286 2525 5632 2559
tri 5632 2525 5666 2559 nw
rect 5745 2525 5836 2559
rect 5866 2525 6212 2559
tri 6212 2525 6246 2559 nw
tri 6328 2525 6362 2559 ne
rect 6362 2525 6416 2559
rect 6446 2525 6792 2559
tri 6792 2525 6826 2559 nw
tri 6908 2525 6942 2559 ne
rect 6942 2525 6952 2559
rect -91 2423 253 2437
rect 285 2423 833 2437
rect 865 2423 1413 2437
rect 1445 2423 1993 2437
rect 2025 2423 2573 2437
rect 2605 2423 3153 2437
rect 3185 2423 3733 2437
rect 3765 2423 4313 2437
rect 4345 2423 4893 2437
rect 4925 2423 5473 2437
rect 5505 2423 6053 2437
rect 6085 2423 6633 2437
rect 6665 2423 6925 2437
rect -91 2379 253 2393
rect 285 2379 833 2393
rect 865 2379 1413 2393
rect 1445 2379 1993 2393
rect 2025 2379 2573 2393
rect 2605 2379 3153 2393
rect 3185 2379 3733 2393
rect 3765 2379 4313 2393
rect 4345 2379 4893 2393
rect 4925 2379 5473 2393
rect 5505 2379 6053 2393
rect 6085 2379 6633 2393
rect 6665 2379 6925 2393
tri 428 2315 462 2349 se
rect 462 2315 512 2349
tri 512 2315 546 2349 sw
tri 1008 2315 1042 2349 se
rect 1042 2315 1092 2349
tri 1092 2315 1126 2349 sw
tri 1588 2315 1622 2349 se
rect 1622 2315 1672 2349
tri 1672 2315 1706 2349 sw
tri 2168 2315 2202 2349 se
rect 2202 2315 2252 2349
tri 2252 2315 2286 2349 sw
tri 2748 2315 2782 2349 se
rect 2782 2315 2832 2349
tri 2832 2315 2866 2349 sw
tri 3328 2315 3362 2349 se
rect 3362 2315 3412 2349
tri 3412 2315 3446 2349 sw
tri 3908 2315 3942 2349 se
rect 3942 2315 3992 2349
tri 3992 2315 4026 2349 sw
tri 4488 2315 4522 2349 se
rect 4522 2315 4572 2349
tri 4572 2315 4606 2349 sw
tri 5068 2315 5102 2349 se
rect 5102 2315 5152 2349
tri 5152 2315 5186 2349 sw
tri 5648 2315 5682 2349 se
rect 5682 2315 5732 2349
tri 5732 2315 5766 2349 sw
tri 6228 2315 6262 2349 se
rect 6262 2315 6312 2349
tri 6312 2315 6346 2349 sw
tri 6808 2315 6842 2349 se
rect 6842 2315 6892 2349
tri 6892 2315 6926 2349 sw
tri 402 2289 428 2315 se
rect 428 2289 446 2315
tri 446 2289 472 2315 nw
tri 502 2289 528 2315 ne
rect 528 2289 546 2315
tri 546 2289 572 2315 sw
tri 982 2289 1008 2315 se
rect 1008 2289 1026 2315
tri 1026 2289 1052 2315 nw
tri 1082 2289 1108 2315 ne
rect 1108 2289 1126 2315
tri 1126 2289 1152 2315 sw
tri 1562 2289 1588 2315 se
rect 1588 2289 1606 2315
tri 1606 2289 1632 2315 nw
tri 1662 2289 1688 2315 ne
rect 1688 2289 1706 2315
tri 1706 2289 1732 2315 sw
tri 2142 2289 2168 2315 se
rect 2168 2289 2186 2315
tri 2186 2289 2212 2315 nw
tri 2242 2289 2268 2315 ne
rect 2268 2289 2286 2315
tri 2286 2289 2312 2315 sw
tri 2722 2289 2748 2315 se
rect 2748 2289 2766 2315
tri 2766 2289 2792 2315 nw
tri 2822 2289 2848 2315 ne
rect 2848 2289 2866 2315
tri 2866 2289 2892 2315 sw
tri 3302 2289 3328 2315 se
rect 3328 2289 3346 2315
tri 3346 2289 3372 2315 nw
tri 3402 2289 3428 2315 ne
rect 3428 2289 3446 2315
tri 3446 2289 3472 2315 sw
tri 3882 2289 3908 2315 se
rect 3908 2289 3926 2315
tri 3926 2289 3952 2315 nw
tri 3982 2289 4008 2315 ne
rect 4008 2289 4026 2315
tri 4026 2289 4052 2315 sw
tri 4462 2289 4488 2315 se
rect 4488 2289 4506 2315
tri 4506 2289 4532 2315 nw
tri 4562 2289 4588 2315 ne
rect 4588 2289 4606 2315
tri 4606 2289 4632 2315 sw
tri 5042 2289 5068 2315 se
rect 5068 2289 5086 2315
tri 5086 2289 5112 2315 nw
tri 5142 2289 5168 2315 ne
rect 5168 2289 5186 2315
tri 5186 2289 5212 2315 sw
tri 5622 2289 5648 2315 se
rect 5648 2289 5666 2315
tri 5666 2289 5692 2315 nw
tri 5722 2289 5748 2315 ne
rect 5748 2289 5766 2315
tri 5766 2289 5792 2315 sw
tri 6202 2289 6228 2315 se
rect 6228 2289 6246 2315
tri 6246 2289 6272 2315 nw
tri 6302 2289 6328 2315 ne
rect 6328 2289 6346 2315
tri 6346 2289 6372 2315 sw
tri 6782 2289 6808 2315 se
rect 6808 2289 6826 2315
tri 6826 2289 6852 2315 nw
tri 6882 2289 6908 2315 ne
rect 6908 2289 6926 2315
tri 6926 2289 6952 2315 sw
rect -91 2255 36 2289
rect 66 2255 412 2289
tri 412 2255 446 2289 nw
tri 528 2255 562 2289 ne
rect 562 2255 616 2289
rect 646 2255 992 2289
tri 992 2255 1026 2289 nw
rect 1105 2255 1196 2289
rect 1226 2255 1572 2289
tri 1572 2255 1606 2289 nw
tri 1688 2255 1722 2289 ne
rect 1722 2255 1776 2289
rect 1806 2255 2152 2289
tri 2152 2255 2186 2289 nw
rect 2265 2255 2356 2289
rect 2386 2255 2732 2289
tri 2732 2255 2766 2289 nw
tri 2848 2255 2882 2289 ne
rect 2882 2255 2936 2289
rect 2966 2255 3312 2289
tri 3312 2255 3346 2289 nw
rect 3425 2255 3516 2289
rect 3546 2255 3892 2289
tri 3892 2255 3926 2289 nw
tri 4008 2255 4042 2289 ne
rect 4042 2255 4096 2289
rect 4126 2255 4472 2289
tri 4472 2255 4506 2289 nw
rect 4585 2255 4676 2289
rect 4706 2255 5052 2289
tri 5052 2255 5086 2289 nw
tri 5168 2255 5202 2289 ne
rect 5202 2255 5256 2289
rect 5286 2255 5632 2289
tri 5632 2255 5666 2289 nw
rect 5745 2255 5836 2289
rect 5866 2255 6212 2289
tri 6212 2255 6246 2289 nw
tri 6328 2255 6362 2289 ne
rect 6362 2255 6416 2289
rect 6446 2255 6792 2289
tri 6792 2255 6826 2289 nw
tri 6908 2255 6942 2289 ne
rect 6942 2255 6952 2289
rect -91 2153 253 2167
rect 285 2153 833 2167
rect 865 2153 1413 2167
rect 1445 2153 1993 2167
rect 2025 2153 2573 2167
rect 2605 2153 3153 2167
rect 3185 2153 3733 2167
rect 3765 2153 4313 2167
rect 4345 2153 4893 2167
rect 4925 2153 5473 2167
rect 5505 2153 6053 2167
rect 6085 2153 6633 2167
rect 6665 2153 6925 2167
rect -91 2109 253 2123
rect 285 2109 833 2123
rect 865 2109 1413 2123
rect 1445 2109 1993 2123
rect 2025 2109 2573 2123
rect 2605 2109 3153 2123
rect 3185 2109 3733 2123
rect 3765 2109 4313 2123
rect 4345 2109 4893 2123
rect 4925 2109 5473 2123
rect 5505 2109 6053 2123
rect 6085 2109 6633 2123
rect 6665 2109 6925 2123
tri 428 2045 462 2079 se
rect 462 2045 512 2079
tri 512 2045 546 2079 sw
tri 1008 2045 1042 2079 se
rect 1042 2045 1092 2079
tri 1092 2045 1126 2079 sw
tri 1588 2045 1622 2079 se
rect 1622 2045 1672 2079
tri 1672 2045 1706 2079 sw
tri 2168 2045 2202 2079 se
rect 2202 2045 2252 2079
tri 2252 2045 2286 2079 sw
tri 2748 2045 2782 2079 se
rect 2782 2045 2832 2079
tri 2832 2045 2866 2079 sw
tri 3328 2045 3362 2079 se
rect 3362 2045 3412 2079
tri 3412 2045 3446 2079 sw
tri 3908 2045 3942 2079 se
rect 3942 2045 3992 2079
tri 3992 2045 4026 2079 sw
tri 4488 2045 4522 2079 se
rect 4522 2045 4572 2079
tri 4572 2045 4606 2079 sw
tri 5068 2045 5102 2079 se
rect 5102 2045 5152 2079
tri 5152 2045 5186 2079 sw
tri 5648 2045 5682 2079 se
rect 5682 2045 5732 2079
tri 5732 2045 5766 2079 sw
tri 6228 2045 6262 2079 se
rect 6262 2045 6312 2079
tri 6312 2045 6346 2079 sw
tri 6808 2045 6842 2079 se
rect 6842 2045 6892 2079
tri 6892 2045 6926 2079 sw
tri 402 2019 428 2045 se
rect 428 2019 446 2045
tri 446 2019 472 2045 nw
tri 502 2019 528 2045 ne
rect 528 2019 546 2045
tri 546 2019 572 2045 sw
tri 982 2019 1008 2045 se
rect 1008 2019 1026 2045
tri 1026 2019 1052 2045 nw
tri 1082 2019 1108 2045 ne
rect 1108 2019 1126 2045
tri 1126 2019 1152 2045 sw
tri 1562 2019 1588 2045 se
rect 1588 2019 1606 2045
tri 1606 2019 1632 2045 nw
tri 1662 2019 1688 2045 ne
rect 1688 2019 1706 2045
tri 1706 2019 1732 2045 sw
tri 2142 2019 2168 2045 se
rect 2168 2019 2186 2045
tri 2186 2019 2212 2045 nw
tri 2242 2019 2268 2045 ne
rect 2268 2019 2286 2045
tri 2286 2019 2312 2045 sw
tri 2722 2019 2748 2045 se
rect 2748 2019 2766 2045
tri 2766 2019 2792 2045 nw
tri 2822 2019 2848 2045 ne
rect 2848 2019 2866 2045
tri 2866 2019 2892 2045 sw
tri 3302 2019 3328 2045 se
rect 3328 2019 3346 2045
tri 3346 2019 3372 2045 nw
tri 3402 2019 3428 2045 ne
rect 3428 2019 3446 2045
tri 3446 2019 3472 2045 sw
tri 3882 2019 3908 2045 se
rect 3908 2019 3926 2045
tri 3926 2019 3952 2045 nw
tri 3982 2019 4008 2045 ne
rect 4008 2019 4026 2045
tri 4026 2019 4052 2045 sw
tri 4462 2019 4488 2045 se
rect 4488 2019 4506 2045
tri 4506 2019 4532 2045 nw
tri 4562 2019 4588 2045 ne
rect 4588 2019 4606 2045
tri 4606 2019 4632 2045 sw
tri 5042 2019 5068 2045 se
rect 5068 2019 5086 2045
tri 5086 2019 5112 2045 nw
tri 5142 2019 5168 2045 ne
rect 5168 2019 5186 2045
tri 5186 2019 5212 2045 sw
tri 5622 2019 5648 2045 se
rect 5648 2019 5666 2045
tri 5666 2019 5692 2045 nw
tri 5722 2019 5748 2045 ne
rect 5748 2019 5766 2045
tri 5766 2019 5792 2045 sw
tri 6202 2019 6228 2045 se
rect 6228 2019 6246 2045
tri 6246 2019 6272 2045 nw
tri 6302 2019 6328 2045 ne
rect 6328 2019 6346 2045
tri 6346 2019 6372 2045 sw
tri 6782 2019 6808 2045 se
rect 6808 2019 6826 2045
tri 6826 2019 6852 2045 nw
tri 6882 2019 6908 2045 ne
rect 6908 2019 6926 2045
tri 6926 2019 6952 2045 sw
rect -91 1985 36 2019
rect 66 1985 412 2019
tri 412 1985 446 2019 nw
tri 528 1985 562 2019 ne
rect 562 1985 616 2019
rect 646 1985 992 2019
tri 992 1985 1026 2019 nw
rect 1105 1985 1196 2019
rect 1226 1985 1572 2019
tri 1572 1985 1606 2019 nw
tri 1688 1985 1722 2019 ne
rect 1722 1985 1776 2019
rect 1806 1985 2152 2019
tri 2152 1985 2186 2019 nw
rect 2265 1985 2356 2019
rect 2386 1985 2732 2019
tri 2732 1985 2766 2019 nw
tri 2848 1985 2882 2019 ne
rect 2882 1985 2936 2019
rect 2966 1985 3312 2019
tri 3312 1985 3346 2019 nw
rect 3425 1985 3516 2019
rect 3546 1985 3892 2019
tri 3892 1985 3926 2019 nw
tri 4008 1985 4042 2019 ne
rect 4042 1985 4096 2019
rect 4126 1985 4472 2019
tri 4472 1985 4506 2019 nw
rect 4585 1985 4676 2019
rect 4706 1985 5052 2019
tri 5052 1985 5086 2019 nw
tri 5168 1985 5202 2019 ne
rect 5202 1985 5256 2019
rect 5286 1985 5632 2019
tri 5632 1985 5666 2019 nw
rect 5745 1985 5836 2019
rect 5866 1985 6212 2019
tri 6212 1985 6246 2019 nw
tri 6328 1985 6362 2019 ne
rect 6362 1985 6416 2019
rect 6446 1985 6792 2019
tri 6792 1985 6826 2019 nw
tri 6908 1985 6942 2019 ne
rect 6942 1985 6952 2019
rect -91 1883 253 1897
rect 285 1883 833 1897
rect 865 1883 1413 1897
rect 1445 1883 1993 1897
rect 2025 1883 2573 1897
rect 2605 1883 3153 1897
rect 3185 1883 3733 1897
rect 3765 1883 4313 1897
rect 4345 1883 4893 1897
rect 4925 1883 5473 1897
rect 5505 1883 6053 1897
rect 6085 1883 6633 1897
rect 6665 1883 6925 1897
rect -91 1839 253 1853
rect 285 1839 833 1853
rect 865 1839 1413 1853
rect 1445 1839 1993 1853
rect 2025 1839 2573 1853
rect 2605 1839 3153 1853
rect 3185 1839 3733 1853
rect 3765 1839 4313 1853
rect 4345 1839 4893 1853
rect 4925 1839 5473 1853
rect 5505 1839 6053 1853
rect 6085 1839 6633 1853
rect 6665 1839 6925 1853
tri 428 1775 462 1809 se
rect 462 1775 512 1809
tri 512 1775 546 1809 sw
tri 1008 1775 1042 1809 se
rect 1042 1775 1092 1809
tri 1092 1775 1126 1809 sw
tri 1588 1775 1622 1809 se
rect 1622 1775 1672 1809
tri 1672 1775 1706 1809 sw
tri 2168 1775 2202 1809 se
rect 2202 1775 2252 1809
tri 2252 1775 2286 1809 sw
tri 2748 1775 2782 1809 se
rect 2782 1775 2832 1809
tri 2832 1775 2866 1809 sw
tri 3328 1775 3362 1809 se
rect 3362 1775 3412 1809
tri 3412 1775 3446 1809 sw
tri 3908 1775 3942 1809 se
rect 3942 1775 3992 1809
tri 3992 1775 4026 1809 sw
tri 4488 1775 4522 1809 se
rect 4522 1775 4572 1809
tri 4572 1775 4606 1809 sw
tri 5068 1775 5102 1809 se
rect 5102 1775 5152 1809
tri 5152 1775 5186 1809 sw
tri 5648 1775 5682 1809 se
rect 5682 1775 5732 1809
tri 5732 1775 5766 1809 sw
tri 6228 1775 6262 1809 se
rect 6262 1775 6312 1809
tri 6312 1775 6346 1809 sw
tri 6808 1775 6842 1809 se
rect 6842 1775 6892 1809
tri 6892 1775 6926 1809 sw
tri 402 1749 428 1775 se
rect 428 1749 446 1775
tri 446 1749 472 1775 nw
tri 502 1749 528 1775 ne
rect 528 1749 546 1775
tri 546 1749 572 1775 sw
tri 982 1749 1008 1775 se
rect 1008 1749 1026 1775
tri 1026 1749 1052 1775 nw
tri 1082 1749 1108 1775 ne
rect 1108 1749 1126 1775
tri 1126 1749 1152 1775 sw
tri 1562 1749 1588 1775 se
rect 1588 1749 1606 1775
tri 1606 1749 1632 1775 nw
tri 1662 1749 1688 1775 ne
rect 1688 1749 1706 1775
tri 1706 1749 1732 1775 sw
tri 2142 1749 2168 1775 se
rect 2168 1749 2186 1775
tri 2186 1749 2212 1775 nw
tri 2242 1749 2268 1775 ne
rect 2268 1749 2286 1775
tri 2286 1749 2312 1775 sw
tri 2722 1749 2748 1775 se
rect 2748 1749 2766 1775
tri 2766 1749 2792 1775 nw
tri 2822 1749 2848 1775 ne
rect 2848 1749 2866 1775
tri 2866 1749 2892 1775 sw
tri 3302 1749 3328 1775 se
rect 3328 1749 3346 1775
tri 3346 1749 3372 1775 nw
tri 3402 1749 3428 1775 ne
rect 3428 1749 3446 1775
tri 3446 1749 3472 1775 sw
tri 3882 1749 3908 1775 se
rect 3908 1749 3926 1775
tri 3926 1749 3952 1775 nw
tri 3982 1749 4008 1775 ne
rect 4008 1749 4026 1775
tri 4026 1749 4052 1775 sw
tri 4462 1749 4488 1775 se
rect 4488 1749 4506 1775
tri 4506 1749 4532 1775 nw
tri 4562 1749 4588 1775 ne
rect 4588 1749 4606 1775
tri 4606 1749 4632 1775 sw
tri 5042 1749 5068 1775 se
rect 5068 1749 5086 1775
tri 5086 1749 5112 1775 nw
tri 5142 1749 5168 1775 ne
rect 5168 1749 5186 1775
tri 5186 1749 5212 1775 sw
tri 5622 1749 5648 1775 se
rect 5648 1749 5666 1775
tri 5666 1749 5692 1775 nw
tri 5722 1749 5748 1775 ne
rect 5748 1749 5766 1775
tri 5766 1749 5792 1775 sw
tri 6202 1749 6228 1775 se
rect 6228 1749 6246 1775
tri 6246 1749 6272 1775 nw
tri 6302 1749 6328 1775 ne
rect 6328 1749 6346 1775
tri 6346 1749 6372 1775 sw
tri 6782 1749 6808 1775 se
rect 6808 1749 6826 1775
tri 6826 1749 6852 1775 nw
tri 6882 1749 6908 1775 ne
rect 6908 1749 6926 1775
tri 6926 1749 6952 1775 sw
rect -91 1715 36 1749
rect 66 1715 412 1749
tri 412 1715 446 1749 nw
tri 528 1715 562 1749 ne
rect 562 1715 616 1749
rect 646 1715 992 1749
tri 992 1715 1026 1749 nw
rect 1105 1715 1196 1749
rect 1226 1715 1572 1749
tri 1572 1715 1606 1749 nw
tri 1688 1715 1722 1749 ne
rect 1722 1715 1776 1749
rect 1806 1715 2152 1749
tri 2152 1715 2186 1749 nw
rect 2265 1715 2356 1749
rect 2386 1715 2732 1749
tri 2732 1715 2766 1749 nw
tri 2848 1715 2882 1749 ne
rect 2882 1715 2936 1749
rect 2966 1715 3312 1749
tri 3312 1715 3346 1749 nw
rect 3425 1715 3516 1749
rect 3546 1715 3892 1749
tri 3892 1715 3926 1749 nw
tri 4008 1715 4042 1749 ne
rect 4042 1715 4096 1749
rect 4126 1715 4472 1749
tri 4472 1715 4506 1749 nw
rect 4585 1715 4676 1749
rect 4706 1715 5052 1749
tri 5052 1715 5086 1749 nw
tri 5168 1715 5202 1749 ne
rect 5202 1715 5256 1749
rect 5286 1715 5632 1749
tri 5632 1715 5666 1749 nw
rect 5745 1715 5836 1749
rect 5866 1715 6212 1749
tri 6212 1715 6246 1749 nw
tri 6328 1715 6362 1749 ne
rect 6362 1715 6416 1749
rect 6446 1715 6792 1749
tri 6792 1715 6826 1749 nw
tri 6908 1715 6942 1749 ne
rect 6942 1715 6952 1749
rect -91 1613 253 1627
rect 285 1613 833 1627
rect 865 1613 1413 1627
rect 1445 1613 1993 1627
rect 2025 1613 2573 1627
rect 2605 1613 3153 1627
rect 3185 1613 3733 1627
rect 3765 1613 4313 1627
rect 4345 1613 4893 1627
rect 4925 1613 5473 1627
rect 5505 1613 6053 1627
rect 6085 1613 6633 1627
rect 6665 1613 6925 1627
rect -91 1569 253 1583
rect 285 1569 833 1583
rect 865 1569 1413 1583
rect 1445 1569 1993 1583
rect 2025 1569 2573 1583
rect 2605 1569 3153 1583
rect 3185 1569 3733 1583
rect 3765 1569 4313 1583
rect 4345 1569 4893 1583
rect 4925 1569 5473 1583
rect 5505 1569 6053 1583
rect 6085 1569 6633 1583
rect 6665 1569 6925 1583
tri 428 1505 462 1539 se
rect 462 1505 512 1539
tri 512 1505 546 1539 sw
tri 1008 1505 1042 1539 se
rect 1042 1505 1092 1539
tri 1092 1505 1126 1539 sw
tri 1588 1505 1622 1539 se
rect 1622 1505 1672 1539
tri 1672 1505 1706 1539 sw
tri 2168 1505 2202 1539 se
rect 2202 1505 2252 1539
tri 2252 1505 2286 1539 sw
tri 2748 1505 2782 1539 se
rect 2782 1505 2832 1539
tri 2832 1505 2866 1539 sw
tri 3328 1505 3362 1539 se
rect 3362 1505 3412 1539
tri 3412 1505 3446 1539 sw
tri 3908 1505 3942 1539 se
rect 3942 1505 3992 1539
tri 3992 1505 4026 1539 sw
tri 4488 1505 4522 1539 se
rect 4522 1505 4572 1539
tri 4572 1505 4606 1539 sw
tri 5068 1505 5102 1539 se
rect 5102 1505 5152 1539
tri 5152 1505 5186 1539 sw
tri 5648 1505 5682 1539 se
rect 5682 1505 5732 1539
tri 5732 1505 5766 1539 sw
tri 6228 1505 6262 1539 se
rect 6262 1505 6312 1539
tri 6312 1505 6346 1539 sw
tri 6808 1505 6842 1539 se
rect 6842 1505 6892 1539
tri 6892 1505 6926 1539 sw
tri 402 1479 428 1505 se
rect 428 1479 446 1505
tri 446 1479 472 1505 nw
tri 502 1479 528 1505 ne
rect 528 1479 546 1505
tri 546 1479 572 1505 sw
tri 982 1479 1008 1505 se
rect 1008 1479 1026 1505
tri 1026 1479 1052 1505 nw
tri 1082 1479 1108 1505 ne
rect 1108 1479 1126 1505
tri 1126 1479 1152 1505 sw
tri 1562 1479 1588 1505 se
rect 1588 1479 1606 1505
tri 1606 1479 1632 1505 nw
tri 1662 1479 1688 1505 ne
rect 1688 1479 1706 1505
tri 1706 1479 1732 1505 sw
tri 2142 1479 2168 1505 se
rect 2168 1479 2186 1505
tri 2186 1479 2212 1505 nw
tri 2242 1479 2268 1505 ne
rect 2268 1479 2286 1505
tri 2286 1479 2312 1505 sw
tri 2722 1479 2748 1505 se
rect 2748 1479 2766 1505
tri 2766 1479 2792 1505 nw
tri 2822 1479 2848 1505 ne
rect 2848 1479 2866 1505
tri 2866 1479 2892 1505 sw
tri 3302 1479 3328 1505 se
rect 3328 1479 3346 1505
tri 3346 1479 3372 1505 nw
tri 3402 1479 3428 1505 ne
rect 3428 1479 3446 1505
tri 3446 1479 3472 1505 sw
tri 3882 1479 3908 1505 se
rect 3908 1479 3926 1505
tri 3926 1479 3952 1505 nw
tri 3982 1479 4008 1505 ne
rect 4008 1479 4026 1505
tri 4026 1479 4052 1505 sw
tri 4462 1479 4488 1505 se
rect 4488 1479 4506 1505
tri 4506 1479 4532 1505 nw
tri 4562 1479 4588 1505 ne
rect 4588 1479 4606 1505
tri 4606 1479 4632 1505 sw
tri 5042 1479 5068 1505 se
rect 5068 1479 5086 1505
tri 5086 1479 5112 1505 nw
tri 5142 1479 5168 1505 ne
rect 5168 1479 5186 1505
tri 5186 1479 5212 1505 sw
tri 5622 1479 5648 1505 se
rect 5648 1479 5666 1505
tri 5666 1479 5692 1505 nw
tri 5722 1479 5748 1505 ne
rect 5748 1479 5766 1505
tri 5766 1479 5792 1505 sw
tri 6202 1479 6228 1505 se
rect 6228 1479 6246 1505
tri 6246 1479 6272 1505 nw
tri 6302 1479 6328 1505 ne
rect 6328 1479 6346 1505
tri 6346 1479 6372 1505 sw
tri 6782 1479 6808 1505 se
rect 6808 1479 6826 1505
tri 6826 1479 6852 1505 nw
tri 6882 1479 6908 1505 ne
rect 6908 1479 6926 1505
tri 6926 1479 6952 1505 sw
rect -91 1445 36 1479
rect 66 1445 412 1479
tri 412 1445 446 1479 nw
tri 528 1445 562 1479 ne
rect 562 1445 616 1479
rect 646 1445 992 1479
tri 992 1445 1026 1479 nw
rect 1105 1445 1196 1479
rect 1226 1445 1572 1479
tri 1572 1445 1606 1479 nw
tri 1688 1445 1722 1479 ne
rect 1722 1445 1776 1479
rect 1806 1445 2152 1479
tri 2152 1445 2186 1479 nw
rect 2265 1445 2356 1479
rect 2386 1445 2732 1479
tri 2732 1445 2766 1479 nw
tri 2848 1445 2882 1479 ne
rect 2882 1445 2936 1479
rect 2966 1445 3312 1479
tri 3312 1445 3346 1479 nw
rect 3425 1445 3516 1479
rect 3546 1445 3892 1479
tri 3892 1445 3926 1479 nw
tri 4008 1445 4042 1479 ne
rect 4042 1445 4096 1479
rect 4126 1445 4472 1479
tri 4472 1445 4506 1479 nw
rect 4585 1445 4676 1479
rect 4706 1445 5052 1479
tri 5052 1445 5086 1479 nw
tri 5168 1445 5202 1479 ne
rect 5202 1445 5256 1479
rect 5286 1445 5632 1479
tri 5632 1445 5666 1479 nw
rect 5745 1445 5836 1479
rect 5866 1445 6212 1479
tri 6212 1445 6246 1479 nw
tri 6328 1445 6362 1479 ne
rect 6362 1445 6416 1479
rect 6446 1445 6792 1479
tri 6792 1445 6826 1479 nw
tri 6908 1445 6942 1479 ne
rect 6942 1445 6952 1479
rect -91 1343 253 1357
rect 285 1343 833 1357
rect 865 1343 1413 1357
rect 1445 1343 1993 1357
rect 2025 1343 2573 1357
rect 2605 1343 3153 1357
rect 3185 1343 3733 1357
rect 3765 1343 4313 1357
rect 4345 1343 4893 1357
rect 4925 1343 5473 1357
rect 5505 1343 6053 1357
rect 6085 1343 6633 1357
rect 6665 1343 6925 1357
rect -91 1299 253 1313
rect 285 1299 833 1313
rect 865 1299 1413 1313
rect 1445 1299 1993 1313
rect 2025 1299 2573 1313
rect 2605 1299 3153 1313
rect 3185 1299 3733 1313
rect 3765 1299 4313 1313
rect 4345 1299 4893 1313
rect 4925 1299 5473 1313
rect 5505 1299 6053 1313
rect 6085 1299 6633 1313
rect 6665 1299 6925 1313
tri 428 1235 462 1269 se
rect 462 1235 512 1269
tri 512 1235 546 1269 sw
tri 1008 1235 1042 1269 se
rect 1042 1235 1092 1269
tri 1092 1235 1126 1269 sw
tri 1588 1235 1622 1269 se
rect 1622 1235 1672 1269
tri 1672 1235 1706 1269 sw
tri 2168 1235 2202 1269 se
rect 2202 1235 2252 1269
tri 2252 1235 2286 1269 sw
tri 2748 1235 2782 1269 se
rect 2782 1235 2832 1269
tri 2832 1235 2866 1269 sw
tri 3328 1235 3362 1269 se
rect 3362 1235 3412 1269
tri 3412 1235 3446 1269 sw
tri 3908 1235 3942 1269 se
rect 3942 1235 3992 1269
tri 3992 1235 4026 1269 sw
tri 4488 1235 4522 1269 se
rect 4522 1235 4572 1269
tri 4572 1235 4606 1269 sw
tri 5068 1235 5102 1269 se
rect 5102 1235 5152 1269
tri 5152 1235 5186 1269 sw
tri 5648 1235 5682 1269 se
rect 5682 1235 5732 1269
tri 5732 1235 5766 1269 sw
tri 6228 1235 6262 1269 se
rect 6262 1235 6312 1269
tri 6312 1235 6346 1269 sw
tri 6808 1235 6842 1269 se
rect 6842 1235 6892 1269
tri 6892 1235 6926 1269 sw
tri 402 1209 428 1235 se
rect 428 1209 446 1235
tri 446 1209 472 1235 nw
tri 502 1209 528 1235 ne
rect 528 1209 546 1235
tri 546 1209 572 1235 sw
tri 982 1209 1008 1235 se
rect 1008 1209 1026 1235
tri 1026 1209 1052 1235 nw
tri 1082 1209 1108 1235 ne
rect 1108 1209 1126 1235
tri 1126 1209 1152 1235 sw
tri 1562 1209 1588 1235 se
rect 1588 1209 1606 1235
tri 1606 1209 1632 1235 nw
tri 1662 1209 1688 1235 ne
rect 1688 1209 1706 1235
tri 1706 1209 1732 1235 sw
tri 2142 1209 2168 1235 se
rect 2168 1209 2186 1235
tri 2186 1209 2212 1235 nw
tri 2242 1209 2268 1235 ne
rect 2268 1209 2286 1235
tri 2286 1209 2312 1235 sw
tri 2722 1209 2748 1235 se
rect 2748 1209 2766 1235
tri 2766 1209 2792 1235 nw
tri 2822 1209 2848 1235 ne
rect 2848 1209 2866 1235
tri 2866 1209 2892 1235 sw
tri 3302 1209 3328 1235 se
rect 3328 1209 3346 1235
tri 3346 1209 3372 1235 nw
tri 3402 1209 3428 1235 ne
rect 3428 1209 3446 1235
tri 3446 1209 3472 1235 sw
tri 3882 1209 3908 1235 se
rect 3908 1209 3926 1235
tri 3926 1209 3952 1235 nw
tri 3982 1209 4008 1235 ne
rect 4008 1209 4026 1235
tri 4026 1209 4052 1235 sw
tri 4462 1209 4488 1235 se
rect 4488 1209 4506 1235
tri 4506 1209 4532 1235 nw
tri 4562 1209 4588 1235 ne
rect 4588 1209 4606 1235
tri 4606 1209 4632 1235 sw
tri 5042 1209 5068 1235 se
rect 5068 1209 5086 1235
tri 5086 1209 5112 1235 nw
tri 5142 1209 5168 1235 ne
rect 5168 1209 5186 1235
tri 5186 1209 5212 1235 sw
tri 5622 1209 5648 1235 se
rect 5648 1209 5666 1235
tri 5666 1209 5692 1235 nw
tri 5722 1209 5748 1235 ne
rect 5748 1209 5766 1235
tri 5766 1209 5792 1235 sw
tri 6202 1209 6228 1235 se
rect 6228 1209 6246 1235
tri 6246 1209 6272 1235 nw
tri 6302 1209 6328 1235 ne
rect 6328 1209 6346 1235
tri 6346 1209 6372 1235 sw
tri 6782 1209 6808 1235 se
rect 6808 1209 6826 1235
tri 6826 1209 6852 1235 nw
tri 6882 1209 6908 1235 ne
rect 6908 1209 6926 1235
tri 6926 1209 6952 1235 sw
rect -91 1175 36 1209
rect 66 1175 412 1209
tri 412 1175 446 1209 nw
tri 528 1175 562 1209 ne
rect 562 1175 616 1209
rect 646 1175 992 1209
tri 992 1175 1026 1209 nw
rect 1105 1175 1196 1209
rect 1226 1175 1572 1209
tri 1572 1175 1606 1209 nw
tri 1688 1175 1722 1209 ne
rect 1722 1175 1776 1209
rect 1806 1175 2152 1209
tri 2152 1175 2186 1209 nw
rect 2265 1175 2356 1209
rect 2386 1175 2732 1209
tri 2732 1175 2766 1209 nw
tri 2848 1175 2882 1209 ne
rect 2882 1175 2936 1209
rect 2966 1175 3312 1209
tri 3312 1175 3346 1209 nw
rect 3425 1175 3516 1209
rect 3546 1175 3892 1209
tri 3892 1175 3926 1209 nw
tri 4008 1175 4042 1209 ne
rect 4042 1175 4096 1209
rect 4126 1175 4472 1209
tri 4472 1175 4506 1209 nw
rect 4585 1175 4676 1209
rect 4706 1175 5052 1209
tri 5052 1175 5086 1209 nw
tri 5168 1175 5202 1209 ne
rect 5202 1175 5256 1209
rect 5286 1175 5632 1209
tri 5632 1175 5666 1209 nw
rect 5745 1175 5836 1209
rect 5866 1175 6212 1209
tri 6212 1175 6246 1209 nw
tri 6328 1175 6362 1209 ne
rect 6362 1175 6416 1209
rect 6446 1175 6792 1209
tri 6792 1175 6826 1209 nw
tri 6908 1175 6942 1209 ne
rect 6942 1175 6952 1209
rect -91 1073 253 1087
rect 285 1073 833 1087
rect 865 1073 1413 1087
rect 1445 1073 1993 1087
rect 2025 1073 2573 1087
rect 2605 1073 3153 1087
rect 3185 1073 3733 1087
rect 3765 1073 4313 1087
rect 4345 1073 4893 1087
rect 4925 1073 5473 1087
rect 5505 1073 6053 1087
rect 6085 1073 6633 1087
rect 6665 1073 6925 1087
rect -91 1029 253 1043
rect 285 1029 833 1043
rect 865 1029 1413 1043
rect 1445 1029 1993 1043
rect 2025 1029 2573 1043
rect 2605 1029 3153 1043
rect 3185 1029 3733 1043
rect 3765 1029 4313 1043
rect 4345 1029 4893 1043
rect 4925 1029 5473 1043
rect 5505 1029 6053 1043
rect 6085 1029 6633 1043
rect 6665 1029 6925 1043
tri 428 965 462 999 se
rect 462 965 512 999
tri 512 965 546 999 sw
tri 1008 965 1042 999 se
rect 1042 965 1092 999
tri 1092 965 1126 999 sw
tri 1588 965 1622 999 se
rect 1622 965 1672 999
tri 1672 965 1706 999 sw
tri 2168 965 2202 999 se
rect 2202 965 2252 999
tri 2252 965 2286 999 sw
tri 2748 965 2782 999 se
rect 2782 965 2832 999
tri 2832 965 2866 999 sw
tri 3328 965 3362 999 se
rect 3362 965 3412 999
tri 3412 965 3446 999 sw
tri 3908 965 3942 999 se
rect 3942 965 3992 999
tri 3992 965 4026 999 sw
tri 4488 965 4522 999 se
rect 4522 965 4572 999
tri 4572 965 4606 999 sw
tri 5068 965 5102 999 se
rect 5102 965 5152 999
tri 5152 965 5186 999 sw
tri 5648 965 5682 999 se
rect 5682 965 5732 999
tri 5732 965 5766 999 sw
tri 6228 965 6262 999 se
rect 6262 965 6312 999
tri 6312 965 6346 999 sw
tri 6808 965 6842 999 se
rect 6842 965 6892 999
tri 6892 965 6926 999 sw
tri 402 939 428 965 se
rect 428 939 446 965
tri 446 939 472 965 nw
tri 502 939 528 965 ne
rect 528 939 546 965
tri 546 939 572 965 sw
tri 982 939 1008 965 se
rect 1008 939 1026 965
tri 1026 939 1052 965 nw
tri 1082 939 1108 965 ne
rect 1108 939 1126 965
tri 1126 939 1152 965 sw
tri 1562 939 1588 965 se
rect 1588 939 1606 965
tri 1606 939 1632 965 nw
tri 1662 939 1688 965 ne
rect 1688 939 1706 965
tri 1706 939 1732 965 sw
tri 2142 939 2168 965 se
rect 2168 939 2186 965
tri 2186 939 2212 965 nw
tri 2242 939 2268 965 ne
rect 2268 939 2286 965
tri 2286 939 2312 965 sw
tri 2722 939 2748 965 se
rect 2748 939 2766 965
tri 2766 939 2792 965 nw
tri 2822 939 2848 965 ne
rect 2848 939 2866 965
tri 2866 939 2892 965 sw
tri 3302 939 3328 965 se
rect 3328 939 3346 965
tri 3346 939 3372 965 nw
tri 3402 939 3428 965 ne
rect 3428 939 3446 965
tri 3446 939 3472 965 sw
tri 3882 939 3908 965 se
rect 3908 939 3926 965
tri 3926 939 3952 965 nw
tri 3982 939 4008 965 ne
rect 4008 939 4026 965
tri 4026 939 4052 965 sw
tri 4462 939 4488 965 se
rect 4488 939 4506 965
tri 4506 939 4532 965 nw
tri 4562 939 4588 965 ne
rect 4588 939 4606 965
tri 4606 939 4632 965 sw
tri 5042 939 5068 965 se
rect 5068 939 5086 965
tri 5086 939 5112 965 nw
tri 5142 939 5168 965 ne
rect 5168 939 5186 965
tri 5186 939 5212 965 sw
tri 5622 939 5648 965 se
rect 5648 939 5666 965
tri 5666 939 5692 965 nw
tri 5722 939 5748 965 ne
rect 5748 939 5766 965
tri 5766 939 5792 965 sw
tri 6202 939 6228 965 se
rect 6228 939 6246 965
tri 6246 939 6272 965 nw
tri 6302 939 6328 965 ne
rect 6328 939 6346 965
tri 6346 939 6372 965 sw
tri 6782 939 6808 965 se
rect 6808 939 6826 965
tri 6826 939 6852 965 nw
tri 6882 939 6908 965 ne
rect 6908 939 6926 965
tri 6926 939 6952 965 sw
rect -91 905 36 939
rect 66 905 412 939
tri 412 905 446 939 nw
tri 528 905 562 939 ne
rect 562 905 616 939
rect 646 905 992 939
tri 992 905 1026 939 nw
rect 1105 905 1196 939
rect 1226 905 1572 939
tri 1572 905 1606 939 nw
tri 1688 905 1722 939 ne
rect 1722 905 1776 939
rect 1806 905 2152 939
tri 2152 905 2186 939 nw
rect 2265 905 2356 939
rect 2386 905 2732 939
tri 2732 905 2766 939 nw
tri 2848 905 2882 939 ne
rect 2882 905 2936 939
rect 2966 905 3312 939
tri 3312 905 3346 939 nw
rect 3425 905 3516 939
rect 3546 905 3892 939
tri 3892 905 3926 939 nw
tri 4008 905 4042 939 ne
rect 4042 905 4096 939
rect 4126 905 4472 939
tri 4472 905 4506 939 nw
rect 4585 905 4676 939
rect 4706 905 5052 939
tri 5052 905 5086 939 nw
tri 5168 905 5202 939 ne
rect 5202 905 5256 939
rect 5286 905 5632 939
tri 5632 905 5666 939 nw
rect 5745 905 5836 939
rect 5866 905 6212 939
tri 6212 905 6246 939 nw
tri 6328 905 6362 939 ne
rect 6362 905 6416 939
rect 6446 905 6792 939
tri 6792 905 6826 939 nw
tri 6908 905 6942 939 ne
rect 6942 905 6952 939
rect -91 803 253 817
rect 285 803 833 817
rect 865 803 1413 817
rect 1445 803 1993 817
rect 2025 803 2573 817
rect 2605 803 3153 817
rect 3185 803 3733 817
rect 3765 803 4313 817
rect 4345 803 4893 817
rect 4925 803 5473 817
rect 5505 803 6053 817
rect 6085 803 6633 817
rect 6665 803 6925 817
rect -91 759 253 773
rect 285 759 833 773
rect 865 759 1413 773
rect 1445 759 1993 773
rect 2025 759 2573 773
rect 2605 759 3153 773
rect 3185 759 3733 773
rect 3765 759 4313 773
rect 4345 759 4893 773
rect 4925 759 5473 773
rect 5505 759 6053 773
rect 6085 759 6633 773
rect 6665 759 6925 773
tri 428 695 462 729 se
rect 462 695 512 729
tri 512 695 546 729 sw
tri 1008 695 1042 729 se
rect 1042 695 1092 729
tri 1092 695 1126 729 sw
tri 1588 695 1622 729 se
rect 1622 695 1672 729
tri 1672 695 1706 729 sw
tri 2168 695 2202 729 se
rect 2202 695 2252 729
tri 2252 695 2286 729 sw
tri 2748 695 2782 729 se
rect 2782 695 2832 729
tri 2832 695 2866 729 sw
tri 3328 695 3362 729 se
rect 3362 695 3412 729
tri 3412 695 3446 729 sw
tri 3908 695 3942 729 se
rect 3942 695 3992 729
tri 3992 695 4026 729 sw
tri 4488 695 4522 729 se
rect 4522 695 4572 729
tri 4572 695 4606 729 sw
tri 5068 695 5102 729 se
rect 5102 695 5152 729
tri 5152 695 5186 729 sw
tri 5648 695 5682 729 se
rect 5682 695 5732 729
tri 5732 695 5766 729 sw
tri 6228 695 6262 729 se
rect 6262 695 6312 729
tri 6312 695 6346 729 sw
tri 6808 695 6842 729 se
rect 6842 695 6892 729
tri 6892 695 6926 729 sw
tri 402 669 428 695 se
rect 428 669 446 695
tri 446 669 472 695 nw
tri 502 669 528 695 ne
rect 528 669 546 695
tri 546 669 572 695 sw
tri 982 669 1008 695 se
rect 1008 669 1026 695
tri 1026 669 1052 695 nw
tri 1082 669 1108 695 ne
rect 1108 669 1126 695
tri 1126 669 1152 695 sw
tri 1562 669 1588 695 se
rect 1588 669 1606 695
tri 1606 669 1632 695 nw
tri 1662 669 1688 695 ne
rect 1688 669 1706 695
tri 1706 669 1732 695 sw
tri 2142 669 2168 695 se
rect 2168 669 2186 695
tri 2186 669 2212 695 nw
tri 2242 669 2268 695 ne
rect 2268 669 2286 695
tri 2286 669 2312 695 sw
tri 2722 669 2748 695 se
rect 2748 669 2766 695
tri 2766 669 2792 695 nw
tri 2822 669 2848 695 ne
rect 2848 669 2866 695
tri 2866 669 2892 695 sw
tri 3302 669 3328 695 se
rect 3328 669 3346 695
tri 3346 669 3372 695 nw
tri 3402 669 3428 695 ne
rect 3428 669 3446 695
tri 3446 669 3472 695 sw
tri 3882 669 3908 695 se
rect 3908 669 3926 695
tri 3926 669 3952 695 nw
tri 3982 669 4008 695 ne
rect 4008 669 4026 695
tri 4026 669 4052 695 sw
tri 4462 669 4488 695 se
rect 4488 669 4506 695
tri 4506 669 4532 695 nw
tri 4562 669 4588 695 ne
rect 4588 669 4606 695
tri 4606 669 4632 695 sw
tri 5042 669 5068 695 se
rect 5068 669 5086 695
tri 5086 669 5112 695 nw
tri 5142 669 5168 695 ne
rect 5168 669 5186 695
tri 5186 669 5212 695 sw
tri 5622 669 5648 695 se
rect 5648 669 5666 695
tri 5666 669 5692 695 nw
tri 5722 669 5748 695 ne
rect 5748 669 5766 695
tri 5766 669 5792 695 sw
tri 6202 669 6228 695 se
rect 6228 669 6246 695
tri 6246 669 6272 695 nw
tri 6302 669 6328 695 ne
rect 6328 669 6346 695
tri 6346 669 6372 695 sw
tri 6782 669 6808 695 se
rect 6808 669 6826 695
tri 6826 669 6852 695 nw
tri 6882 669 6908 695 ne
rect 6908 669 6926 695
tri 6926 669 6952 695 sw
rect -91 635 36 669
rect 66 635 412 669
tri 412 635 446 669 nw
tri 528 635 562 669 ne
rect 562 635 616 669
rect 646 635 992 669
tri 992 635 1026 669 nw
rect 1105 635 1196 669
rect 1226 635 1572 669
tri 1572 635 1606 669 nw
tri 1688 635 1722 669 ne
rect 1722 635 1776 669
rect 1806 635 2152 669
tri 2152 635 2186 669 nw
rect 2265 635 2356 669
rect 2386 635 2732 669
tri 2732 635 2766 669 nw
tri 2848 635 2882 669 ne
rect 2882 635 2936 669
rect 2966 635 3312 669
tri 3312 635 3346 669 nw
rect 3425 635 3516 669
rect 3546 635 3892 669
tri 3892 635 3926 669 nw
tri 4008 635 4042 669 ne
rect 4042 635 4096 669
rect 4126 635 4472 669
tri 4472 635 4506 669 nw
rect 4585 635 4676 669
rect 4706 635 5052 669
tri 5052 635 5086 669 nw
tri 5168 635 5202 669 ne
rect 5202 635 5256 669
rect 5286 635 5632 669
tri 5632 635 5666 669 nw
rect 5745 635 5836 669
rect 5866 635 6212 669
tri 6212 635 6246 669 nw
tri 6328 635 6362 669 ne
rect 6362 635 6416 669
rect 6446 635 6792 669
tri 6792 635 6826 669 nw
tri 6908 635 6942 669 ne
rect 6942 635 6952 669
rect -91 533 253 547
rect 285 533 833 547
rect 865 533 1413 547
rect 1445 533 1993 547
rect 2025 533 2573 547
rect 2605 533 3153 547
rect 3185 533 3733 547
rect 3765 533 4313 547
rect 4345 533 4893 547
rect 4925 533 5473 547
rect 5505 533 6053 547
rect 6085 533 6633 547
rect 6665 533 6925 547
rect -91 489 253 503
rect 285 489 833 503
rect 865 489 1413 503
rect 1445 489 1993 503
rect 2025 489 2573 503
rect 2605 489 3153 503
rect 3185 489 3733 503
rect 3765 489 4313 503
rect 4345 489 4893 503
rect 4925 489 5473 503
rect 5505 489 6053 503
rect 6085 489 6633 503
rect 6665 489 6925 503
tri 428 425 462 459 se
rect 462 425 512 459
tri 512 425 546 459 sw
tri 1008 425 1042 459 se
rect 1042 425 1092 459
tri 1092 425 1126 459 sw
tri 1588 425 1622 459 se
rect 1622 425 1672 459
tri 1672 425 1706 459 sw
tri 2168 425 2202 459 se
rect 2202 425 2252 459
tri 2252 425 2286 459 sw
tri 2748 425 2782 459 se
rect 2782 425 2832 459
tri 2832 425 2866 459 sw
tri 3328 425 3362 459 se
rect 3362 425 3412 459
tri 3412 425 3446 459 sw
tri 3908 425 3942 459 se
rect 3942 425 3992 459
tri 3992 425 4026 459 sw
tri 4488 425 4522 459 se
rect 4522 425 4572 459
tri 4572 425 4606 459 sw
tri 5068 425 5102 459 se
rect 5102 425 5152 459
tri 5152 425 5186 459 sw
tri 5648 425 5682 459 se
rect 5682 425 5732 459
tri 5732 425 5766 459 sw
tri 6228 425 6262 459 se
rect 6262 425 6312 459
tri 6312 425 6346 459 sw
tri 6808 425 6842 459 se
rect 6842 425 6892 459
tri 6892 425 6926 459 sw
tri 402 399 428 425 se
rect 428 399 446 425
tri 446 399 472 425 nw
tri 502 399 528 425 ne
rect 528 399 546 425
tri 546 399 572 425 sw
tri 982 399 1008 425 se
rect 1008 399 1026 425
tri 1026 399 1052 425 nw
tri 1082 399 1108 425 ne
rect 1108 399 1126 425
tri 1126 399 1152 425 sw
tri 1562 399 1588 425 se
rect 1588 399 1606 425
tri 1606 399 1632 425 nw
tri 1662 399 1688 425 ne
rect 1688 399 1706 425
tri 1706 399 1732 425 sw
tri 2142 399 2168 425 se
rect 2168 399 2186 425
tri 2186 399 2212 425 nw
tri 2242 399 2268 425 ne
rect 2268 399 2286 425
tri 2286 399 2312 425 sw
tri 2722 399 2748 425 se
rect 2748 399 2766 425
tri 2766 399 2792 425 nw
tri 2822 399 2848 425 ne
rect 2848 399 2866 425
tri 2866 399 2892 425 sw
tri 3302 399 3328 425 se
rect 3328 399 3346 425
tri 3346 399 3372 425 nw
tri 3402 399 3428 425 ne
rect 3428 399 3446 425
tri 3446 399 3472 425 sw
tri 3882 399 3908 425 se
rect 3908 399 3926 425
tri 3926 399 3952 425 nw
tri 3982 399 4008 425 ne
rect 4008 399 4026 425
tri 4026 399 4052 425 sw
tri 4462 399 4488 425 se
rect 4488 399 4506 425
tri 4506 399 4532 425 nw
tri 4562 399 4588 425 ne
rect 4588 399 4606 425
tri 4606 399 4632 425 sw
tri 5042 399 5068 425 se
rect 5068 399 5086 425
tri 5086 399 5112 425 nw
tri 5142 399 5168 425 ne
rect 5168 399 5186 425
tri 5186 399 5212 425 sw
tri 5622 399 5648 425 se
rect 5648 399 5666 425
tri 5666 399 5692 425 nw
tri 5722 399 5748 425 ne
rect 5748 399 5766 425
tri 5766 399 5792 425 sw
tri 6202 399 6228 425 se
rect 6228 399 6246 425
tri 6246 399 6272 425 nw
tri 6302 399 6328 425 ne
rect 6328 399 6346 425
tri 6346 399 6372 425 sw
tri 6782 399 6808 425 se
rect 6808 399 6826 425
tri 6826 399 6852 425 nw
tri 6882 399 6908 425 ne
rect 6908 399 6926 425
tri 6926 399 6952 425 sw
rect -91 365 36 399
rect 66 365 412 399
tri 412 365 446 399 nw
tri 528 365 562 399 ne
rect 562 365 616 399
rect 646 365 992 399
tri 992 365 1026 399 nw
rect 1105 365 1196 399
rect 1226 365 1572 399
tri 1572 365 1606 399 nw
tri 1688 365 1722 399 ne
rect 1722 365 1776 399
rect 1806 365 2152 399
tri 2152 365 2186 399 nw
rect 2265 365 2356 399
rect 2386 365 2732 399
tri 2732 365 2766 399 nw
tri 2848 365 2882 399 ne
rect 2882 365 2936 399
rect 2966 365 3312 399
tri 3312 365 3346 399 nw
rect 3425 365 3516 399
rect 3546 365 3892 399
tri 3892 365 3926 399 nw
tri 4008 365 4042 399 ne
rect 4042 365 4096 399
rect 4126 365 4472 399
tri 4472 365 4506 399 nw
rect 4585 365 4676 399
rect 4706 365 5052 399
tri 5052 365 5086 399 nw
tri 5168 365 5202 399 ne
rect 5202 365 5256 399
rect 5286 365 5632 399
tri 5632 365 5666 399 nw
rect 5745 365 5836 399
rect 5866 365 6212 399
tri 6212 365 6246 399 nw
tri 6328 365 6362 399 ne
rect 6362 365 6416 399
rect 6446 365 6792 399
tri 6792 365 6826 399 nw
tri 6908 365 6942 399 ne
rect 6942 365 6952 399
rect -91 263 253 277
rect 285 263 833 277
rect 865 263 1413 277
rect 1445 263 1993 277
rect 2025 263 2573 277
rect 2605 263 3153 277
rect 3185 263 3733 277
rect 3765 263 4313 277
rect 4345 263 4893 277
rect 4925 263 5473 277
rect 5505 263 6053 277
rect 6085 263 6633 277
rect 6665 263 6925 277
rect -91 219 253 233
rect 285 219 833 233
rect 865 219 1413 233
rect 1445 219 1993 233
rect 2025 219 2573 233
rect 2605 219 3153 233
rect 3185 219 3733 233
rect 3765 219 4313 233
rect 4345 219 4893 233
rect 4925 219 5473 233
rect 5505 219 6053 233
rect 6085 219 6633 233
rect 6665 219 6925 233
tri 428 155 462 189 se
rect 462 155 512 189
tri 512 155 546 189 sw
tri 1008 155 1042 189 se
rect 1042 155 1092 189
tri 1092 155 1126 189 sw
tri 1588 155 1622 189 se
rect 1622 155 1672 189
tri 1672 155 1706 189 sw
tri 2168 155 2202 189 se
rect 2202 155 2252 189
tri 2252 155 2286 189 sw
tri 2748 155 2782 189 se
rect 2782 155 2832 189
tri 2832 155 2866 189 sw
tri 3328 155 3362 189 se
rect 3362 155 3412 189
tri 3412 155 3446 189 sw
tri 3908 155 3942 189 se
rect 3942 155 3992 189
tri 3992 155 4026 189 sw
tri 4488 155 4522 189 se
rect 4522 155 4572 189
tri 4572 155 4606 189 sw
tri 5068 155 5102 189 se
rect 5102 155 5152 189
tri 5152 155 5186 189 sw
tri 5648 155 5682 189 se
rect 5682 155 5732 189
tri 5732 155 5766 189 sw
tri 6228 155 6262 189 se
rect 6262 155 6312 189
tri 6312 155 6346 189 sw
tri 6808 155 6842 189 se
rect 6842 155 6892 189
tri 6892 155 6926 189 sw
tri 402 129 428 155 se
rect 428 129 446 155
tri 446 129 472 155 nw
tri 502 129 528 155 ne
rect 528 129 546 155
tri 546 129 572 155 sw
tri 982 129 1008 155 se
rect 1008 129 1026 155
tri 1026 129 1052 155 nw
tri 1082 129 1108 155 ne
rect 1108 129 1126 155
tri 1126 129 1152 155 sw
tri 1562 129 1588 155 se
rect 1588 129 1606 155
tri 1606 129 1632 155 nw
tri 1662 129 1688 155 ne
rect 1688 129 1706 155
tri 1706 129 1732 155 sw
tri 2142 129 2168 155 se
rect 2168 129 2186 155
tri 2186 129 2212 155 nw
tri 2242 129 2268 155 ne
rect 2268 129 2286 155
tri 2286 129 2312 155 sw
tri 2722 129 2748 155 se
rect 2748 129 2766 155
tri 2766 129 2792 155 nw
tri 2822 129 2848 155 ne
rect 2848 129 2866 155
tri 2866 129 2892 155 sw
tri 3302 129 3328 155 se
rect 3328 129 3346 155
tri 3346 129 3372 155 nw
tri 3402 129 3428 155 ne
rect 3428 129 3446 155
tri 3446 129 3472 155 sw
tri 3882 129 3908 155 se
rect 3908 129 3926 155
tri 3926 129 3952 155 nw
tri 3982 129 4008 155 ne
rect 4008 129 4026 155
tri 4026 129 4052 155 sw
tri 4462 129 4488 155 se
rect 4488 129 4506 155
tri 4506 129 4532 155 nw
tri 4562 129 4588 155 ne
rect 4588 129 4606 155
tri 4606 129 4632 155 sw
tri 5042 129 5068 155 se
rect 5068 129 5086 155
tri 5086 129 5112 155 nw
tri 5142 129 5168 155 ne
rect 5168 129 5186 155
tri 5186 129 5212 155 sw
tri 5622 129 5648 155 se
rect 5648 129 5666 155
tri 5666 129 5692 155 nw
tri 5722 129 5748 155 ne
rect 5748 129 5766 155
tri 5766 129 5792 155 sw
tri 6202 129 6228 155 se
rect 6228 129 6246 155
tri 6246 129 6272 155 nw
tri 6302 129 6328 155 ne
rect 6328 129 6346 155
tri 6346 129 6372 155 sw
tri 6782 129 6808 155 se
rect 6808 129 6826 155
tri 6826 129 6852 155 nw
tri 6882 129 6908 155 ne
rect 6908 129 6926 155
tri 6926 129 6952 155 sw
rect -91 95 36 129
rect 66 95 412 129
tri 412 95 446 129 nw
tri 528 95 562 129 ne
rect 562 95 616 129
rect 646 95 992 129
tri 992 95 1026 129 nw
rect 1105 95 1196 129
rect 1226 95 1572 129
tri 1572 95 1606 129 nw
tri 1688 95 1722 129 ne
rect 1722 95 1776 129
rect 1806 95 2152 129
tri 2152 95 2186 129 nw
rect 2265 95 2356 129
rect 2386 95 2732 129
tri 2732 95 2766 129 nw
tri 2848 95 2882 129 ne
rect 2882 95 2936 129
rect 2966 95 3312 129
tri 3312 95 3346 129 nw
rect 3425 95 3516 129
rect 3546 95 3892 129
tri 3892 95 3926 129 nw
tri 4008 95 4042 129 ne
rect 4042 95 4096 129
rect 4126 95 4472 129
tri 4472 95 4506 129 nw
rect 4585 95 4676 129
rect 4706 95 5052 129
tri 5052 95 5086 129 nw
tri 5168 95 5202 129 ne
rect 5202 95 5256 129
rect 5286 95 5632 129
tri 5632 95 5666 129 nw
rect 5745 95 5836 129
rect 5866 95 6212 129
tri 6212 95 6246 129 nw
tri 6328 95 6362 129 ne
rect 6362 95 6416 129
rect 6446 95 6792 129
tri 6792 95 6826 129 nw
tri 6908 95 6942 129 ne
rect 6942 95 6952 129
rect -91 -7 253 7
rect 285 -7 833 7
rect 865 -7 1413 7
rect 1445 -7 1993 7
rect 2025 -7 2573 7
rect 2605 -7 3153 7
rect 3185 -7 3733 7
rect 3765 -7 4313 7
rect 4345 -7 4893 7
rect 4925 -7 5473 7
rect 5505 -7 6053 7
rect 6085 -7 6633 7
rect 6665 -7 6925 7
<< via1 >>
rect 472 4145 502 4179
rect 1052 4145 1082 4179
rect 1632 4146 1662 4179
rect 1632 4145 1662 4146
rect 2212 4145 2242 4179
rect 2792 4146 2822 4179
rect 2792 4145 2822 4146
rect 3372 4145 3402 4179
rect 3952 4146 3982 4179
rect 3952 4145 3982 4146
rect 4532 4145 4562 4179
rect 5112 4146 5142 4179
rect 5112 4145 5142 4146
rect 5692 4145 5722 4179
rect 6272 4146 6302 4179
rect 6272 4145 6302 4146
rect 6852 4145 6882 4179
rect 472 3876 502 3909
rect 472 3875 502 3876
rect 1052 3875 1082 3909
rect 1632 3876 1662 3909
rect 1632 3875 1662 3876
rect 2212 3875 2242 3909
rect 2792 3876 2822 3909
rect 2792 3875 2822 3876
rect 3372 3875 3402 3909
rect 3952 3876 3982 3909
rect 3952 3875 3982 3876
rect 4532 3875 4562 3909
rect 5112 3876 5142 3909
rect 5112 3875 5142 3876
rect 5692 3875 5722 3909
rect 6272 3876 6302 3909
rect 6272 3875 6302 3876
rect 6852 3875 6882 3909
rect 472 3606 502 3639
rect 472 3605 502 3606
rect 1052 3605 1082 3639
rect 1632 3606 1662 3639
rect 1632 3605 1662 3606
rect 2212 3605 2242 3639
rect 2792 3606 2822 3639
rect 2792 3605 2822 3606
rect 3372 3605 3402 3639
rect 3952 3606 3982 3639
rect 3952 3605 3982 3606
rect 4532 3605 4562 3639
rect 5112 3606 5142 3639
rect 5112 3605 5142 3606
rect 5692 3605 5722 3639
rect 6272 3606 6302 3639
rect 6272 3605 6302 3606
rect 6852 3605 6882 3639
rect 472 3336 502 3369
rect 472 3335 502 3336
rect 1052 3335 1082 3369
rect 1632 3336 1662 3369
rect 1632 3335 1662 3336
rect 2212 3335 2242 3369
rect 2792 3336 2822 3369
rect 2792 3335 2822 3336
rect 3372 3335 3402 3369
rect 3952 3336 3982 3369
rect 3952 3335 3982 3336
rect 4532 3335 4562 3369
rect 5112 3336 5142 3369
rect 5112 3335 5142 3336
rect 5692 3335 5722 3369
rect 6272 3336 6302 3369
rect 6272 3335 6302 3336
rect 6852 3335 6882 3369
rect 472 3066 502 3099
rect 472 3065 502 3066
rect 1052 3065 1082 3099
rect 1632 3066 1662 3099
rect 1632 3065 1662 3066
rect 2212 3065 2242 3099
rect 2792 3066 2822 3099
rect 2792 3065 2822 3066
rect 3372 3065 3402 3099
rect 3952 3066 3982 3099
rect 3952 3065 3982 3066
rect 4532 3065 4562 3099
rect 5112 3066 5142 3099
rect 5112 3065 5142 3066
rect 5692 3065 5722 3099
rect 6272 3066 6302 3099
rect 6272 3065 6302 3066
rect 6852 3065 6882 3099
rect 472 2796 502 2829
rect 472 2795 502 2796
rect 1052 2795 1082 2829
rect 1632 2796 1662 2829
rect 1632 2795 1662 2796
rect 2212 2795 2242 2829
rect 2792 2796 2822 2829
rect 2792 2795 2822 2796
rect 3372 2795 3402 2829
rect 3952 2796 3982 2829
rect 3952 2795 3982 2796
rect 4532 2795 4562 2829
rect 5112 2796 5142 2829
rect 5112 2795 5142 2796
rect 5692 2795 5722 2829
rect 6272 2796 6302 2829
rect 6272 2795 6302 2796
rect 6852 2795 6882 2829
rect 472 2526 502 2559
rect 472 2525 502 2526
rect 1052 2525 1082 2559
rect 1632 2526 1662 2559
rect 1632 2525 1662 2526
rect 2212 2525 2242 2559
rect 2792 2526 2822 2559
rect 2792 2525 2822 2526
rect 3372 2525 3402 2559
rect 3952 2526 3982 2559
rect 3952 2525 3982 2526
rect 4532 2525 4562 2559
rect 5112 2526 5142 2559
rect 5112 2525 5142 2526
rect 5692 2525 5722 2559
rect 6272 2526 6302 2559
rect 6272 2525 6302 2526
rect 6852 2525 6882 2559
rect 472 2256 502 2289
rect 472 2255 502 2256
rect 1052 2255 1082 2289
rect 1632 2256 1662 2289
rect 1632 2255 1662 2256
rect 2212 2255 2242 2289
rect 2792 2256 2822 2289
rect 2792 2255 2822 2256
rect 3372 2255 3402 2289
rect 3952 2256 3982 2289
rect 3952 2255 3982 2256
rect 4532 2255 4562 2289
rect 5112 2256 5142 2289
rect 5112 2255 5142 2256
rect 5692 2255 5722 2289
rect 6272 2256 6302 2289
rect 6272 2255 6302 2256
rect 6852 2255 6882 2289
rect 472 1986 502 2019
rect 472 1985 502 1986
rect 1052 1985 1082 2019
rect 1632 1986 1662 2019
rect 1632 1985 1662 1986
rect 2212 1985 2242 2019
rect 2792 1986 2822 2019
rect 2792 1985 2822 1986
rect 3372 1985 3402 2019
rect 3952 1986 3982 2019
rect 3952 1985 3982 1986
rect 4532 1985 4562 2019
rect 5112 1986 5142 2019
rect 5112 1985 5142 1986
rect 5692 1985 5722 2019
rect 6272 1986 6302 2019
rect 6272 1985 6302 1986
rect 6852 1985 6882 2019
rect 472 1716 502 1749
rect 472 1715 502 1716
rect 1052 1715 1082 1749
rect 1632 1716 1662 1749
rect 1632 1715 1662 1716
rect 2212 1715 2242 1749
rect 2792 1716 2822 1749
rect 2792 1715 2822 1716
rect 3372 1715 3402 1749
rect 3952 1716 3982 1749
rect 3952 1715 3982 1716
rect 4532 1715 4562 1749
rect 5112 1716 5142 1749
rect 5112 1715 5142 1716
rect 5692 1715 5722 1749
rect 6272 1716 6302 1749
rect 6272 1715 6302 1716
rect 6852 1715 6882 1749
rect 472 1446 502 1479
rect 472 1445 502 1446
rect 1052 1445 1082 1479
rect 1632 1446 1662 1479
rect 1632 1445 1662 1446
rect 2212 1445 2242 1479
rect 2792 1446 2822 1479
rect 2792 1445 2822 1446
rect 3372 1445 3402 1479
rect 3952 1446 3982 1479
rect 3952 1445 3982 1446
rect 4532 1445 4562 1479
rect 5112 1446 5142 1479
rect 5112 1445 5142 1446
rect 5692 1445 5722 1479
rect 6272 1446 6302 1479
rect 6272 1445 6302 1446
rect 6852 1445 6882 1479
rect 472 1176 502 1209
rect 472 1175 502 1176
rect 1052 1175 1082 1209
rect 1632 1176 1662 1209
rect 1632 1175 1662 1176
rect 2212 1175 2242 1209
rect 2792 1176 2822 1209
rect 2792 1175 2822 1176
rect 3372 1175 3402 1209
rect 3952 1176 3982 1209
rect 3952 1175 3982 1176
rect 4532 1175 4562 1209
rect 5112 1176 5142 1209
rect 5112 1175 5142 1176
rect 5692 1175 5722 1209
rect 6272 1176 6302 1209
rect 6272 1175 6302 1176
rect 6852 1175 6882 1209
rect 472 906 502 939
rect 472 905 502 906
rect 1052 905 1082 939
rect 1632 906 1662 939
rect 1632 905 1662 906
rect 2212 905 2242 939
rect 2792 906 2822 939
rect 2792 905 2822 906
rect 3372 905 3402 939
rect 3952 906 3982 939
rect 3952 905 3982 906
rect 4532 905 4562 939
rect 5112 906 5142 939
rect 5112 905 5142 906
rect 5692 905 5722 939
rect 6272 906 6302 939
rect 6272 905 6302 906
rect 6852 905 6882 939
rect 472 636 502 669
rect 472 635 502 636
rect 1052 635 1082 669
rect 1632 636 1662 669
rect 1632 635 1662 636
rect 2212 635 2242 669
rect 2792 636 2822 669
rect 2792 635 2822 636
rect 3372 635 3402 669
rect 3952 636 3982 669
rect 3952 635 3982 636
rect 4532 635 4562 669
rect 5112 636 5142 669
rect 5112 635 5142 636
rect 5692 635 5722 669
rect 6272 636 6302 669
rect 6272 635 6302 636
rect 6852 635 6882 669
rect 472 366 502 399
rect 472 365 502 366
rect 1052 365 1082 399
rect 1632 366 1662 399
rect 1632 365 1662 366
rect 2212 365 2242 399
rect 2792 366 2822 399
rect 2792 365 2822 366
rect 3372 365 3402 399
rect 3952 366 3982 399
rect 3952 365 3982 366
rect 4532 365 4562 399
rect 5112 366 5142 399
rect 5112 365 5142 366
rect 5692 365 5722 399
rect 6272 366 6302 399
rect 6272 365 6302 366
rect 6852 365 6882 399
rect 472 96 502 129
rect 472 95 502 96
rect 1052 95 1082 129
rect 1632 96 1662 129
rect 1632 95 1662 96
rect 2212 95 2242 129
rect 2792 96 2822 129
rect 2792 95 2822 96
rect 3372 95 3402 129
rect 3952 96 3982 129
rect 3952 95 3982 96
rect 4532 95 4562 129
rect 5112 96 5142 129
rect 5112 95 5142 96
rect 5692 95 5722 129
rect 6272 96 6302 129
rect 6272 95 6302 96
rect 6852 95 6882 129
<< metal2 >>
rect -91 4145 472 4179
rect 502 4145 1052 4179
rect 1082 4145 1632 4179
rect 1662 4145 2212 4179
rect 2242 4145 2792 4179
rect 2822 4145 3372 4179
rect 3402 4145 3952 4179
rect 3982 4145 4532 4179
rect 4562 4145 5112 4179
rect 5142 4145 5692 4179
rect 5722 4145 6272 4179
rect 6302 4145 6852 4179
rect 6882 4145 6952 4179
rect -91 3875 472 3909
rect 502 3875 1052 3909
rect 1082 3875 1632 3909
rect 1662 3875 2212 3909
rect 2242 3875 2792 3909
rect 2822 3875 3372 3909
rect 3402 3875 3952 3909
rect 3982 3875 4532 3909
rect 4562 3875 5112 3909
rect 5142 3875 5692 3909
rect 5722 3875 6272 3909
rect 6302 3875 6852 3909
rect 6882 3875 6952 3909
rect -91 3605 472 3639
rect 502 3605 1052 3639
rect 1082 3605 1632 3639
rect 1662 3605 2212 3639
rect 2242 3605 2792 3639
rect 2822 3605 3372 3639
rect 3402 3605 3952 3639
rect 3982 3605 4532 3639
rect 4562 3605 5112 3639
rect 5142 3605 5692 3639
rect 5722 3605 6272 3639
rect 6302 3605 6852 3639
rect 6882 3605 6952 3639
rect -91 3335 472 3369
rect 502 3335 1052 3369
rect 1082 3335 1632 3369
rect 1662 3335 2212 3369
rect 2242 3335 2792 3369
rect 2822 3335 3372 3369
rect 3402 3335 3952 3369
rect 3982 3335 4532 3369
rect 4562 3335 5112 3369
rect 5142 3335 5692 3369
rect 5722 3335 6272 3369
rect 6302 3335 6852 3369
rect 6882 3335 6952 3369
rect -91 3065 472 3099
rect 502 3065 1052 3099
rect 1082 3065 1632 3099
rect 1662 3065 2212 3099
rect 2242 3065 2792 3099
rect 2822 3065 3372 3099
rect 3402 3065 3952 3099
rect 3982 3065 4532 3099
rect 4562 3065 5112 3099
rect 5142 3065 5692 3099
rect 5722 3065 6272 3099
rect 6302 3065 6852 3099
rect 6882 3065 6952 3099
rect -91 2795 472 2829
rect 502 2795 1052 2829
rect 1082 2795 1632 2829
rect 1662 2795 2212 2829
rect 2242 2795 2792 2829
rect 2822 2795 3372 2829
rect 3402 2795 3952 2829
rect 3982 2795 4532 2829
rect 4562 2795 5112 2829
rect 5142 2795 5692 2829
rect 5722 2795 6272 2829
rect 6302 2795 6852 2829
rect 6882 2795 6952 2829
rect -91 2525 472 2559
rect 502 2525 1052 2559
rect 1082 2525 1632 2559
rect 1662 2525 2212 2559
rect 2242 2525 2792 2559
rect 2822 2525 3372 2559
rect 3402 2525 3952 2559
rect 3982 2525 4532 2559
rect 4562 2525 5112 2559
rect 5142 2525 5692 2559
rect 5722 2525 6272 2559
rect 6302 2525 6852 2559
rect 6882 2525 6952 2559
rect -91 2255 472 2289
rect 502 2255 1052 2289
rect 1082 2255 1632 2289
rect 1662 2255 2212 2289
rect 2242 2255 2792 2289
rect 2822 2255 3372 2289
rect 3402 2255 3952 2289
rect 3982 2255 4532 2289
rect 4562 2255 5112 2289
rect 5142 2255 5692 2289
rect 5722 2255 6272 2289
rect 6302 2255 6852 2289
rect 6882 2255 6952 2289
rect -91 1985 472 2019
rect 502 1985 1052 2019
rect 1082 1985 1632 2019
rect 1662 1985 2212 2019
rect 2242 1985 2792 2019
rect 2822 1985 3372 2019
rect 3402 1985 3952 2019
rect 3982 1985 4532 2019
rect 4562 1985 5112 2019
rect 5142 1985 5692 2019
rect 5722 1985 6272 2019
rect 6302 1985 6852 2019
rect 6882 1985 6952 2019
rect -91 1715 472 1749
rect 502 1715 1052 1749
rect 1082 1715 1632 1749
rect 1662 1715 2212 1749
rect 2242 1715 2792 1749
rect 2822 1715 3372 1749
rect 3402 1715 3952 1749
rect 3982 1715 4532 1749
rect 4562 1715 5112 1749
rect 5142 1715 5692 1749
rect 5722 1715 6272 1749
rect 6302 1715 6852 1749
rect 6882 1715 6952 1749
rect -91 1445 472 1479
rect 502 1445 1052 1479
rect 1082 1445 1632 1479
rect 1662 1445 2212 1479
rect 2242 1445 2792 1479
rect 2822 1445 3372 1479
rect 3402 1445 3952 1479
rect 3982 1445 4532 1479
rect 4562 1445 5112 1479
rect 5142 1445 5692 1479
rect 5722 1445 6272 1479
rect 6302 1445 6852 1479
rect 6882 1445 6952 1479
rect -91 1175 472 1209
rect 502 1175 1052 1209
rect 1082 1175 1632 1209
rect 1662 1175 2212 1209
rect 2242 1175 2792 1209
rect 2822 1175 3372 1209
rect 3402 1175 3952 1209
rect 3982 1175 4532 1209
rect 4562 1175 5112 1209
rect 5142 1175 5692 1209
rect 5722 1175 6272 1209
rect 6302 1175 6852 1209
rect 6882 1175 6952 1209
rect -91 905 472 939
rect 502 905 1052 939
rect 1082 905 1632 939
rect 1662 905 2212 939
rect 2242 905 2792 939
rect 2822 905 3372 939
rect 3402 905 3952 939
rect 3982 905 4532 939
rect 4562 905 5112 939
rect 5142 905 5692 939
rect 5722 905 6272 939
rect 6302 905 6852 939
rect 6882 905 6952 939
rect -91 635 472 669
rect 502 635 1052 669
rect 1082 635 1632 669
rect 1662 635 2212 669
rect 2242 635 2792 669
rect 2822 635 3372 669
rect 3402 635 3952 669
rect 3982 635 4532 669
rect 4562 635 5112 669
rect 5142 635 5692 669
rect 5722 635 6272 669
rect 6302 635 6852 669
rect 6882 635 6952 669
rect -91 365 472 399
rect 502 365 1052 399
rect 1082 365 1632 399
rect 1662 365 2212 399
rect 2242 365 2792 399
rect 2822 365 3372 399
rect 3402 365 3952 399
rect 3982 365 4532 399
rect 4562 365 5112 399
rect 5142 365 5692 399
rect 5722 365 6272 399
rect 6302 365 6852 399
rect 6882 365 6952 399
rect -91 95 472 129
rect 502 95 1052 129
rect 1082 95 1632 129
rect 1662 95 2212 129
rect 2242 95 2792 129
rect 2822 95 3372 129
rect 3402 95 3952 129
rect 3982 95 4532 129
rect 4562 95 5112 129
rect 5142 95 5692 129
rect 5722 95 6272 129
rect 6302 95 6852 129
rect 6882 95 6952 129
<< labels >>
rlabel corelocali 530 -55 545 -7 1 RBL0_0
port 6 ns signal output
rlabel corelocali -7 -55 8 -7 1 RBL1_0
port 7 ns signal output
rlabel corelocali 429 -55 444 -7 1 WBL_0
port 8 ns signal input
rlabel corelocali 94 -55 109 -7 1 WBLb_0
port 9 ns signal input
rlabel corelocali 1110 -55 1125 -7 1 RBL0_1
port 55 ns signal output
rlabel corelocali 573 -55 588 -7 1 RBL1_1
port 56 ns signal output
rlabel corelocali 1009 -55 1024 -7 1 WBL_1
port 57 ns signal input
rlabel corelocali 674 -55 689 -7 1 WBLb_1
port 58 ns signal input
rlabel corelocali 1690 -55 1705 -7 1 RBL0_2
port 59 ns signal output
rlabel corelocali 1153 -55 1168 -7 1 RBL1_2
port 60 ns signal output
rlabel corelocali 1589 -55 1604 -7 1 WBL_2
port 61 ns signal input
rlabel corelocali 1254 -55 1269 -7 1 WBLb_2
port 62 ns signal input
rlabel corelocali 2270 -55 2285 -7 1 RBL0_3
port 63 ns signal output
rlabel corelocali 1733 -55 1748 -7 1 RBL1_3
port 64 ns signal output
rlabel corelocali 2169 -55 2184 -7 1 WBL_3
port 65 ns signal input
rlabel corelocali 1834 -55 1849 -7 1 WBLb_3
port 66 ns signal input
rlabel corelocali 2850 -55 2865 -7 1 RBL0_4
port 67 ns signal output
rlabel corelocali 2313 -55 2328 -7 1 RBL1_4
port 68 ns signal output
rlabel corelocali 2749 -55 2764 -7 1 WBL_4
port 69 ns signal input
rlabel corelocali 2414 -55 2429 -7 1 WBLb_4
port 70 ns signal input
rlabel corelocali 3430 -55 3445 -7 1 RBL0_5
port 71 ns signal output
rlabel corelocali 2893 -55 2908 -7 1 RBL1_5
port 72 ns signal output
rlabel corelocali 3329 -55 3344 -7 1 WBL_5
port 73 ns signal input
rlabel corelocali 2994 -55 3009 -7 1 WBLb_5
port 74 ns signal input
rlabel corelocali 4010 -55 4025 -7 1 RBL0_6
port 75 ns signal output
rlabel corelocali 3473 -55 3488 -7 1 RBL1_6
port 76 ns signal output
rlabel corelocali 3909 -55 3924 -7 1 WBL_6
port 77 ns signal input
rlabel corelocali 3574 -55 3589 -7 1 WBLb_6
port 78 ns signal input
rlabel corelocali 4590 -55 4605 -7 1 RBL0_7
port 79 ns signal output
rlabel corelocali 4053 -55 4068 -7 1 RBL1_7
port 80 ns signal output
rlabel corelocali 4489 -55 4504 -7 1 WBL_7
port 81 ns signal input
rlabel corelocali 4154 -55 4169 -7 1 WBLb_7
port 82 ns signal input
rlabel corelocali 5170 -55 5185 -7 1 RBL0_8
port 83 ns signal output
rlabel corelocali 4633 -55 4648 -7 1 RBL1_8
port 84 ns signal output
rlabel corelocali 5069 -55 5084 -7 1 WBL_8
port 85 ns signal input
rlabel corelocali 4734 -55 4749 -7 1 WBLb_8
port 86 ns signal input
rlabel corelocali 5750 -55 5765 -7 1 RBL0_9
port 87 ns signal output
rlabel corelocali 5213 -55 5228 -7 1 RBL1_9
port 88 ns signal output
rlabel corelocali 5649 -55 5664 -7 1 WBL_9
port 89 ns signal input
rlabel corelocali 5314 -55 5329 -7 1 WBLb_9
port 90 ns signal input
rlabel corelocali 6330 -55 6345 -7 1 RBL0_10
port 91 ns signal output
rlabel corelocali 5793 -55 5808 -7 1 RBL1_10
port 92 ns signal output
rlabel corelocali 6229 -55 6244 -7 1 WBL_10
port 93 ns signal input
rlabel corelocali 5894 -55 5909 -7 1 WBLb_10
port 94 ns signal input
rlabel corelocali 6910 -55 6925 -7 1 RBL0_11
port 95 ns signal output
rlabel corelocali 6373 -55 6388 -7 1 RBL1_11
port 96 ns signal output
rlabel corelocali 6809 -55 6824 -7 1 WBL_11
port 97 ns signal input
rlabel corelocali 6474 -55 6489 -7 1 WBLb_11
port 98 ns signal input
rlabel metal1 -91 219 -43 233 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 -7 -43 7 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 489 -43 503 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 263 -43 277 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 759 -43 773 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 533 -43 547 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 1029 -43 1043 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 803 -43 817 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 1299 -43 1313 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 1073 -43 1087 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 1569 -43 1583 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 1343 -43 1357 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 1839 -43 1853 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 1613 -43 1627 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 2109 -43 2123 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 1883 -43 1897 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 2379 -43 2393 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 2153 -43 2167 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 2649 -43 2663 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 2423 -43 2437 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 2919 -43 2933 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 2693 -43 2707 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 3189 -43 3203 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 2963 -43 2977 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 3459 -43 3473 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 3233 -43 3247 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 3729 -43 3743 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 3503 -43 3517 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 3999 -43 4013 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 3773 -43 3787 1 GND
port 2 ew ground bidirectional abutment
rlabel metal1 -91 4269 -43 4283 1 VDD
port 1 ew power bidirectional abutment
rlabel metal1 -91 4043 -43 4057 1 GND
port 2 ew ground bidirectional abutment
rlabel polycont -91 233 -43 263 1 WWL_0
port 3 ew signal input
rlabel metal2 -91 95 -67 129 1 RWL0_0
port 4 ew signal input
rlabel metal1 -67 95 -43 129 1 RWL1_0
port 5 ew signal input
rlabel polycont -91 503 -43 533 1 WWL_1
port 10 ew signal input
rlabel metal2 -91 365 -67 399 1 RWL0_1
port 11 ew signal input
rlabel metal1 -67 365 -43 399 1 RWL1_1
port 12 ew signal input
rlabel polycont -91 773 -43 803 1 WWL_2
port 13 ew signal input
rlabel metal2 -91 635 -67 669 1 RWL0_2
port 14 ew signal input
rlabel metal1 -67 635 -43 669 1 RWL1_2
port 15 ew signal input
rlabel polycont -91 1043 -43 1073 1 WWL_3
port 16 ew signal input
rlabel metal2 -91 905 -67 939 1 RWL0_3
port 17 ew signal input
rlabel metal1 -67 905 -43 939 1 RWL1_3
port 18 ew signal input
rlabel polycont -91 1313 -43 1343 1 WWL_4
port 19 ew signal input
rlabel metal2 -91 1175 -67 1209 1 RWL0_4
port 20 ew signal input
rlabel metal1 -67 1175 -43 1209 1 RWL1_4
port 21 ew signal input
rlabel polycont -91 1583 -43 1613 1 WWL_5
port 22 ew signal input
rlabel metal2 -91 1445 -67 1479 1 RWL0_5
port 23 ew signal input
rlabel metal1 -67 1445 -43 1479 1 RWL1_5
port 24 ew signal input
rlabel polycont -91 1853 -43 1883 1 WWL_6
port 25 ew signal input
rlabel metal2 -91 1715 -67 1749 1 RWL0_6
port 26 ew signal input
rlabel metal1 -67 1715 -43 1749 1 RWL1_6
port 27 ew signal input
rlabel polycont -91 2123 -43 2153 1 WWL_7
port 28 ew signal input
rlabel metal2 -91 1985 -67 2019 1 RWL0_7
port 29 ew signal input
rlabel metal1 -67 1985 -43 2019 1 RWL1_7
port 30 ew signal input
rlabel polycont -91 2393 -43 2423 1 WWL_8
port 31 ew signal input
rlabel metal2 -91 2255 -67 2289 1 RWL0_8
port 32 ew signal input
rlabel metal1 -67 2255 -43 2289 1 RWL1_8
port 33 ew signal input
rlabel polycont -91 2663 -43 2693 1 WWL_9
port 34 ew signal input
rlabel metal2 -91 2525 -67 2559 1 RWL0_9
port 35 ew signal input
rlabel metal1 -67 2525 -43 2559 1 RWL1_9
port 36 ew signal input
rlabel polycont -91 2933 -43 2963 1 WWL_10
port 37 ew signal input
rlabel metal2 -91 2795 -67 2829 1 RWL0_10
port 38 ew signal input
rlabel metal1 -67 2795 -43 2829 1 RWL1_10
port 39 ew signal input
rlabel polycont -91 3203 -43 3233 1 WWL_11
port 40 ew signal input
rlabel metal2 -91 3065 -67 3099 1 RWL0_11
port 41 ew signal input
rlabel metal1 -67 3065 -43 3099 1 RWL1_11
port 42 ew signal input
rlabel polycont -91 3473 -43 3503 1 WWL_12
port 43 ew signal input
rlabel metal2 -91 3335 -67 3369 1 RWL0_12
port 44 ew signal input
rlabel metal1 -67 3335 -43 3369 1 RWL1_12
port 45 ew signal input
rlabel polycont -91 3743 -43 3773 1 WWL_13
port 46 ew signal input
rlabel metal2 -91 3605 -67 3639 1 RWL0_13
port 47 ew signal input
rlabel metal1 -67 3605 -43 3639 1 RWL1_13
port 48 ew signal input
rlabel polycont -91 4013 -43 4043 1 WWL_14
port 49 ew signal input
rlabel metal2 -91 3875 -67 3909 1 RWL0_14
port 50 ew signal input
rlabel metal1 -67 3875 -43 3909 1 RWL1_14
port 51 ew signal input
rlabel polycont -91 4283 -43 4313 1 WWL_15
port 52 ew signal input
rlabel metal2 -91 4145 -67 4179 1 RWL0_15
port 53 ew signal input
rlabel metal1 -67 4145 -43 4179 1 RWL1_15
port 54 ew signal input
<< end >>
