magic
tech sky130A
magscale 1 2
timestamp 1668118531
<< error_p >>
rect 14 2158 27 2174
rect 116 2172 129 2174
rect 82 2158 97 2172
rect 106 2158 136 2172
rect 197 2170 350 2216
rect 179 2158 371 2170
rect 414 2158 444 2172
rect 450 2158 463 2174
rect 551 2158 564 2174
rect 594 2158 607 2174
rect 696 2172 709 2174
rect 662 2158 677 2172
rect 686 2158 716 2172
rect 777 2170 930 2216
rect 759 2158 951 2170
rect 994 2158 1024 2172
rect 1030 2158 1043 2174
rect 1131 2158 1144 2174
rect 1174 2158 1187 2174
rect 1276 2172 1289 2174
rect 1242 2158 1257 2172
rect 1266 2158 1296 2172
rect 1357 2170 1510 2216
rect 1339 2158 1531 2170
rect 1574 2158 1604 2172
rect 1610 2158 1623 2174
rect 1711 2158 1724 2174
rect 1754 2158 1767 2174
rect 1822 2158 1837 2172
rect 3494 2158 3507 2174
rect 3596 2172 3609 2174
rect 3562 2158 3577 2172
rect 3586 2158 3616 2172
rect 3677 2170 3830 2216
rect 3659 2158 3851 2170
rect 3894 2158 3924 2172
rect 3930 2158 3943 2174
rect 4031 2158 4044 2174
rect 4074 2158 4087 2174
rect 4176 2172 4189 2174
rect 4142 2158 4157 2172
rect 4166 2158 4196 2172
rect 4257 2170 4410 2216
rect 4239 2158 4431 2170
rect 4474 2158 4504 2172
rect 4510 2158 4523 2174
rect 4611 2158 4624 2174
rect 4654 2158 4667 2174
rect 4756 2172 4769 2174
rect 4722 2158 4737 2172
rect 4746 2158 4776 2172
rect 4837 2170 4990 2216
rect 4819 2158 5011 2170
rect 5054 2158 5084 2172
rect 5090 2158 5103 2174
rect 5191 2158 5204 2174
rect 5234 2158 5247 2174
rect 5336 2172 5349 2174
rect 5302 2158 5317 2172
rect 5326 2158 5356 2172
rect 5417 2170 5570 2216
rect 5399 2158 5591 2170
rect 5634 2158 5664 2172
rect 5670 2158 5683 2174
rect 5771 2158 5784 2174
rect 5814 2158 5827 2174
rect 5916 2172 5929 2174
rect 5882 2158 5897 2172
rect 5906 2158 5936 2172
rect 5997 2170 6150 2216
rect 5979 2158 6171 2170
rect 6214 2158 6244 2172
rect 6250 2158 6263 2174
rect 6351 2158 6364 2174
rect 6394 2158 6407 2174
rect 6496 2172 6509 2174
rect 6462 2158 6477 2172
rect 6486 2158 6516 2172
rect 6577 2170 6730 2216
rect 6559 2158 6751 2170
rect 6794 2158 6824 2172
rect 6830 2158 6843 2174
rect 6931 2158 6944 2174
rect -1 2144 1837 2158
rect 3481 2144 6944 2158
rect 14 2040 27 2144
rect 72 2122 73 2132
rect 88 2122 101 2132
rect 72 2118 101 2122
rect 106 2118 136 2144
rect 154 2130 170 2132
rect 242 2130 295 2144
rect 243 2128 307 2130
rect 350 2128 365 2144
rect 414 2141 444 2144
rect 414 2138 450 2141
rect 380 2130 396 2132
rect 154 2118 169 2122
rect 72 2116 169 2118
rect 197 2116 365 2128
rect 381 2118 396 2122
rect 414 2119 453 2138
rect 472 2132 479 2133
rect 478 2125 479 2132
rect 462 2122 463 2125
rect 478 2122 491 2125
rect 414 2118 444 2119
rect 453 2118 459 2119
rect 462 2118 491 2122
rect 381 2117 491 2118
rect 381 2116 497 2117
rect 56 2108 107 2116
rect 56 2096 81 2108
rect 88 2096 107 2108
rect 138 2108 188 2116
rect 138 2100 154 2108
rect 161 2106 188 2108
rect 197 2106 418 2116
rect 161 2096 418 2106
rect 447 2108 497 2116
rect 447 2099 463 2108
rect 56 2088 107 2096
rect 154 2088 418 2096
rect 444 2096 463 2099
rect 470 2096 497 2108
rect 444 2088 497 2096
rect 72 2080 73 2088
rect 88 2080 101 2088
rect 72 2072 88 2080
rect 69 2065 88 2068
rect 69 2056 91 2065
rect 42 2046 91 2056
rect 42 2040 72 2046
rect 91 2041 96 2046
rect 14 2024 88 2040
rect 106 2032 136 2088
rect 171 2078 379 2088
rect 414 2084 459 2088
rect 462 2087 463 2088
rect 478 2087 491 2088
rect 197 2048 386 2078
rect 212 2045 386 2048
rect 205 2042 386 2045
rect 14 2022 27 2024
rect 42 2022 76 2024
rect 14 2006 88 2022
rect 115 2018 128 2032
rect 143 2018 159 2034
rect 205 2029 216 2042
rect -2 1984 -1 2000
rect 14 1984 27 2006
rect 42 1984 72 2006
rect 115 2002 177 2018
rect 205 2011 216 2027
rect 221 2022 231 2042
rect 241 2022 255 2042
rect 258 2029 267 2042
rect 283 2029 292 2042
rect 221 2011 255 2022
rect 258 2011 267 2027
rect 283 2011 292 2027
rect 299 2022 309 2042
rect 319 2022 333 2042
rect 334 2029 345 2042
rect 299 2011 333 2022
rect 334 2011 345 2027
rect 391 2018 407 2034
rect 414 2032 444 2084
rect 478 2080 479 2087
rect 463 2072 479 2080
rect 450 2040 463 2059
rect 478 2040 508 2056
rect 450 2024 524 2040
rect 450 2022 463 2024
rect 478 2022 512 2024
rect 115 2000 128 2002
rect 143 2000 177 2002
rect 115 1984 177 2000
rect 221 1995 237 2002
rect 299 1995 329 2006
rect 377 2002 423 2018
rect 450 2006 524 2022
rect 377 2000 411 2002
rect 376 1984 423 2000
rect 450 1984 463 2006
rect 478 1984 508 2006
rect 535 1984 536 2000
rect 551 1984 564 2144
rect 594 2040 607 2144
rect 652 2122 653 2132
rect 668 2122 681 2132
rect 652 2118 681 2122
rect 686 2118 716 2144
rect 734 2130 750 2132
rect 822 2130 875 2144
rect 823 2128 887 2130
rect 930 2128 945 2144
rect 994 2141 1024 2144
rect 994 2138 1030 2141
rect 960 2130 976 2132
rect 734 2118 749 2122
rect 652 2116 749 2118
rect 777 2116 945 2128
rect 961 2118 976 2122
rect 994 2119 1033 2138
rect 1052 2132 1059 2133
rect 1058 2125 1059 2132
rect 1042 2122 1043 2125
rect 1058 2122 1071 2125
rect 994 2118 1024 2119
rect 1033 2118 1039 2119
rect 1042 2118 1071 2122
rect 961 2117 1071 2118
rect 961 2116 1077 2117
rect 636 2108 687 2116
rect 636 2096 661 2108
rect 668 2096 687 2108
rect 718 2108 768 2116
rect 718 2100 734 2108
rect 741 2106 768 2108
rect 777 2106 998 2116
rect 741 2096 998 2106
rect 1027 2108 1077 2116
rect 1027 2099 1043 2108
rect 636 2088 687 2096
rect 734 2088 998 2096
rect 1024 2096 1043 2099
rect 1050 2096 1077 2108
rect 1024 2088 1077 2096
rect 652 2080 653 2088
rect 668 2080 681 2088
rect 652 2072 668 2080
rect 649 2065 668 2068
rect 649 2056 671 2065
rect 622 2046 671 2056
rect 622 2040 652 2046
rect 671 2041 676 2046
rect 594 2024 668 2040
rect 686 2032 716 2088
rect 751 2078 959 2088
rect 994 2084 1039 2088
rect 1042 2087 1043 2088
rect 1058 2087 1071 2088
rect 777 2048 966 2078
rect 792 2045 966 2048
rect 785 2042 966 2045
rect 594 2022 607 2024
rect 622 2022 656 2024
rect 594 2006 668 2022
rect 695 2018 708 2032
rect 723 2018 739 2034
rect 785 2029 796 2042
rect 578 1984 579 2000
rect 594 1984 607 2006
rect 622 1984 652 2006
rect 695 2002 757 2018
rect 785 2011 796 2027
rect 801 2022 811 2042
rect 821 2022 835 2042
rect 838 2029 847 2042
rect 863 2029 872 2042
rect 801 2011 835 2022
rect 838 2011 847 2027
rect 863 2011 872 2027
rect 879 2022 889 2042
rect 899 2022 913 2042
rect 914 2029 925 2042
rect 879 2011 913 2022
rect 914 2011 925 2027
rect 971 2018 987 2034
rect 994 2032 1024 2084
rect 1058 2080 1059 2087
rect 1043 2072 1059 2080
rect 1030 2040 1043 2059
rect 1058 2040 1088 2056
rect 1030 2024 1104 2040
rect 1030 2022 1043 2024
rect 1058 2022 1092 2024
rect 695 2000 708 2002
rect 723 2000 757 2002
rect 695 1984 757 2000
rect 801 1995 817 2002
rect 879 1995 909 2006
rect 957 2002 1003 2018
rect 1030 2006 1104 2022
rect 957 2000 991 2002
rect 956 1984 1003 2000
rect 1030 1984 1043 2006
rect 1058 1984 1088 2006
rect 1115 1984 1116 2000
rect 1131 1984 1144 2144
rect 1174 2040 1187 2144
rect 1232 2122 1233 2132
rect 1248 2122 1261 2132
rect 1232 2118 1261 2122
rect 1266 2118 1296 2144
rect 1314 2130 1330 2132
rect 1402 2130 1455 2144
rect 1403 2128 1467 2130
rect 1510 2128 1525 2144
rect 1574 2141 1604 2144
rect 1574 2138 1610 2141
rect 1540 2130 1556 2132
rect 1314 2118 1329 2122
rect 1232 2116 1329 2118
rect 1357 2116 1525 2128
rect 1541 2118 1556 2122
rect 1574 2119 1613 2138
rect 1632 2132 1639 2133
rect 1638 2125 1639 2132
rect 1622 2122 1623 2125
rect 1638 2122 1651 2125
rect 1574 2118 1604 2119
rect 1613 2118 1619 2119
rect 1622 2118 1651 2122
rect 1541 2117 1651 2118
rect 1541 2116 1657 2117
rect 1216 2108 1267 2116
rect 1216 2096 1241 2108
rect 1248 2096 1267 2108
rect 1298 2108 1348 2116
rect 1298 2100 1314 2108
rect 1321 2106 1348 2108
rect 1357 2106 1578 2116
rect 1321 2096 1578 2106
rect 1607 2108 1657 2116
rect 1607 2099 1623 2108
rect 1216 2088 1267 2096
rect 1314 2088 1578 2096
rect 1604 2096 1623 2099
rect 1630 2096 1657 2108
rect 1604 2088 1657 2096
rect 1232 2080 1233 2088
rect 1248 2080 1261 2088
rect 1232 2072 1248 2080
rect 1229 2065 1248 2068
rect 1229 2056 1251 2065
rect 1202 2046 1251 2056
rect 1202 2040 1232 2046
rect 1251 2041 1256 2046
rect 1174 2024 1248 2040
rect 1266 2032 1296 2088
rect 1331 2078 1539 2088
rect 1574 2084 1619 2088
rect 1622 2087 1623 2088
rect 1638 2087 1651 2088
rect 1357 2048 1546 2078
rect 1372 2045 1546 2048
rect 1365 2042 1546 2045
rect 1174 2022 1187 2024
rect 1202 2022 1236 2024
rect 1174 2006 1248 2022
rect 1275 2018 1288 2032
rect 1303 2018 1319 2034
rect 1365 2029 1376 2042
rect 1158 1984 1159 2000
rect 1174 1984 1187 2006
rect 1202 1984 1232 2006
rect 1275 2002 1337 2018
rect 1365 2011 1376 2027
rect 1381 2022 1391 2042
rect 1401 2022 1415 2042
rect 1418 2029 1427 2042
rect 1443 2029 1452 2042
rect 1381 2011 1415 2022
rect 1418 2011 1427 2027
rect 1443 2011 1452 2027
rect 1459 2022 1469 2042
rect 1479 2022 1493 2042
rect 1494 2029 1505 2042
rect 1459 2011 1493 2022
rect 1494 2011 1505 2027
rect 1551 2018 1567 2034
rect 1574 2032 1604 2084
rect 1638 2080 1639 2087
rect 1623 2072 1639 2080
rect 1610 2040 1623 2059
rect 1638 2040 1668 2056
rect 1610 2024 1684 2040
rect 1610 2022 1623 2024
rect 1638 2022 1672 2024
rect 1275 2000 1288 2002
rect 1303 2000 1337 2002
rect 1275 1984 1337 2000
rect 1381 1995 1397 2002
rect 1459 1995 1489 2006
rect 1537 2002 1583 2018
rect 1610 2006 1684 2022
rect 1537 2000 1571 2002
rect 1536 1984 1583 2000
rect 1610 1984 1623 2006
rect 1638 1984 1668 2006
rect 1695 1984 1696 2000
rect 1711 1984 1724 2144
rect 1754 2040 1767 2144
rect 1812 2122 1813 2132
rect 1828 2122 1837 2132
rect 1812 2116 1837 2122
rect 1796 2108 1837 2116
rect 1796 2096 1821 2108
rect 1828 2096 1837 2108
rect 1796 2088 1837 2096
rect 1812 2080 1813 2088
rect 1828 2080 1837 2088
rect 1812 2072 1828 2080
rect 1809 2065 1828 2068
rect 1809 2056 1831 2065
rect 1782 2046 1831 2056
rect 1782 2040 1812 2046
rect 1831 2041 1836 2046
rect 3494 2040 3507 2144
rect 3552 2122 3553 2132
rect 3568 2122 3581 2132
rect 3552 2118 3581 2122
rect 3586 2118 3616 2144
rect 3634 2130 3650 2132
rect 3722 2130 3775 2144
rect 3723 2128 3787 2130
rect 3830 2128 3845 2144
rect 3894 2141 3924 2144
rect 3894 2138 3930 2141
rect 3860 2130 3876 2132
rect 3634 2118 3649 2122
rect 3552 2116 3649 2118
rect 3677 2116 3845 2128
rect 3861 2118 3876 2122
rect 3894 2119 3933 2138
rect 3952 2132 3959 2133
rect 3958 2125 3959 2132
rect 3942 2122 3943 2125
rect 3958 2122 3971 2125
rect 3894 2118 3924 2119
rect 3933 2118 3939 2119
rect 3942 2118 3971 2122
rect 3861 2117 3971 2118
rect 3861 2116 3977 2117
rect 3536 2108 3587 2116
rect 3536 2096 3561 2108
rect 3568 2096 3587 2108
rect 3618 2108 3668 2116
rect 3618 2100 3634 2108
rect 3641 2106 3668 2108
rect 3677 2106 3898 2116
rect 3641 2096 3898 2106
rect 3927 2108 3977 2116
rect 3927 2099 3943 2108
rect 3536 2088 3587 2096
rect 3634 2088 3898 2096
rect 3924 2096 3943 2099
rect 3950 2096 3977 2108
rect 3924 2088 3977 2096
rect 3552 2080 3553 2088
rect 3568 2080 3581 2088
rect 3552 2072 3568 2080
rect 3549 2065 3568 2068
rect 3549 2056 3571 2065
rect 3522 2046 3571 2056
rect 3522 2040 3552 2046
rect 3571 2041 3576 2046
rect 1754 2024 1828 2040
rect 3494 2024 3568 2040
rect 3586 2032 3616 2088
rect 3651 2078 3859 2088
rect 3894 2084 3939 2088
rect 3942 2087 3943 2088
rect 3958 2087 3971 2088
rect 3677 2048 3866 2078
rect 3692 2045 3866 2048
rect 3685 2042 3866 2045
rect 1754 2022 1767 2024
rect 1782 2022 1816 2024
rect 3494 2022 3507 2024
rect 3522 2022 3556 2024
rect 1754 2006 1828 2022
rect 3494 2006 3568 2022
rect 3595 2018 3608 2032
rect 3623 2018 3639 2034
rect 3685 2029 3696 2042
rect 1738 1984 1739 2000
rect 1754 1984 1767 2006
rect 1782 1984 1812 2006
rect 3494 1984 3507 2006
rect 3522 1984 3552 2006
rect 3595 2002 3657 2018
rect 3685 2011 3696 2027
rect 3701 2022 3711 2042
rect 3721 2022 3735 2042
rect 3738 2029 3747 2042
rect 3763 2029 3772 2042
rect 3701 2011 3735 2022
rect 3738 2011 3747 2027
rect 3763 2011 3772 2027
rect 3779 2022 3789 2042
rect 3799 2022 3813 2042
rect 3814 2029 3825 2042
rect 3779 2011 3813 2022
rect 3814 2011 3825 2027
rect 3871 2018 3887 2034
rect 3894 2032 3924 2084
rect 3958 2080 3959 2087
rect 3943 2072 3959 2080
rect 3930 2040 3943 2059
rect 3958 2040 3988 2056
rect 3930 2024 4004 2040
rect 3930 2022 3943 2024
rect 3958 2022 3992 2024
rect 3595 2000 3608 2002
rect 3623 2000 3657 2002
rect 3595 1984 3657 2000
rect 3701 1995 3717 2002
rect 3779 1995 3809 2006
rect 3857 2002 3903 2018
rect 3930 2006 4004 2022
rect 3857 2000 3891 2002
rect 3856 1984 3903 2000
rect 3930 1984 3943 2006
rect 3958 1984 3988 2006
rect 4015 1984 4016 2000
rect 4031 1984 4044 2144
rect 4074 2040 4087 2144
rect 4132 2122 4133 2132
rect 4148 2122 4161 2132
rect 4132 2118 4161 2122
rect 4166 2118 4196 2144
rect 4214 2130 4230 2132
rect 4302 2130 4355 2144
rect 4303 2128 4367 2130
rect 4410 2128 4425 2144
rect 4474 2141 4504 2144
rect 4474 2138 4510 2141
rect 4440 2130 4456 2132
rect 4214 2118 4229 2122
rect 4132 2116 4229 2118
rect 4257 2116 4425 2128
rect 4441 2118 4456 2122
rect 4474 2119 4513 2138
rect 4532 2132 4539 2133
rect 4538 2125 4539 2132
rect 4522 2122 4523 2125
rect 4538 2122 4551 2125
rect 4474 2118 4504 2119
rect 4513 2118 4519 2119
rect 4522 2118 4551 2122
rect 4441 2117 4551 2118
rect 4441 2116 4557 2117
rect 4116 2108 4167 2116
rect 4116 2096 4141 2108
rect 4148 2096 4167 2108
rect 4198 2108 4248 2116
rect 4198 2100 4214 2108
rect 4221 2106 4248 2108
rect 4257 2106 4478 2116
rect 4221 2096 4478 2106
rect 4507 2108 4557 2116
rect 4507 2099 4523 2108
rect 4116 2088 4167 2096
rect 4214 2088 4478 2096
rect 4504 2096 4523 2099
rect 4530 2096 4557 2108
rect 4504 2088 4557 2096
rect 4132 2080 4133 2088
rect 4148 2080 4161 2088
rect 4132 2072 4148 2080
rect 4129 2065 4148 2068
rect 4129 2056 4151 2065
rect 4102 2046 4151 2056
rect 4102 2040 4132 2046
rect 4151 2041 4156 2046
rect 4074 2024 4148 2040
rect 4166 2032 4196 2088
rect 4231 2078 4439 2088
rect 4474 2084 4519 2088
rect 4522 2087 4523 2088
rect 4538 2087 4551 2088
rect 4257 2048 4446 2078
rect 4272 2045 4446 2048
rect 4265 2042 4446 2045
rect 4074 2022 4087 2024
rect 4102 2022 4136 2024
rect 4074 2006 4148 2022
rect 4175 2018 4188 2032
rect 4203 2018 4219 2034
rect 4265 2029 4276 2042
rect 4058 1984 4059 2000
rect 4074 1984 4087 2006
rect 4102 1984 4132 2006
rect 4175 2002 4237 2018
rect 4265 2011 4276 2027
rect 4281 2022 4291 2042
rect 4301 2022 4315 2042
rect 4318 2029 4327 2042
rect 4343 2029 4352 2042
rect 4281 2011 4315 2022
rect 4318 2011 4327 2027
rect 4343 2011 4352 2027
rect 4359 2022 4369 2042
rect 4379 2022 4393 2042
rect 4394 2029 4405 2042
rect 4359 2011 4393 2022
rect 4394 2011 4405 2027
rect 4451 2018 4467 2034
rect 4474 2032 4504 2084
rect 4538 2080 4539 2087
rect 4523 2072 4539 2080
rect 4510 2040 4523 2059
rect 4538 2040 4568 2056
rect 4510 2024 4584 2040
rect 4510 2022 4523 2024
rect 4538 2022 4572 2024
rect 4175 2000 4188 2002
rect 4203 2000 4237 2002
rect 4175 1984 4237 2000
rect 4281 1995 4297 2002
rect 4359 1995 4389 2006
rect 4437 2002 4483 2018
rect 4510 2006 4584 2022
rect 4437 2000 4471 2002
rect 4436 1984 4483 2000
rect 4510 1984 4523 2006
rect 4538 1984 4568 2006
rect 4595 1984 4596 2000
rect 4611 1984 4624 2144
rect 4654 2040 4667 2144
rect 4712 2122 4713 2132
rect 4728 2122 4741 2132
rect 4712 2118 4741 2122
rect 4746 2118 4776 2144
rect 4794 2130 4810 2132
rect 4882 2130 4935 2144
rect 4883 2128 4947 2130
rect 4990 2128 5005 2144
rect 5054 2141 5084 2144
rect 5054 2138 5090 2141
rect 5020 2130 5036 2132
rect 4794 2118 4809 2122
rect 4712 2116 4809 2118
rect 4837 2116 5005 2128
rect 5021 2118 5036 2122
rect 5054 2119 5093 2138
rect 5112 2132 5119 2133
rect 5118 2125 5119 2132
rect 5102 2122 5103 2125
rect 5118 2122 5131 2125
rect 5054 2118 5084 2119
rect 5093 2118 5099 2119
rect 5102 2118 5131 2122
rect 5021 2117 5131 2118
rect 5021 2116 5137 2117
rect 4696 2108 4747 2116
rect 4696 2096 4721 2108
rect 4728 2096 4747 2108
rect 4778 2108 4828 2116
rect 4778 2100 4794 2108
rect 4801 2106 4828 2108
rect 4837 2106 5058 2116
rect 4801 2096 5058 2106
rect 5087 2108 5137 2116
rect 5087 2099 5103 2108
rect 4696 2088 4747 2096
rect 4794 2088 5058 2096
rect 5084 2096 5103 2099
rect 5110 2096 5137 2108
rect 5084 2088 5137 2096
rect 4712 2080 4713 2088
rect 4728 2080 4741 2088
rect 4712 2072 4728 2080
rect 4709 2065 4728 2068
rect 4709 2056 4731 2065
rect 4682 2046 4731 2056
rect 4682 2040 4712 2046
rect 4731 2041 4736 2046
rect 4654 2024 4728 2040
rect 4746 2032 4776 2088
rect 4811 2078 5019 2088
rect 5054 2084 5099 2088
rect 5102 2087 5103 2088
rect 5118 2087 5131 2088
rect 4837 2048 5026 2078
rect 4852 2045 5026 2048
rect 4845 2042 5026 2045
rect 4654 2022 4667 2024
rect 4682 2022 4716 2024
rect 4654 2006 4728 2022
rect 4755 2018 4768 2032
rect 4783 2018 4799 2034
rect 4845 2029 4856 2042
rect 4638 1984 4639 2000
rect 4654 1984 4667 2006
rect 4682 1984 4712 2006
rect 4755 2002 4817 2018
rect 4845 2011 4856 2027
rect 4861 2022 4871 2042
rect 4881 2022 4895 2042
rect 4898 2029 4907 2042
rect 4923 2029 4932 2042
rect 4861 2011 4895 2022
rect 4898 2011 4907 2027
rect 4923 2011 4932 2027
rect 4939 2022 4949 2042
rect 4959 2022 4973 2042
rect 4974 2029 4985 2042
rect 4939 2011 4973 2022
rect 4974 2011 4985 2027
rect 5031 2018 5047 2034
rect 5054 2032 5084 2084
rect 5118 2080 5119 2087
rect 5103 2072 5119 2080
rect 5090 2040 5103 2059
rect 5118 2040 5148 2056
rect 5090 2024 5164 2040
rect 5090 2022 5103 2024
rect 5118 2022 5152 2024
rect 4755 2000 4768 2002
rect 4783 2000 4817 2002
rect 4755 1984 4817 2000
rect 4861 1995 4877 2002
rect 4939 1995 4969 2006
rect 5017 2002 5063 2018
rect 5090 2006 5164 2022
rect 5017 2000 5051 2002
rect 5016 1984 5063 2000
rect 5090 1984 5103 2006
rect 5118 1984 5148 2006
rect 5175 1984 5176 2000
rect 5191 1984 5204 2144
rect 5234 2040 5247 2144
rect 5292 2122 5293 2132
rect 5308 2122 5321 2132
rect 5292 2118 5321 2122
rect 5326 2118 5356 2144
rect 5374 2130 5390 2132
rect 5462 2130 5515 2144
rect 5463 2128 5527 2130
rect 5570 2128 5585 2144
rect 5634 2141 5664 2144
rect 5634 2138 5670 2141
rect 5600 2130 5616 2132
rect 5374 2118 5389 2122
rect 5292 2116 5389 2118
rect 5417 2116 5585 2128
rect 5601 2118 5616 2122
rect 5634 2119 5673 2138
rect 5692 2132 5699 2133
rect 5698 2125 5699 2132
rect 5682 2122 5683 2125
rect 5698 2122 5711 2125
rect 5634 2118 5664 2119
rect 5673 2118 5679 2119
rect 5682 2118 5711 2122
rect 5601 2117 5711 2118
rect 5601 2116 5717 2117
rect 5276 2108 5327 2116
rect 5276 2096 5301 2108
rect 5308 2096 5327 2108
rect 5358 2108 5408 2116
rect 5358 2100 5374 2108
rect 5381 2106 5408 2108
rect 5417 2106 5638 2116
rect 5381 2096 5638 2106
rect 5667 2108 5717 2116
rect 5667 2099 5683 2108
rect 5276 2088 5327 2096
rect 5374 2088 5638 2096
rect 5664 2096 5683 2099
rect 5690 2096 5717 2108
rect 5664 2088 5717 2096
rect 5292 2080 5293 2088
rect 5308 2080 5321 2088
rect 5292 2072 5308 2080
rect 5289 2065 5308 2068
rect 5289 2056 5311 2065
rect 5262 2046 5311 2056
rect 5262 2040 5292 2046
rect 5311 2041 5316 2046
rect 5234 2024 5308 2040
rect 5326 2032 5356 2088
rect 5391 2078 5599 2088
rect 5634 2084 5679 2088
rect 5682 2087 5683 2088
rect 5698 2087 5711 2088
rect 5417 2048 5606 2078
rect 5432 2045 5606 2048
rect 5425 2042 5606 2045
rect 5234 2022 5247 2024
rect 5262 2022 5296 2024
rect 5234 2006 5308 2022
rect 5335 2018 5348 2032
rect 5363 2018 5379 2034
rect 5425 2029 5436 2042
rect 5218 1984 5219 2000
rect 5234 1984 5247 2006
rect 5262 1984 5292 2006
rect 5335 2002 5397 2018
rect 5425 2011 5436 2027
rect 5441 2022 5451 2042
rect 5461 2022 5475 2042
rect 5478 2029 5487 2042
rect 5503 2029 5512 2042
rect 5441 2011 5475 2022
rect 5478 2011 5487 2027
rect 5503 2011 5512 2027
rect 5519 2022 5529 2042
rect 5539 2022 5553 2042
rect 5554 2029 5565 2042
rect 5519 2011 5553 2022
rect 5554 2011 5565 2027
rect 5611 2018 5627 2034
rect 5634 2032 5664 2084
rect 5698 2080 5699 2087
rect 5683 2072 5699 2080
rect 5670 2040 5683 2059
rect 5698 2040 5728 2056
rect 5670 2024 5744 2040
rect 5670 2022 5683 2024
rect 5698 2022 5732 2024
rect 5335 2000 5348 2002
rect 5363 2000 5397 2002
rect 5335 1984 5397 2000
rect 5441 1995 5457 2002
rect 5519 1995 5549 2006
rect 5597 2002 5643 2018
rect 5670 2006 5744 2022
rect 5597 2000 5631 2002
rect 5596 1984 5643 2000
rect 5670 1984 5683 2006
rect 5698 1984 5728 2006
rect 5755 1984 5756 2000
rect 5771 1984 5784 2144
rect 5814 2040 5827 2144
rect 5872 2122 5873 2132
rect 5888 2122 5901 2132
rect 5872 2118 5901 2122
rect 5906 2118 5936 2144
rect 5954 2130 5970 2132
rect 6042 2130 6095 2144
rect 6043 2128 6107 2130
rect 6150 2128 6165 2144
rect 6214 2141 6244 2144
rect 6214 2138 6250 2141
rect 6180 2130 6196 2132
rect 5954 2118 5969 2122
rect 5872 2116 5969 2118
rect 5997 2116 6165 2128
rect 6181 2118 6196 2122
rect 6214 2119 6253 2138
rect 6272 2132 6279 2133
rect 6278 2125 6279 2132
rect 6262 2122 6263 2125
rect 6278 2122 6291 2125
rect 6214 2118 6244 2119
rect 6253 2118 6259 2119
rect 6262 2118 6291 2122
rect 6181 2117 6291 2118
rect 6181 2116 6297 2117
rect 5856 2108 5907 2116
rect 5856 2096 5881 2108
rect 5888 2096 5907 2108
rect 5938 2108 5988 2116
rect 5938 2100 5954 2108
rect 5961 2106 5988 2108
rect 5997 2106 6218 2116
rect 5961 2096 6218 2106
rect 6247 2108 6297 2116
rect 6247 2099 6263 2108
rect 5856 2088 5907 2096
rect 5954 2088 6218 2096
rect 6244 2096 6263 2099
rect 6270 2096 6297 2108
rect 6244 2088 6297 2096
rect 5872 2080 5873 2088
rect 5888 2080 5901 2088
rect 5872 2072 5888 2080
rect 5869 2065 5888 2068
rect 5869 2056 5891 2065
rect 5842 2046 5891 2056
rect 5842 2040 5872 2046
rect 5891 2041 5896 2046
rect 5814 2024 5888 2040
rect 5906 2032 5936 2088
rect 5971 2078 6179 2088
rect 6214 2084 6259 2088
rect 6262 2087 6263 2088
rect 6278 2087 6291 2088
rect 5997 2048 6186 2078
rect 6012 2045 6186 2048
rect 6005 2042 6186 2045
rect 5814 2022 5827 2024
rect 5842 2022 5876 2024
rect 5814 2006 5888 2022
rect 5915 2018 5928 2032
rect 5943 2018 5959 2034
rect 6005 2029 6016 2042
rect 5798 1984 5799 2000
rect 5814 1984 5827 2006
rect 5842 1984 5872 2006
rect 5915 2002 5977 2018
rect 6005 2011 6016 2027
rect 6021 2022 6031 2042
rect 6041 2022 6055 2042
rect 6058 2029 6067 2042
rect 6083 2029 6092 2042
rect 6021 2011 6055 2022
rect 6058 2011 6067 2027
rect 6083 2011 6092 2027
rect 6099 2022 6109 2042
rect 6119 2022 6133 2042
rect 6134 2029 6145 2042
rect 6099 2011 6133 2022
rect 6134 2011 6145 2027
rect 6191 2018 6207 2034
rect 6214 2032 6244 2084
rect 6278 2080 6279 2087
rect 6263 2072 6279 2080
rect 6250 2040 6263 2059
rect 6278 2040 6308 2056
rect 6250 2024 6324 2040
rect 6250 2022 6263 2024
rect 6278 2022 6312 2024
rect 5915 2000 5928 2002
rect 5943 2000 5977 2002
rect 5915 1984 5977 2000
rect 6021 1995 6037 2002
rect 6099 1995 6129 2006
rect 6177 2002 6223 2018
rect 6250 2006 6324 2022
rect 6177 2000 6211 2002
rect 6176 1984 6223 2000
rect 6250 1984 6263 2006
rect 6278 1984 6308 2006
rect 6335 1984 6336 2000
rect 6351 1984 6364 2144
rect 6394 2040 6407 2144
rect 6452 2122 6453 2132
rect 6468 2122 6481 2132
rect 6452 2118 6481 2122
rect 6486 2118 6516 2144
rect 6534 2130 6550 2132
rect 6622 2130 6675 2144
rect 6623 2128 6687 2130
rect 6730 2128 6745 2144
rect 6794 2141 6824 2144
rect 6794 2138 6830 2141
rect 6760 2130 6776 2132
rect 6534 2118 6549 2122
rect 6452 2116 6549 2118
rect 6577 2116 6745 2128
rect 6761 2118 6776 2122
rect 6794 2119 6833 2138
rect 6852 2132 6859 2133
rect 6858 2125 6859 2132
rect 6842 2122 6843 2125
rect 6858 2122 6871 2125
rect 6794 2118 6824 2119
rect 6833 2118 6839 2119
rect 6842 2118 6871 2122
rect 6761 2117 6871 2118
rect 6761 2116 6877 2117
rect 6436 2108 6487 2116
rect 6436 2096 6461 2108
rect 6468 2096 6487 2108
rect 6518 2108 6568 2116
rect 6518 2100 6534 2108
rect 6541 2106 6568 2108
rect 6577 2106 6798 2116
rect 6541 2096 6798 2106
rect 6827 2108 6877 2116
rect 6827 2099 6843 2108
rect 6436 2088 6487 2096
rect 6534 2088 6798 2096
rect 6824 2096 6843 2099
rect 6850 2096 6877 2108
rect 6824 2088 6877 2096
rect 6452 2080 6453 2088
rect 6468 2080 6481 2088
rect 6452 2072 6468 2080
rect 6449 2065 6468 2068
rect 6449 2056 6471 2065
rect 6422 2046 6471 2056
rect 6422 2040 6452 2046
rect 6471 2041 6476 2046
rect 6394 2024 6468 2040
rect 6486 2032 6516 2088
rect 6551 2078 6759 2088
rect 6794 2084 6839 2088
rect 6842 2087 6843 2088
rect 6858 2087 6871 2088
rect 6577 2048 6766 2078
rect 6592 2045 6766 2048
rect 6585 2042 6766 2045
rect 6394 2022 6407 2024
rect 6422 2022 6456 2024
rect 6394 2006 6468 2022
rect 6495 2018 6508 2032
rect 6523 2018 6539 2034
rect 6585 2029 6596 2042
rect 6378 1984 6379 2000
rect 6394 1984 6407 2006
rect 6422 1984 6452 2006
rect 6495 2002 6557 2018
rect 6585 2011 6596 2027
rect 6601 2022 6611 2042
rect 6621 2022 6635 2042
rect 6638 2029 6647 2042
rect 6663 2029 6672 2042
rect 6601 2011 6635 2022
rect 6638 2011 6647 2027
rect 6663 2011 6672 2027
rect 6679 2022 6689 2042
rect 6699 2022 6713 2042
rect 6714 2029 6725 2042
rect 6679 2011 6713 2022
rect 6714 2011 6725 2027
rect 6771 2018 6787 2034
rect 6794 2032 6824 2084
rect 6858 2080 6859 2087
rect 6843 2072 6859 2080
rect 6830 2040 6843 2059
rect 6858 2040 6888 2056
rect 6830 2024 6904 2040
rect 6830 2022 6843 2024
rect 6858 2022 6892 2024
rect 6495 2000 6508 2002
rect 6523 2000 6557 2002
rect 6495 1984 6557 2000
rect 6601 1995 6617 2002
rect 6679 1995 6709 2006
rect 6757 2002 6803 2018
rect 6830 2006 6904 2022
rect 6757 2000 6791 2002
rect 6756 1984 6803 2000
rect 6830 1984 6843 2006
rect 6858 1984 6888 2006
rect 6915 1984 6916 2000
rect 6931 1984 6944 2144
rect -8 1976 33 1984
rect -8 1950 7 1976
rect 14 1950 33 1976
rect 97 1972 159 1984
rect 171 1972 246 1984
rect 304 1972 379 1984
rect 391 1972 422 1984
rect 428 1972 463 1984
rect 97 1970 259 1972
rect -8 1942 33 1950
rect 115 1946 128 1970
rect 143 1968 158 1970
rect -2 1932 -1 1942
rect 14 1932 27 1942
rect 42 1932 72 1946
rect 115 1932 158 1946
rect 182 1943 189 1950
rect 192 1946 259 1970
rect 291 1970 463 1972
rect 261 1948 289 1952
rect 291 1948 371 1970
rect 392 1968 407 1970
rect 261 1946 371 1948
rect 192 1942 371 1946
rect 165 1932 195 1942
rect 197 1932 350 1942
rect 358 1932 388 1942
rect 392 1932 422 1946
rect 450 1932 463 1970
rect 535 1976 570 1984
rect 535 1950 536 1976
rect 543 1950 570 1976
rect 478 1932 508 1946
rect 535 1942 570 1950
rect 572 1976 613 1984
rect 572 1950 587 1976
rect 594 1950 613 1976
rect 677 1972 739 1984
rect 751 1972 826 1984
rect 884 1972 959 1984
rect 971 1972 1002 1984
rect 1008 1972 1043 1984
rect 677 1970 839 1972
rect 572 1942 613 1950
rect 695 1946 708 1970
rect 723 1968 738 1970
rect 535 1932 536 1942
rect 551 1932 564 1942
rect 578 1932 579 1942
rect 594 1932 607 1942
rect 622 1932 652 1946
rect 695 1932 738 1946
rect 762 1943 769 1950
rect 772 1946 839 1970
rect 871 1970 1043 1972
rect 841 1948 869 1952
rect 871 1948 951 1970
rect 972 1968 987 1970
rect 841 1946 951 1948
rect 772 1942 951 1946
rect 745 1932 775 1942
rect 777 1932 930 1942
rect 938 1932 968 1942
rect 972 1932 1002 1946
rect 1030 1932 1043 1970
rect 1115 1976 1150 1984
rect 1115 1950 1116 1976
rect 1123 1950 1150 1976
rect 1058 1932 1088 1946
rect 1115 1942 1150 1950
rect 1152 1976 1193 1984
rect 1152 1950 1167 1976
rect 1174 1950 1193 1976
rect 1257 1972 1319 1984
rect 1331 1972 1406 1984
rect 1464 1972 1539 1984
rect 1551 1972 1582 1984
rect 1588 1972 1623 1984
rect 1257 1970 1419 1972
rect 1152 1942 1193 1950
rect 1275 1946 1288 1970
rect 1303 1968 1318 1970
rect 1115 1932 1116 1942
rect 1131 1932 1144 1942
rect 1158 1932 1159 1942
rect 1174 1932 1187 1942
rect 1202 1932 1232 1946
rect 1275 1932 1318 1946
rect 1342 1943 1349 1950
rect 1352 1946 1419 1970
rect 1451 1970 1623 1972
rect 1421 1948 1449 1952
rect 1451 1948 1531 1970
rect 1552 1968 1567 1970
rect 1421 1946 1531 1948
rect 1352 1942 1531 1946
rect 1325 1932 1355 1942
rect 1357 1932 1510 1942
rect 1518 1932 1548 1942
rect 1552 1932 1582 1946
rect 1610 1932 1623 1970
rect 1695 1976 1730 1984
rect 1695 1950 1696 1976
rect 1703 1950 1730 1976
rect 1638 1932 1668 1946
rect 1695 1942 1730 1950
rect 1732 1976 1773 1984
rect 1732 1950 1747 1976
rect 1754 1950 1773 1976
rect 1732 1942 1773 1950
rect 3481 1976 3513 1984
rect 3481 1950 3487 1976
rect 3494 1950 3513 1976
rect 3577 1972 3639 1984
rect 3651 1972 3726 1984
rect 3784 1972 3859 1984
rect 3871 1972 3902 1984
rect 3908 1972 3943 1984
rect 3577 1970 3739 1972
rect 1695 1932 1696 1942
rect 1711 1932 1724 1942
rect 1738 1932 1739 1942
rect 1754 1932 1767 1942
rect 1782 1932 1812 1946
rect 3481 1942 3513 1950
rect 3595 1946 3608 1970
rect 3623 1968 3638 1970
rect 3494 1932 3507 1942
rect 3522 1932 3552 1946
rect 3595 1932 3638 1946
rect 3662 1943 3669 1950
rect 3672 1946 3739 1970
rect 3771 1970 3943 1972
rect 3741 1948 3769 1952
rect 3771 1948 3851 1970
rect 3872 1968 3887 1970
rect 3741 1946 3851 1948
rect 3672 1942 3851 1946
rect 3645 1932 3675 1942
rect 3677 1932 3830 1942
rect 3838 1932 3868 1942
rect 3872 1932 3902 1946
rect 3930 1932 3943 1970
rect 4015 1976 4050 1984
rect 4015 1950 4016 1976
rect 4023 1950 4050 1976
rect 3958 1932 3988 1946
rect 4015 1942 4050 1950
rect 4052 1976 4093 1984
rect 4052 1950 4067 1976
rect 4074 1950 4093 1976
rect 4157 1972 4219 1984
rect 4231 1972 4306 1984
rect 4364 1972 4439 1984
rect 4451 1972 4482 1984
rect 4488 1972 4523 1984
rect 4157 1970 4319 1972
rect 4052 1942 4093 1950
rect 4175 1946 4188 1970
rect 4203 1968 4218 1970
rect 4015 1932 4016 1942
rect 4031 1932 4044 1942
rect 4058 1932 4059 1942
rect 4074 1932 4087 1942
rect 4102 1932 4132 1946
rect 4175 1932 4218 1946
rect 4242 1943 4249 1950
rect 4252 1946 4319 1970
rect 4351 1970 4523 1972
rect 4321 1948 4349 1952
rect 4351 1948 4431 1970
rect 4452 1968 4467 1970
rect 4321 1946 4431 1948
rect 4252 1942 4431 1946
rect 4225 1932 4255 1942
rect 4257 1932 4410 1942
rect 4418 1932 4448 1942
rect 4452 1932 4482 1946
rect 4510 1932 4523 1970
rect 4595 1976 4630 1984
rect 4595 1950 4596 1976
rect 4603 1950 4630 1976
rect 4538 1932 4568 1946
rect 4595 1942 4630 1950
rect 4632 1976 4673 1984
rect 4632 1950 4647 1976
rect 4654 1950 4673 1976
rect 4737 1972 4799 1984
rect 4811 1972 4886 1984
rect 4944 1972 5019 1984
rect 5031 1972 5062 1984
rect 5068 1972 5103 1984
rect 4737 1970 4899 1972
rect 4632 1942 4673 1950
rect 4755 1946 4768 1970
rect 4783 1968 4798 1970
rect 4595 1932 4596 1942
rect 4611 1932 4624 1942
rect 4638 1932 4639 1942
rect 4654 1932 4667 1942
rect 4682 1932 4712 1946
rect 4755 1932 4798 1946
rect 4822 1943 4829 1950
rect 4832 1946 4899 1970
rect 4931 1970 5103 1972
rect 4901 1948 4929 1952
rect 4931 1948 5011 1970
rect 5032 1968 5047 1970
rect 4901 1946 5011 1948
rect 4832 1942 5011 1946
rect 4805 1932 4835 1942
rect 4837 1932 4990 1942
rect 4998 1932 5028 1942
rect 5032 1932 5062 1946
rect 5090 1932 5103 1970
rect 5175 1976 5210 1984
rect 5175 1950 5176 1976
rect 5183 1950 5210 1976
rect 5118 1932 5148 1946
rect 5175 1942 5210 1950
rect 5212 1976 5253 1984
rect 5212 1950 5227 1976
rect 5234 1950 5253 1976
rect 5317 1972 5379 1984
rect 5391 1972 5466 1984
rect 5524 1972 5599 1984
rect 5611 1972 5642 1984
rect 5648 1972 5683 1984
rect 5317 1970 5479 1972
rect 5212 1942 5253 1950
rect 5335 1946 5348 1970
rect 5363 1968 5378 1970
rect 5175 1932 5176 1942
rect 5191 1932 5204 1942
rect 5218 1932 5219 1942
rect 5234 1932 5247 1942
rect 5262 1932 5292 1946
rect 5335 1932 5378 1946
rect 5402 1943 5409 1950
rect 5412 1946 5479 1970
rect 5511 1970 5683 1972
rect 5481 1948 5509 1952
rect 5511 1948 5591 1970
rect 5612 1968 5627 1970
rect 5481 1946 5591 1948
rect 5412 1942 5591 1946
rect 5385 1932 5415 1942
rect 5417 1932 5570 1942
rect 5578 1932 5608 1942
rect 5612 1932 5642 1946
rect 5670 1932 5683 1970
rect 5755 1976 5790 1984
rect 5755 1950 5756 1976
rect 5763 1950 5790 1976
rect 5698 1932 5728 1946
rect 5755 1942 5790 1950
rect 5792 1976 5833 1984
rect 5792 1950 5807 1976
rect 5814 1950 5833 1976
rect 5897 1972 5959 1984
rect 5971 1972 6046 1984
rect 6104 1972 6179 1984
rect 6191 1972 6222 1984
rect 6228 1972 6263 1984
rect 5897 1970 6059 1972
rect 5792 1942 5833 1950
rect 5915 1946 5928 1970
rect 5943 1968 5958 1970
rect 5755 1932 5756 1942
rect 5771 1932 5784 1942
rect 5798 1932 5799 1942
rect 5814 1932 5827 1942
rect 5842 1932 5872 1946
rect 5915 1932 5958 1946
rect 5982 1943 5989 1950
rect 5992 1946 6059 1970
rect 6091 1970 6263 1972
rect 6061 1948 6089 1952
rect 6091 1948 6171 1970
rect 6192 1968 6207 1970
rect 6061 1946 6171 1948
rect 5992 1942 6171 1946
rect 5965 1932 5995 1942
rect 5997 1932 6150 1942
rect 6158 1932 6188 1942
rect 6192 1932 6222 1946
rect 6250 1932 6263 1970
rect 6335 1976 6370 1984
rect 6335 1950 6336 1976
rect 6343 1950 6370 1976
rect 6278 1932 6308 1946
rect 6335 1942 6370 1950
rect 6372 1976 6413 1984
rect 6372 1950 6387 1976
rect 6394 1950 6413 1976
rect 6477 1972 6539 1984
rect 6551 1972 6626 1984
rect 6684 1972 6759 1984
rect 6771 1972 6802 1984
rect 6808 1972 6843 1984
rect 6477 1970 6639 1972
rect 6372 1942 6413 1950
rect 6495 1946 6508 1970
rect 6523 1968 6538 1970
rect 6335 1932 6336 1942
rect 6351 1932 6364 1942
rect 6378 1932 6379 1942
rect 6394 1932 6407 1942
rect 6422 1932 6452 1946
rect 6495 1932 6538 1946
rect 6562 1943 6569 1950
rect 6572 1946 6639 1970
rect 6671 1970 6843 1972
rect 6641 1948 6669 1952
rect 6671 1948 6751 1970
rect 6772 1968 6787 1970
rect 6641 1946 6751 1948
rect 6572 1942 6751 1946
rect 6545 1932 6575 1942
rect 6577 1932 6730 1942
rect 6738 1932 6768 1942
rect 6772 1932 6802 1946
rect 6830 1932 6843 1970
rect 6915 1976 6950 1984
rect 6915 1950 6916 1976
rect 6923 1950 6950 1976
rect 6858 1932 6888 1946
rect 6915 1942 6950 1950
rect 6915 1932 6916 1942
rect 6931 1932 6944 1942
rect -2 1926 1837 1932
rect -1 1918 1837 1926
rect 3481 1918 6944 1932
rect 14 1888 27 1918
rect 42 1900 72 1918
rect 115 1904 129 1918
rect 165 1904 385 1918
rect 116 1902 129 1904
rect 82 1890 97 1902
rect 79 1888 101 1890
rect 106 1888 136 1902
rect 197 1900 350 1904
rect 179 1888 371 1900
rect 414 1888 444 1902
rect 450 1888 463 1918
rect 478 1900 508 1918
rect 551 1888 564 1918
rect 594 1888 607 1918
rect 622 1900 652 1918
rect 695 1904 709 1918
rect 745 1904 965 1918
rect 696 1902 709 1904
rect 662 1890 677 1902
rect 659 1888 681 1890
rect 686 1888 716 1902
rect 777 1900 930 1904
rect 759 1888 951 1900
rect 994 1888 1024 1902
rect 1030 1888 1043 1918
rect 1058 1900 1088 1918
rect 1131 1888 1144 1918
rect 1174 1888 1187 1918
rect 1202 1900 1232 1918
rect 1275 1904 1289 1918
rect 1325 1904 1545 1918
rect 1276 1902 1289 1904
rect 1242 1890 1257 1902
rect 1239 1888 1261 1890
rect 1266 1888 1296 1902
rect 1357 1900 1510 1904
rect 1339 1888 1531 1900
rect 1574 1888 1604 1902
rect 1610 1888 1623 1918
rect 1638 1900 1668 1918
rect 1711 1888 1724 1918
rect 1754 1888 1767 1918
rect 1782 1900 1812 1918
rect 1822 1890 1837 1902
rect 1819 1888 1837 1890
rect 3494 1888 3507 1918
rect 3522 1900 3552 1918
rect 3595 1904 3609 1918
rect 3645 1904 3865 1918
rect 3596 1902 3609 1904
rect 3562 1890 3577 1902
rect 3559 1888 3581 1890
rect 3586 1888 3616 1902
rect 3677 1900 3830 1904
rect 3659 1888 3851 1900
rect 3894 1888 3924 1902
rect 3930 1888 3943 1918
rect 3958 1900 3988 1918
rect 4031 1888 4044 1918
rect 4074 1888 4087 1918
rect 4102 1900 4132 1918
rect 4175 1904 4189 1918
rect 4225 1904 4445 1918
rect 4176 1902 4189 1904
rect 4142 1890 4157 1902
rect 4139 1888 4161 1890
rect 4166 1888 4196 1902
rect 4257 1900 4410 1904
rect 4239 1888 4431 1900
rect 4474 1888 4504 1902
rect 4510 1888 4523 1918
rect 4538 1900 4568 1918
rect 4611 1888 4624 1918
rect 4654 1888 4667 1918
rect 4682 1900 4712 1918
rect 4755 1904 4769 1918
rect 4805 1904 5025 1918
rect 4756 1902 4769 1904
rect 4722 1890 4737 1902
rect 4719 1888 4741 1890
rect 4746 1888 4776 1902
rect 4837 1900 4990 1904
rect 4819 1888 5011 1900
rect 5054 1888 5084 1902
rect 5090 1888 5103 1918
rect 5118 1900 5148 1918
rect 5191 1888 5204 1918
rect 5234 1888 5247 1918
rect 5262 1900 5292 1918
rect 5335 1904 5349 1918
rect 5385 1904 5605 1918
rect 5336 1902 5349 1904
rect 5302 1890 5317 1902
rect 5299 1888 5321 1890
rect 5326 1888 5356 1902
rect 5417 1900 5570 1904
rect 5399 1888 5591 1900
rect 5634 1888 5664 1902
rect 5670 1888 5683 1918
rect 5698 1900 5728 1918
rect 5771 1888 5784 1918
rect 5814 1888 5827 1918
rect 5842 1900 5872 1918
rect 5915 1904 5929 1918
rect 5965 1904 6185 1918
rect 5916 1902 5929 1904
rect 5882 1890 5897 1902
rect 5879 1888 5901 1890
rect 5906 1888 5936 1902
rect 5997 1900 6150 1904
rect 5979 1888 6171 1900
rect 6214 1888 6244 1902
rect 6250 1888 6263 1918
rect 6278 1900 6308 1918
rect 6351 1888 6364 1918
rect 6394 1888 6407 1918
rect 6422 1900 6452 1918
rect 6495 1904 6509 1918
rect 6545 1904 6765 1918
rect 6496 1902 6509 1904
rect 6462 1890 6477 1902
rect 6459 1888 6481 1890
rect 6486 1888 6516 1902
rect 6577 1900 6730 1904
rect 6559 1888 6751 1900
rect 6794 1888 6824 1902
rect 6830 1888 6843 1918
rect 6858 1900 6888 1918
rect 6931 1888 6944 1918
rect -1 1874 1837 1888
rect 3481 1874 6944 1888
rect 14 1770 27 1874
rect 72 1852 73 1862
rect 88 1852 101 1862
rect 72 1848 101 1852
rect 106 1848 136 1874
rect 154 1860 170 1862
rect 242 1860 295 1874
rect 243 1858 307 1860
rect 350 1858 365 1874
rect 414 1871 444 1874
rect 414 1868 450 1871
rect 380 1860 396 1862
rect 154 1848 169 1852
rect 72 1846 169 1848
rect 197 1846 365 1858
rect 381 1848 396 1852
rect 414 1849 453 1868
rect 472 1862 479 1863
rect 478 1855 479 1862
rect 462 1852 463 1855
rect 478 1852 491 1855
rect 414 1848 444 1849
rect 453 1848 459 1849
rect 462 1848 491 1852
rect 381 1847 491 1848
rect 381 1846 497 1847
rect 56 1838 107 1846
rect 56 1826 81 1838
rect 88 1826 107 1838
rect 138 1838 188 1846
rect 138 1830 154 1838
rect 161 1836 188 1838
rect 197 1836 418 1846
rect 161 1826 418 1836
rect 447 1838 497 1846
rect 447 1829 463 1838
rect 56 1818 107 1826
rect 154 1818 418 1826
rect 444 1826 463 1829
rect 470 1826 497 1838
rect 444 1818 497 1826
rect 72 1810 73 1818
rect 88 1810 101 1818
rect 72 1802 88 1810
rect 69 1795 88 1798
rect 69 1786 91 1795
rect 42 1776 91 1786
rect 42 1770 72 1776
rect 91 1771 96 1776
rect 14 1754 88 1770
rect 106 1762 136 1818
rect 171 1808 379 1818
rect 414 1814 459 1818
rect 462 1817 463 1818
rect 478 1817 491 1818
rect 197 1778 386 1808
rect 212 1775 386 1778
rect 205 1772 386 1775
rect 14 1752 27 1754
rect 42 1752 76 1754
rect 14 1736 88 1752
rect 115 1748 128 1762
rect 143 1748 159 1764
rect 205 1759 216 1772
rect -2 1714 -1 1730
rect 14 1714 27 1736
rect 42 1714 72 1736
rect 115 1732 177 1748
rect 205 1741 216 1757
rect 221 1752 231 1772
rect 241 1752 255 1772
rect 258 1759 267 1772
rect 283 1759 292 1772
rect 221 1741 255 1752
rect 258 1741 267 1757
rect 283 1741 292 1757
rect 299 1752 309 1772
rect 319 1752 333 1772
rect 334 1759 345 1772
rect 299 1741 333 1752
rect 334 1741 345 1757
rect 391 1748 407 1764
rect 414 1762 444 1814
rect 478 1810 479 1817
rect 463 1802 479 1810
rect 450 1770 463 1789
rect 478 1770 508 1786
rect 450 1754 524 1770
rect 450 1752 463 1754
rect 478 1752 512 1754
rect 115 1730 128 1732
rect 143 1730 177 1732
rect 115 1714 177 1730
rect 221 1725 237 1732
rect 299 1725 329 1736
rect 377 1732 423 1748
rect 450 1736 524 1752
rect 377 1730 411 1732
rect 376 1714 423 1730
rect 450 1714 463 1736
rect 478 1714 508 1736
rect 535 1714 536 1730
rect 551 1714 564 1874
rect 594 1770 607 1874
rect 652 1852 653 1862
rect 668 1852 681 1862
rect 652 1848 681 1852
rect 686 1848 716 1874
rect 734 1860 750 1862
rect 822 1860 875 1874
rect 823 1858 887 1860
rect 930 1858 945 1874
rect 994 1871 1024 1874
rect 994 1868 1030 1871
rect 960 1860 976 1862
rect 734 1848 749 1852
rect 652 1846 749 1848
rect 777 1846 945 1858
rect 961 1848 976 1852
rect 994 1849 1033 1868
rect 1052 1862 1059 1863
rect 1058 1855 1059 1862
rect 1042 1852 1043 1855
rect 1058 1852 1071 1855
rect 994 1848 1024 1849
rect 1033 1848 1039 1849
rect 1042 1848 1071 1852
rect 961 1847 1071 1848
rect 961 1846 1077 1847
rect 636 1838 687 1846
rect 636 1826 661 1838
rect 668 1826 687 1838
rect 718 1838 768 1846
rect 718 1830 734 1838
rect 741 1836 768 1838
rect 777 1836 998 1846
rect 741 1826 998 1836
rect 1027 1838 1077 1846
rect 1027 1829 1043 1838
rect 636 1818 687 1826
rect 734 1818 998 1826
rect 1024 1826 1043 1829
rect 1050 1826 1077 1838
rect 1024 1818 1077 1826
rect 652 1810 653 1818
rect 668 1810 681 1818
rect 652 1802 668 1810
rect 649 1795 668 1798
rect 649 1786 671 1795
rect 622 1776 671 1786
rect 622 1770 652 1776
rect 671 1771 676 1776
rect 594 1754 668 1770
rect 686 1762 716 1818
rect 751 1808 959 1818
rect 994 1814 1039 1818
rect 1042 1817 1043 1818
rect 1058 1817 1071 1818
rect 777 1778 966 1808
rect 792 1775 966 1778
rect 785 1772 966 1775
rect 594 1752 607 1754
rect 622 1752 656 1754
rect 594 1736 668 1752
rect 695 1748 708 1762
rect 723 1748 739 1764
rect 785 1759 796 1772
rect 578 1714 579 1730
rect 594 1714 607 1736
rect 622 1714 652 1736
rect 695 1732 757 1748
rect 785 1741 796 1757
rect 801 1752 811 1772
rect 821 1752 835 1772
rect 838 1759 847 1772
rect 863 1759 872 1772
rect 801 1741 835 1752
rect 838 1741 847 1757
rect 863 1741 872 1757
rect 879 1752 889 1772
rect 899 1752 913 1772
rect 914 1759 925 1772
rect 879 1741 913 1752
rect 914 1741 925 1757
rect 971 1748 987 1764
rect 994 1762 1024 1814
rect 1058 1810 1059 1817
rect 1043 1802 1059 1810
rect 1030 1770 1043 1789
rect 1058 1770 1088 1786
rect 1030 1754 1104 1770
rect 1030 1752 1043 1754
rect 1058 1752 1092 1754
rect 695 1730 708 1732
rect 723 1730 757 1732
rect 695 1714 757 1730
rect 801 1725 817 1732
rect 879 1725 909 1736
rect 957 1732 1003 1748
rect 1030 1736 1104 1752
rect 957 1730 991 1732
rect 956 1714 1003 1730
rect 1030 1714 1043 1736
rect 1058 1714 1088 1736
rect 1115 1714 1116 1730
rect 1131 1714 1144 1874
rect 1174 1770 1187 1874
rect 1232 1852 1233 1862
rect 1248 1852 1261 1862
rect 1232 1848 1261 1852
rect 1266 1848 1296 1874
rect 1314 1860 1330 1862
rect 1402 1860 1455 1874
rect 1403 1858 1467 1860
rect 1510 1858 1525 1874
rect 1574 1871 1604 1874
rect 1574 1868 1610 1871
rect 1540 1860 1556 1862
rect 1314 1848 1329 1852
rect 1232 1846 1329 1848
rect 1357 1846 1525 1858
rect 1541 1848 1556 1852
rect 1574 1849 1613 1868
rect 1632 1862 1639 1863
rect 1638 1855 1639 1862
rect 1622 1852 1623 1855
rect 1638 1852 1651 1855
rect 1574 1848 1604 1849
rect 1613 1848 1619 1849
rect 1622 1848 1651 1852
rect 1541 1847 1651 1848
rect 1541 1846 1657 1847
rect 1216 1838 1267 1846
rect 1216 1826 1241 1838
rect 1248 1826 1267 1838
rect 1298 1838 1348 1846
rect 1298 1830 1314 1838
rect 1321 1836 1348 1838
rect 1357 1836 1578 1846
rect 1321 1826 1578 1836
rect 1607 1838 1657 1846
rect 1607 1829 1623 1838
rect 1216 1818 1267 1826
rect 1314 1818 1578 1826
rect 1604 1826 1623 1829
rect 1630 1826 1657 1838
rect 1604 1818 1657 1826
rect 1232 1810 1233 1818
rect 1248 1810 1261 1818
rect 1232 1802 1248 1810
rect 1229 1795 1248 1798
rect 1229 1786 1251 1795
rect 1202 1776 1251 1786
rect 1202 1770 1232 1776
rect 1251 1771 1256 1776
rect 1174 1754 1248 1770
rect 1266 1762 1296 1818
rect 1331 1808 1539 1818
rect 1574 1814 1619 1818
rect 1622 1817 1623 1818
rect 1638 1817 1651 1818
rect 1357 1778 1546 1808
rect 1372 1775 1546 1778
rect 1365 1772 1546 1775
rect 1174 1752 1187 1754
rect 1202 1752 1236 1754
rect 1174 1736 1248 1752
rect 1275 1748 1288 1762
rect 1303 1748 1319 1764
rect 1365 1759 1376 1772
rect 1158 1714 1159 1730
rect 1174 1714 1187 1736
rect 1202 1714 1232 1736
rect 1275 1732 1337 1748
rect 1365 1741 1376 1757
rect 1381 1752 1391 1772
rect 1401 1752 1415 1772
rect 1418 1759 1427 1772
rect 1443 1759 1452 1772
rect 1381 1741 1415 1752
rect 1418 1741 1427 1757
rect 1443 1741 1452 1757
rect 1459 1752 1469 1772
rect 1479 1752 1493 1772
rect 1494 1759 1505 1772
rect 1459 1741 1493 1752
rect 1494 1741 1505 1757
rect 1551 1748 1567 1764
rect 1574 1762 1604 1814
rect 1638 1810 1639 1817
rect 1623 1802 1639 1810
rect 1610 1770 1623 1789
rect 1638 1770 1668 1786
rect 1610 1754 1684 1770
rect 1610 1752 1623 1754
rect 1638 1752 1672 1754
rect 1275 1730 1288 1732
rect 1303 1730 1337 1732
rect 1275 1714 1337 1730
rect 1381 1725 1397 1732
rect 1459 1725 1489 1736
rect 1537 1732 1583 1748
rect 1610 1736 1684 1752
rect 1537 1730 1571 1732
rect 1536 1714 1583 1730
rect 1610 1714 1623 1736
rect 1638 1714 1668 1736
rect 1695 1714 1696 1730
rect 1711 1714 1724 1874
rect 1754 1770 1767 1874
rect 1812 1852 1813 1862
rect 1828 1852 1837 1862
rect 1812 1846 1837 1852
rect 1796 1838 1837 1846
rect 1796 1826 1821 1838
rect 1828 1826 1837 1838
rect 1796 1818 1837 1826
rect 1812 1810 1813 1818
rect 1828 1810 1837 1818
rect 1812 1802 1828 1810
rect 1809 1795 1828 1798
rect 1809 1786 1831 1795
rect 1782 1776 1831 1786
rect 1782 1770 1812 1776
rect 1831 1771 1836 1776
rect 3494 1770 3507 1874
rect 3552 1852 3553 1862
rect 3568 1852 3581 1862
rect 3552 1848 3581 1852
rect 3586 1848 3616 1874
rect 3634 1860 3650 1862
rect 3722 1860 3775 1874
rect 3723 1858 3787 1860
rect 3830 1858 3845 1874
rect 3894 1871 3924 1874
rect 3894 1868 3930 1871
rect 3860 1860 3876 1862
rect 3634 1848 3649 1852
rect 3552 1846 3649 1848
rect 3677 1846 3845 1858
rect 3861 1848 3876 1852
rect 3894 1849 3933 1868
rect 3952 1862 3959 1863
rect 3958 1855 3959 1862
rect 3942 1852 3943 1855
rect 3958 1852 3971 1855
rect 3894 1848 3924 1849
rect 3933 1848 3939 1849
rect 3942 1848 3971 1852
rect 3861 1847 3971 1848
rect 3861 1846 3977 1847
rect 3536 1838 3587 1846
rect 3536 1826 3561 1838
rect 3568 1826 3587 1838
rect 3618 1838 3668 1846
rect 3618 1830 3634 1838
rect 3641 1836 3668 1838
rect 3677 1836 3898 1846
rect 3641 1826 3898 1836
rect 3927 1838 3977 1846
rect 3927 1829 3943 1838
rect 3536 1818 3587 1826
rect 3634 1818 3898 1826
rect 3924 1826 3943 1829
rect 3950 1826 3977 1838
rect 3924 1818 3977 1826
rect 3552 1810 3553 1818
rect 3568 1810 3581 1818
rect 3552 1802 3568 1810
rect 3549 1795 3568 1798
rect 3549 1786 3571 1795
rect 3522 1776 3571 1786
rect 3522 1770 3552 1776
rect 3571 1771 3576 1776
rect 1754 1754 1828 1770
rect 3494 1754 3568 1770
rect 3586 1762 3616 1818
rect 3651 1808 3859 1818
rect 3894 1814 3939 1818
rect 3942 1817 3943 1818
rect 3958 1817 3971 1818
rect 3677 1778 3866 1808
rect 3692 1775 3866 1778
rect 3685 1772 3866 1775
rect 1754 1752 1767 1754
rect 1782 1752 1816 1754
rect 3494 1752 3507 1754
rect 3522 1752 3556 1754
rect 1754 1736 1828 1752
rect 3494 1736 3568 1752
rect 3595 1748 3608 1762
rect 3623 1748 3639 1764
rect 3685 1759 3696 1772
rect 1738 1714 1739 1730
rect 1754 1714 1767 1736
rect 1782 1714 1812 1736
rect 3494 1714 3507 1736
rect 3522 1714 3552 1736
rect 3595 1732 3657 1748
rect 3685 1741 3696 1757
rect 3701 1752 3711 1772
rect 3721 1752 3735 1772
rect 3738 1759 3747 1772
rect 3763 1759 3772 1772
rect 3701 1741 3735 1752
rect 3738 1741 3747 1757
rect 3763 1741 3772 1757
rect 3779 1752 3789 1772
rect 3799 1752 3813 1772
rect 3814 1759 3825 1772
rect 3779 1741 3813 1752
rect 3814 1741 3825 1757
rect 3871 1748 3887 1764
rect 3894 1762 3924 1814
rect 3958 1810 3959 1817
rect 3943 1802 3959 1810
rect 3930 1770 3943 1789
rect 3958 1770 3988 1786
rect 3930 1754 4004 1770
rect 3930 1752 3943 1754
rect 3958 1752 3992 1754
rect 3595 1730 3608 1732
rect 3623 1730 3657 1732
rect 3595 1714 3657 1730
rect 3701 1725 3717 1732
rect 3779 1725 3809 1736
rect 3857 1732 3903 1748
rect 3930 1736 4004 1752
rect 3857 1730 3891 1732
rect 3856 1714 3903 1730
rect 3930 1714 3943 1736
rect 3958 1714 3988 1736
rect 4015 1714 4016 1730
rect 4031 1714 4044 1874
rect 4074 1770 4087 1874
rect 4132 1852 4133 1862
rect 4148 1852 4161 1862
rect 4132 1848 4161 1852
rect 4166 1848 4196 1874
rect 4214 1860 4230 1862
rect 4302 1860 4355 1874
rect 4303 1858 4367 1860
rect 4410 1858 4425 1874
rect 4474 1871 4504 1874
rect 4474 1868 4510 1871
rect 4440 1860 4456 1862
rect 4214 1848 4229 1852
rect 4132 1846 4229 1848
rect 4257 1846 4425 1858
rect 4441 1848 4456 1852
rect 4474 1849 4513 1868
rect 4532 1862 4539 1863
rect 4538 1855 4539 1862
rect 4522 1852 4523 1855
rect 4538 1852 4551 1855
rect 4474 1848 4504 1849
rect 4513 1848 4519 1849
rect 4522 1848 4551 1852
rect 4441 1847 4551 1848
rect 4441 1846 4557 1847
rect 4116 1838 4167 1846
rect 4116 1826 4141 1838
rect 4148 1826 4167 1838
rect 4198 1838 4248 1846
rect 4198 1830 4214 1838
rect 4221 1836 4248 1838
rect 4257 1836 4478 1846
rect 4221 1826 4478 1836
rect 4507 1838 4557 1846
rect 4507 1829 4523 1838
rect 4116 1818 4167 1826
rect 4214 1818 4478 1826
rect 4504 1826 4523 1829
rect 4530 1826 4557 1838
rect 4504 1818 4557 1826
rect 4132 1810 4133 1818
rect 4148 1810 4161 1818
rect 4132 1802 4148 1810
rect 4129 1795 4148 1798
rect 4129 1786 4151 1795
rect 4102 1776 4151 1786
rect 4102 1770 4132 1776
rect 4151 1771 4156 1776
rect 4074 1754 4148 1770
rect 4166 1762 4196 1818
rect 4231 1808 4439 1818
rect 4474 1814 4519 1818
rect 4522 1817 4523 1818
rect 4538 1817 4551 1818
rect 4257 1778 4446 1808
rect 4272 1775 4446 1778
rect 4265 1772 4446 1775
rect 4074 1752 4087 1754
rect 4102 1752 4136 1754
rect 4074 1736 4148 1752
rect 4175 1748 4188 1762
rect 4203 1748 4219 1764
rect 4265 1759 4276 1772
rect 4058 1714 4059 1730
rect 4074 1714 4087 1736
rect 4102 1714 4132 1736
rect 4175 1732 4237 1748
rect 4265 1741 4276 1757
rect 4281 1752 4291 1772
rect 4301 1752 4315 1772
rect 4318 1759 4327 1772
rect 4343 1759 4352 1772
rect 4281 1741 4315 1752
rect 4318 1741 4327 1757
rect 4343 1741 4352 1757
rect 4359 1752 4369 1772
rect 4379 1752 4393 1772
rect 4394 1759 4405 1772
rect 4359 1741 4393 1752
rect 4394 1741 4405 1757
rect 4451 1748 4467 1764
rect 4474 1762 4504 1814
rect 4538 1810 4539 1817
rect 4523 1802 4539 1810
rect 4510 1770 4523 1789
rect 4538 1770 4568 1786
rect 4510 1754 4584 1770
rect 4510 1752 4523 1754
rect 4538 1752 4572 1754
rect 4175 1730 4188 1732
rect 4203 1730 4237 1732
rect 4175 1714 4237 1730
rect 4281 1725 4297 1732
rect 4359 1725 4389 1736
rect 4437 1732 4483 1748
rect 4510 1736 4584 1752
rect 4437 1730 4471 1732
rect 4436 1714 4483 1730
rect 4510 1714 4523 1736
rect 4538 1714 4568 1736
rect 4595 1714 4596 1730
rect 4611 1714 4624 1874
rect 4654 1770 4667 1874
rect 4712 1852 4713 1862
rect 4728 1852 4741 1862
rect 4712 1848 4741 1852
rect 4746 1848 4776 1874
rect 4794 1860 4810 1862
rect 4882 1860 4935 1874
rect 4883 1858 4947 1860
rect 4990 1858 5005 1874
rect 5054 1871 5084 1874
rect 5054 1868 5090 1871
rect 5020 1860 5036 1862
rect 4794 1848 4809 1852
rect 4712 1846 4809 1848
rect 4837 1846 5005 1858
rect 5021 1848 5036 1852
rect 5054 1849 5093 1868
rect 5112 1862 5119 1863
rect 5118 1855 5119 1862
rect 5102 1852 5103 1855
rect 5118 1852 5131 1855
rect 5054 1848 5084 1849
rect 5093 1848 5099 1849
rect 5102 1848 5131 1852
rect 5021 1847 5131 1848
rect 5021 1846 5137 1847
rect 4696 1838 4747 1846
rect 4696 1826 4721 1838
rect 4728 1826 4747 1838
rect 4778 1838 4828 1846
rect 4778 1830 4794 1838
rect 4801 1836 4828 1838
rect 4837 1836 5058 1846
rect 4801 1826 5058 1836
rect 5087 1838 5137 1846
rect 5087 1829 5103 1838
rect 4696 1818 4747 1826
rect 4794 1818 5058 1826
rect 5084 1826 5103 1829
rect 5110 1826 5137 1838
rect 5084 1818 5137 1826
rect 4712 1810 4713 1818
rect 4728 1810 4741 1818
rect 4712 1802 4728 1810
rect 4709 1795 4728 1798
rect 4709 1786 4731 1795
rect 4682 1776 4731 1786
rect 4682 1770 4712 1776
rect 4731 1771 4736 1776
rect 4654 1754 4728 1770
rect 4746 1762 4776 1818
rect 4811 1808 5019 1818
rect 5054 1814 5099 1818
rect 5102 1817 5103 1818
rect 5118 1817 5131 1818
rect 4837 1778 5026 1808
rect 4852 1775 5026 1778
rect 4845 1772 5026 1775
rect 4654 1752 4667 1754
rect 4682 1752 4716 1754
rect 4654 1736 4728 1752
rect 4755 1748 4768 1762
rect 4783 1748 4799 1764
rect 4845 1759 4856 1772
rect 4638 1714 4639 1730
rect 4654 1714 4667 1736
rect 4682 1714 4712 1736
rect 4755 1732 4817 1748
rect 4845 1741 4856 1757
rect 4861 1752 4871 1772
rect 4881 1752 4895 1772
rect 4898 1759 4907 1772
rect 4923 1759 4932 1772
rect 4861 1741 4895 1752
rect 4898 1741 4907 1757
rect 4923 1741 4932 1757
rect 4939 1752 4949 1772
rect 4959 1752 4973 1772
rect 4974 1759 4985 1772
rect 4939 1741 4973 1752
rect 4974 1741 4985 1757
rect 5031 1748 5047 1764
rect 5054 1762 5084 1814
rect 5118 1810 5119 1817
rect 5103 1802 5119 1810
rect 5090 1770 5103 1789
rect 5118 1770 5148 1786
rect 5090 1754 5164 1770
rect 5090 1752 5103 1754
rect 5118 1752 5152 1754
rect 4755 1730 4768 1732
rect 4783 1730 4817 1732
rect 4755 1714 4817 1730
rect 4861 1725 4877 1732
rect 4939 1725 4969 1736
rect 5017 1732 5063 1748
rect 5090 1736 5164 1752
rect 5017 1730 5051 1732
rect 5016 1714 5063 1730
rect 5090 1714 5103 1736
rect 5118 1714 5148 1736
rect 5175 1714 5176 1730
rect 5191 1714 5204 1874
rect 5234 1770 5247 1874
rect 5292 1852 5293 1862
rect 5308 1852 5321 1862
rect 5292 1848 5321 1852
rect 5326 1848 5356 1874
rect 5374 1860 5390 1862
rect 5462 1860 5515 1874
rect 5463 1858 5527 1860
rect 5570 1858 5585 1874
rect 5634 1871 5664 1874
rect 5634 1868 5670 1871
rect 5600 1860 5616 1862
rect 5374 1848 5389 1852
rect 5292 1846 5389 1848
rect 5417 1846 5585 1858
rect 5601 1848 5616 1852
rect 5634 1849 5673 1868
rect 5692 1862 5699 1863
rect 5698 1855 5699 1862
rect 5682 1852 5683 1855
rect 5698 1852 5711 1855
rect 5634 1848 5664 1849
rect 5673 1848 5679 1849
rect 5682 1848 5711 1852
rect 5601 1847 5711 1848
rect 5601 1846 5717 1847
rect 5276 1838 5327 1846
rect 5276 1826 5301 1838
rect 5308 1826 5327 1838
rect 5358 1838 5408 1846
rect 5358 1830 5374 1838
rect 5381 1836 5408 1838
rect 5417 1836 5638 1846
rect 5381 1826 5638 1836
rect 5667 1838 5717 1846
rect 5667 1829 5683 1838
rect 5276 1818 5327 1826
rect 5374 1818 5638 1826
rect 5664 1826 5683 1829
rect 5690 1826 5717 1838
rect 5664 1818 5717 1826
rect 5292 1810 5293 1818
rect 5308 1810 5321 1818
rect 5292 1802 5308 1810
rect 5289 1795 5308 1798
rect 5289 1786 5311 1795
rect 5262 1776 5311 1786
rect 5262 1770 5292 1776
rect 5311 1771 5316 1776
rect 5234 1754 5308 1770
rect 5326 1762 5356 1818
rect 5391 1808 5599 1818
rect 5634 1814 5679 1818
rect 5682 1817 5683 1818
rect 5698 1817 5711 1818
rect 5417 1778 5606 1808
rect 5432 1775 5606 1778
rect 5425 1772 5606 1775
rect 5234 1752 5247 1754
rect 5262 1752 5296 1754
rect 5234 1736 5308 1752
rect 5335 1748 5348 1762
rect 5363 1748 5379 1764
rect 5425 1759 5436 1772
rect 5218 1714 5219 1730
rect 5234 1714 5247 1736
rect 5262 1714 5292 1736
rect 5335 1732 5397 1748
rect 5425 1741 5436 1757
rect 5441 1752 5451 1772
rect 5461 1752 5475 1772
rect 5478 1759 5487 1772
rect 5503 1759 5512 1772
rect 5441 1741 5475 1752
rect 5478 1741 5487 1757
rect 5503 1741 5512 1757
rect 5519 1752 5529 1772
rect 5539 1752 5553 1772
rect 5554 1759 5565 1772
rect 5519 1741 5553 1752
rect 5554 1741 5565 1757
rect 5611 1748 5627 1764
rect 5634 1762 5664 1814
rect 5698 1810 5699 1817
rect 5683 1802 5699 1810
rect 5670 1770 5683 1789
rect 5698 1770 5728 1786
rect 5670 1754 5744 1770
rect 5670 1752 5683 1754
rect 5698 1752 5732 1754
rect 5335 1730 5348 1732
rect 5363 1730 5397 1732
rect 5335 1714 5397 1730
rect 5441 1725 5457 1732
rect 5519 1725 5549 1736
rect 5597 1732 5643 1748
rect 5670 1736 5744 1752
rect 5597 1730 5631 1732
rect 5596 1714 5643 1730
rect 5670 1714 5683 1736
rect 5698 1714 5728 1736
rect 5755 1714 5756 1730
rect 5771 1714 5784 1874
rect 5814 1770 5827 1874
rect 5872 1852 5873 1862
rect 5888 1852 5901 1862
rect 5872 1848 5901 1852
rect 5906 1848 5936 1874
rect 5954 1860 5970 1862
rect 6042 1860 6095 1874
rect 6043 1858 6107 1860
rect 6150 1858 6165 1874
rect 6214 1871 6244 1874
rect 6214 1868 6250 1871
rect 6180 1860 6196 1862
rect 5954 1848 5969 1852
rect 5872 1846 5969 1848
rect 5997 1846 6165 1858
rect 6181 1848 6196 1852
rect 6214 1849 6253 1868
rect 6272 1862 6279 1863
rect 6278 1855 6279 1862
rect 6262 1852 6263 1855
rect 6278 1852 6291 1855
rect 6214 1848 6244 1849
rect 6253 1848 6259 1849
rect 6262 1848 6291 1852
rect 6181 1847 6291 1848
rect 6181 1846 6297 1847
rect 5856 1838 5907 1846
rect 5856 1826 5881 1838
rect 5888 1826 5907 1838
rect 5938 1838 5988 1846
rect 5938 1830 5954 1838
rect 5961 1836 5988 1838
rect 5997 1836 6218 1846
rect 5961 1826 6218 1836
rect 6247 1838 6297 1846
rect 6247 1829 6263 1838
rect 5856 1818 5907 1826
rect 5954 1818 6218 1826
rect 6244 1826 6263 1829
rect 6270 1826 6297 1838
rect 6244 1818 6297 1826
rect 5872 1810 5873 1818
rect 5888 1810 5901 1818
rect 5872 1802 5888 1810
rect 5869 1795 5888 1798
rect 5869 1786 5891 1795
rect 5842 1776 5891 1786
rect 5842 1770 5872 1776
rect 5891 1771 5896 1776
rect 5814 1754 5888 1770
rect 5906 1762 5936 1818
rect 5971 1808 6179 1818
rect 6214 1814 6259 1818
rect 6262 1817 6263 1818
rect 6278 1817 6291 1818
rect 5997 1778 6186 1808
rect 6012 1775 6186 1778
rect 6005 1772 6186 1775
rect 5814 1752 5827 1754
rect 5842 1752 5876 1754
rect 5814 1736 5888 1752
rect 5915 1748 5928 1762
rect 5943 1748 5959 1764
rect 6005 1759 6016 1772
rect 5798 1714 5799 1730
rect 5814 1714 5827 1736
rect 5842 1714 5872 1736
rect 5915 1732 5977 1748
rect 6005 1741 6016 1757
rect 6021 1752 6031 1772
rect 6041 1752 6055 1772
rect 6058 1759 6067 1772
rect 6083 1759 6092 1772
rect 6021 1741 6055 1752
rect 6058 1741 6067 1757
rect 6083 1741 6092 1757
rect 6099 1752 6109 1772
rect 6119 1752 6133 1772
rect 6134 1759 6145 1772
rect 6099 1741 6133 1752
rect 6134 1741 6145 1757
rect 6191 1748 6207 1764
rect 6214 1762 6244 1814
rect 6278 1810 6279 1817
rect 6263 1802 6279 1810
rect 6250 1770 6263 1789
rect 6278 1770 6308 1786
rect 6250 1754 6324 1770
rect 6250 1752 6263 1754
rect 6278 1752 6312 1754
rect 5915 1730 5928 1732
rect 5943 1730 5977 1732
rect 5915 1714 5977 1730
rect 6021 1725 6037 1732
rect 6099 1725 6129 1736
rect 6177 1732 6223 1748
rect 6250 1736 6324 1752
rect 6177 1730 6211 1732
rect 6176 1714 6223 1730
rect 6250 1714 6263 1736
rect 6278 1714 6308 1736
rect 6335 1714 6336 1730
rect 6351 1714 6364 1874
rect 6394 1770 6407 1874
rect 6452 1852 6453 1862
rect 6468 1852 6481 1862
rect 6452 1848 6481 1852
rect 6486 1848 6516 1874
rect 6534 1860 6550 1862
rect 6622 1860 6675 1874
rect 6623 1858 6687 1860
rect 6730 1858 6745 1874
rect 6794 1871 6824 1874
rect 6794 1868 6830 1871
rect 6760 1860 6776 1862
rect 6534 1848 6549 1852
rect 6452 1846 6549 1848
rect 6577 1846 6745 1858
rect 6761 1848 6776 1852
rect 6794 1849 6833 1868
rect 6852 1862 6859 1863
rect 6858 1855 6859 1862
rect 6842 1852 6843 1855
rect 6858 1852 6871 1855
rect 6794 1848 6824 1849
rect 6833 1848 6839 1849
rect 6842 1848 6871 1852
rect 6761 1847 6871 1848
rect 6761 1846 6877 1847
rect 6436 1838 6487 1846
rect 6436 1826 6461 1838
rect 6468 1826 6487 1838
rect 6518 1838 6568 1846
rect 6518 1830 6534 1838
rect 6541 1836 6568 1838
rect 6577 1836 6798 1846
rect 6541 1826 6798 1836
rect 6827 1838 6877 1846
rect 6827 1829 6843 1838
rect 6436 1818 6487 1826
rect 6534 1818 6798 1826
rect 6824 1826 6843 1829
rect 6850 1826 6877 1838
rect 6824 1818 6877 1826
rect 6452 1810 6453 1818
rect 6468 1810 6481 1818
rect 6452 1802 6468 1810
rect 6449 1795 6468 1798
rect 6449 1786 6471 1795
rect 6422 1776 6471 1786
rect 6422 1770 6452 1776
rect 6471 1771 6476 1776
rect 6394 1754 6468 1770
rect 6486 1762 6516 1818
rect 6551 1808 6759 1818
rect 6794 1814 6839 1818
rect 6842 1817 6843 1818
rect 6858 1817 6871 1818
rect 6577 1778 6766 1808
rect 6592 1775 6766 1778
rect 6585 1772 6766 1775
rect 6394 1752 6407 1754
rect 6422 1752 6456 1754
rect 6394 1736 6468 1752
rect 6495 1748 6508 1762
rect 6523 1748 6539 1764
rect 6585 1759 6596 1772
rect 6378 1714 6379 1730
rect 6394 1714 6407 1736
rect 6422 1714 6452 1736
rect 6495 1732 6557 1748
rect 6585 1741 6596 1757
rect 6601 1752 6611 1772
rect 6621 1752 6635 1772
rect 6638 1759 6647 1772
rect 6663 1759 6672 1772
rect 6601 1741 6635 1752
rect 6638 1741 6647 1757
rect 6663 1741 6672 1757
rect 6679 1752 6689 1772
rect 6699 1752 6713 1772
rect 6714 1759 6725 1772
rect 6679 1741 6713 1752
rect 6714 1741 6725 1757
rect 6771 1748 6787 1764
rect 6794 1762 6824 1814
rect 6858 1810 6859 1817
rect 6843 1802 6859 1810
rect 6830 1770 6843 1789
rect 6858 1770 6888 1786
rect 6830 1754 6904 1770
rect 6830 1752 6843 1754
rect 6858 1752 6892 1754
rect 6495 1730 6508 1732
rect 6523 1730 6557 1732
rect 6495 1714 6557 1730
rect 6601 1725 6617 1732
rect 6679 1725 6709 1736
rect 6757 1732 6803 1748
rect 6830 1736 6904 1752
rect 6757 1730 6791 1732
rect 6756 1714 6803 1730
rect 6830 1714 6843 1736
rect 6858 1714 6888 1736
rect 6915 1714 6916 1730
rect 6931 1714 6944 1874
rect -8 1706 33 1714
rect -8 1680 7 1706
rect 14 1680 33 1706
rect 97 1702 159 1714
rect 171 1702 246 1714
rect 304 1702 379 1714
rect 391 1702 422 1714
rect 428 1702 463 1714
rect 97 1700 259 1702
rect -8 1672 33 1680
rect 115 1676 128 1700
rect 143 1698 158 1700
rect -2 1662 -1 1672
rect 14 1662 27 1672
rect 42 1662 72 1676
rect 115 1662 158 1676
rect 182 1673 189 1680
rect 192 1676 259 1700
rect 291 1700 463 1702
rect 261 1678 289 1682
rect 291 1678 371 1700
rect 392 1698 407 1700
rect 261 1676 371 1678
rect 192 1672 371 1676
rect 165 1662 195 1672
rect 197 1662 350 1672
rect 358 1662 388 1672
rect 392 1662 422 1676
rect 450 1662 463 1700
rect 535 1706 570 1714
rect 535 1680 536 1706
rect 543 1680 570 1706
rect 478 1662 508 1676
rect 535 1672 570 1680
rect 572 1706 613 1714
rect 572 1680 587 1706
rect 594 1680 613 1706
rect 677 1702 739 1714
rect 751 1702 826 1714
rect 884 1702 959 1714
rect 971 1702 1002 1714
rect 1008 1702 1043 1714
rect 677 1700 839 1702
rect 572 1672 613 1680
rect 695 1676 708 1700
rect 723 1698 738 1700
rect 535 1662 536 1672
rect 551 1662 564 1672
rect 578 1662 579 1672
rect 594 1662 607 1672
rect 622 1662 652 1676
rect 695 1662 738 1676
rect 762 1673 769 1680
rect 772 1676 839 1700
rect 871 1700 1043 1702
rect 841 1678 869 1682
rect 871 1678 951 1700
rect 972 1698 987 1700
rect 841 1676 951 1678
rect 772 1672 951 1676
rect 745 1662 775 1672
rect 777 1662 930 1672
rect 938 1662 968 1672
rect 972 1662 1002 1676
rect 1030 1662 1043 1700
rect 1115 1706 1150 1714
rect 1115 1680 1116 1706
rect 1123 1680 1150 1706
rect 1058 1662 1088 1676
rect 1115 1672 1150 1680
rect 1152 1706 1193 1714
rect 1152 1680 1167 1706
rect 1174 1680 1193 1706
rect 1257 1702 1319 1714
rect 1331 1702 1406 1714
rect 1464 1702 1539 1714
rect 1551 1702 1582 1714
rect 1588 1702 1623 1714
rect 1257 1700 1419 1702
rect 1152 1672 1193 1680
rect 1275 1676 1288 1700
rect 1303 1698 1318 1700
rect 1115 1662 1116 1672
rect 1131 1662 1144 1672
rect 1158 1662 1159 1672
rect 1174 1662 1187 1672
rect 1202 1662 1232 1676
rect 1275 1662 1318 1676
rect 1342 1673 1349 1680
rect 1352 1676 1419 1700
rect 1451 1700 1623 1702
rect 1421 1678 1449 1682
rect 1451 1678 1531 1700
rect 1552 1698 1567 1700
rect 1421 1676 1531 1678
rect 1352 1672 1531 1676
rect 1325 1662 1355 1672
rect 1357 1662 1510 1672
rect 1518 1662 1548 1672
rect 1552 1662 1582 1676
rect 1610 1662 1623 1700
rect 1695 1706 1730 1714
rect 1695 1680 1696 1706
rect 1703 1680 1730 1706
rect 1638 1662 1668 1676
rect 1695 1672 1730 1680
rect 1732 1706 1773 1714
rect 1732 1680 1747 1706
rect 1754 1680 1773 1706
rect 1732 1672 1773 1680
rect 3481 1706 3513 1714
rect 3481 1680 3487 1706
rect 3494 1680 3513 1706
rect 3577 1702 3639 1714
rect 3651 1702 3726 1714
rect 3784 1702 3859 1714
rect 3871 1702 3902 1714
rect 3908 1702 3943 1714
rect 3577 1700 3739 1702
rect 1695 1662 1696 1672
rect 1711 1662 1724 1672
rect 1738 1662 1739 1672
rect 1754 1662 1767 1672
rect 1782 1662 1812 1676
rect 3481 1672 3513 1680
rect 3595 1676 3608 1700
rect 3623 1698 3638 1700
rect 3494 1662 3507 1672
rect 3522 1662 3552 1676
rect 3595 1662 3638 1676
rect 3662 1673 3669 1680
rect 3672 1676 3739 1700
rect 3771 1700 3943 1702
rect 3741 1678 3769 1682
rect 3771 1678 3851 1700
rect 3872 1698 3887 1700
rect 3741 1676 3851 1678
rect 3672 1672 3851 1676
rect 3645 1662 3675 1672
rect 3677 1662 3830 1672
rect 3838 1662 3868 1672
rect 3872 1662 3902 1676
rect 3930 1662 3943 1700
rect 4015 1706 4050 1714
rect 4015 1680 4016 1706
rect 4023 1680 4050 1706
rect 3958 1662 3988 1676
rect 4015 1672 4050 1680
rect 4052 1706 4093 1714
rect 4052 1680 4067 1706
rect 4074 1680 4093 1706
rect 4157 1702 4219 1714
rect 4231 1702 4306 1714
rect 4364 1702 4439 1714
rect 4451 1702 4482 1714
rect 4488 1702 4523 1714
rect 4157 1700 4319 1702
rect 4052 1672 4093 1680
rect 4175 1676 4188 1700
rect 4203 1698 4218 1700
rect 4015 1662 4016 1672
rect 4031 1662 4044 1672
rect 4058 1662 4059 1672
rect 4074 1662 4087 1672
rect 4102 1662 4132 1676
rect 4175 1662 4218 1676
rect 4242 1673 4249 1680
rect 4252 1676 4319 1700
rect 4351 1700 4523 1702
rect 4321 1678 4349 1682
rect 4351 1678 4431 1700
rect 4452 1698 4467 1700
rect 4321 1676 4431 1678
rect 4252 1672 4431 1676
rect 4225 1662 4255 1672
rect 4257 1662 4410 1672
rect 4418 1662 4448 1672
rect 4452 1662 4482 1676
rect 4510 1662 4523 1700
rect 4595 1706 4630 1714
rect 4595 1680 4596 1706
rect 4603 1680 4630 1706
rect 4538 1662 4568 1676
rect 4595 1672 4630 1680
rect 4632 1706 4673 1714
rect 4632 1680 4647 1706
rect 4654 1680 4673 1706
rect 4737 1702 4799 1714
rect 4811 1702 4886 1714
rect 4944 1702 5019 1714
rect 5031 1702 5062 1714
rect 5068 1702 5103 1714
rect 4737 1700 4899 1702
rect 4755 1682 4768 1700
rect 4783 1698 4798 1700
rect 4632 1672 4673 1680
rect 4756 1676 4768 1682
rect 4595 1662 4596 1672
rect 4611 1662 4624 1672
rect 4638 1662 4639 1672
rect 4654 1662 4667 1672
rect 4682 1662 4712 1676
rect 4756 1662 4798 1676
rect 4822 1673 4829 1680
rect 4832 1676 4899 1700
rect 4931 1700 5103 1702
rect 4901 1678 4929 1682
rect 4931 1678 5011 1700
rect 5032 1698 5047 1700
rect 4901 1676 5011 1678
rect 4832 1672 5011 1676
rect 4805 1662 4835 1672
rect 4837 1662 4990 1672
rect 4998 1662 5028 1672
rect 5032 1662 5062 1676
rect 5090 1662 5103 1700
rect 5175 1706 5210 1714
rect 5175 1680 5176 1706
rect 5183 1680 5210 1706
rect 5118 1662 5148 1676
rect 5175 1672 5210 1680
rect 5212 1706 5253 1714
rect 5212 1680 5227 1706
rect 5234 1680 5253 1706
rect 5317 1702 5379 1714
rect 5391 1702 5466 1714
rect 5524 1702 5599 1714
rect 5611 1702 5642 1714
rect 5648 1702 5683 1714
rect 5317 1700 5479 1702
rect 5335 1682 5348 1700
rect 5363 1698 5378 1700
rect 5212 1672 5253 1680
rect 5336 1676 5348 1682
rect 5175 1662 5176 1672
rect 5191 1662 5204 1672
rect 5218 1662 5219 1672
rect 5234 1662 5247 1672
rect 5262 1662 5292 1676
rect 5336 1662 5378 1676
rect 5402 1673 5409 1680
rect 5412 1676 5479 1700
rect 5511 1700 5683 1702
rect 5481 1678 5509 1682
rect 5511 1678 5591 1700
rect 5612 1698 5627 1700
rect 5481 1676 5591 1678
rect 5412 1672 5591 1676
rect 5385 1662 5415 1672
rect 5417 1662 5570 1672
rect 5578 1662 5608 1672
rect 5612 1662 5642 1676
rect 5670 1662 5683 1700
rect 5755 1706 5790 1714
rect 5755 1680 5756 1706
rect 5763 1680 5790 1706
rect 5698 1662 5728 1676
rect 5755 1672 5790 1680
rect 5792 1706 5833 1714
rect 5792 1680 5807 1706
rect 5814 1680 5833 1706
rect 5897 1702 5959 1714
rect 5971 1702 6046 1714
rect 6104 1702 6179 1714
rect 6191 1702 6222 1714
rect 6228 1702 6263 1714
rect 5897 1700 6059 1702
rect 5915 1682 5928 1700
rect 5943 1698 5958 1700
rect 5792 1672 5833 1680
rect 5916 1676 5928 1682
rect 5755 1662 5756 1672
rect 5771 1662 5784 1672
rect 5798 1662 5799 1672
rect 5814 1662 5827 1672
rect 5842 1662 5872 1676
rect 5916 1662 5958 1676
rect 5982 1673 5989 1680
rect 5992 1676 6059 1700
rect 6091 1700 6263 1702
rect 6061 1678 6089 1682
rect 6091 1678 6171 1700
rect 6192 1698 6207 1700
rect 6061 1676 6171 1678
rect 5992 1672 6171 1676
rect 5965 1662 5995 1672
rect 5997 1662 6150 1672
rect 6158 1662 6188 1672
rect 6192 1662 6222 1676
rect 6250 1662 6263 1700
rect 6335 1706 6370 1714
rect 6335 1680 6336 1706
rect 6343 1680 6370 1706
rect 6278 1662 6308 1676
rect 6335 1672 6370 1680
rect 6372 1706 6413 1714
rect 6372 1680 6387 1706
rect 6394 1680 6413 1706
rect 6477 1702 6539 1714
rect 6551 1702 6626 1714
rect 6684 1702 6759 1714
rect 6771 1702 6802 1714
rect 6808 1702 6843 1714
rect 6477 1700 6639 1702
rect 6495 1682 6508 1700
rect 6523 1698 6538 1700
rect 6372 1672 6413 1680
rect 6496 1676 6508 1682
rect 6335 1662 6336 1672
rect 6351 1662 6364 1672
rect 6378 1662 6379 1672
rect 6394 1662 6407 1672
rect 6422 1662 6452 1676
rect 6496 1662 6538 1676
rect 6562 1673 6569 1680
rect 6572 1676 6639 1700
rect 6671 1700 6843 1702
rect 6641 1678 6669 1682
rect 6671 1678 6751 1700
rect 6772 1698 6787 1700
rect 6641 1676 6751 1678
rect 6572 1672 6751 1676
rect 6545 1662 6575 1672
rect 6577 1662 6730 1672
rect 6738 1662 6768 1672
rect 6772 1662 6802 1676
rect 6830 1662 6843 1700
rect 6915 1706 6950 1714
rect 6915 1680 6916 1706
rect 6923 1680 6950 1706
rect 6858 1662 6888 1676
rect 6915 1672 6950 1680
rect 6915 1662 6916 1672
rect 6931 1662 6944 1672
rect -2 1656 1837 1662
rect -1 1648 1837 1656
rect 3481 1648 6944 1662
rect 14 1618 27 1648
rect 42 1630 72 1648
rect 115 1634 129 1648
rect 165 1634 385 1648
rect 116 1632 129 1634
rect 82 1620 97 1632
rect 79 1618 101 1620
rect 106 1618 136 1632
rect 197 1630 350 1634
rect 179 1618 371 1630
rect 414 1618 444 1632
rect 450 1618 463 1648
rect 478 1630 508 1648
rect 551 1618 564 1648
rect 594 1618 607 1648
rect 622 1630 652 1648
rect 695 1634 709 1648
rect 745 1634 965 1648
rect 696 1632 709 1634
rect 662 1620 677 1632
rect 659 1618 681 1620
rect 686 1618 716 1632
rect 777 1630 930 1634
rect 759 1618 951 1630
rect 994 1618 1024 1632
rect 1030 1618 1043 1648
rect 1058 1630 1088 1648
rect 1131 1618 1144 1648
rect 1174 1618 1187 1648
rect 1202 1630 1232 1648
rect 1275 1634 1289 1648
rect 1325 1634 1545 1648
rect 1276 1632 1289 1634
rect 1242 1620 1257 1632
rect 1239 1618 1261 1620
rect 1266 1618 1296 1632
rect 1357 1630 1510 1634
rect 1339 1618 1531 1630
rect 1574 1618 1604 1632
rect 1610 1618 1623 1648
rect 1638 1630 1668 1648
rect 1711 1618 1724 1648
rect 1754 1618 1767 1648
rect 1782 1630 1812 1648
rect 1822 1620 1837 1632
rect 1819 1618 1837 1620
rect 3494 1618 3507 1648
rect 3522 1630 3552 1648
rect 3595 1634 3609 1648
rect 3645 1634 3865 1648
rect 3596 1632 3609 1634
rect 3562 1620 3577 1632
rect 3559 1618 3581 1620
rect 3586 1618 3616 1632
rect 3677 1630 3830 1634
rect 3659 1618 3851 1630
rect 3894 1618 3924 1632
rect 3930 1618 3943 1648
rect 3958 1630 3988 1648
rect 4031 1618 4044 1648
rect 4074 1618 4087 1648
rect 4102 1630 4132 1648
rect 4175 1634 4189 1648
rect 4225 1634 4445 1648
rect 4176 1632 4189 1634
rect 4142 1620 4157 1632
rect 4139 1618 4161 1620
rect 4166 1618 4196 1632
rect 4257 1630 4410 1634
rect 4239 1618 4431 1630
rect 4474 1618 4504 1632
rect 4510 1618 4523 1648
rect 4538 1630 4568 1648
rect 4611 1618 4624 1648
rect 4654 1618 4667 1648
rect 4682 1630 4712 1648
rect 4756 1632 4769 1648
rect 4805 1634 5025 1648
rect 4722 1620 4737 1632
rect 4719 1618 4741 1620
rect 4746 1618 4776 1632
rect 4837 1630 4990 1634
rect 4819 1618 5011 1630
rect 5054 1618 5084 1632
rect 5090 1618 5103 1648
rect 5118 1630 5148 1648
rect 5191 1618 5204 1648
rect 5234 1618 5247 1648
rect 5262 1630 5292 1648
rect 5336 1632 5349 1648
rect 5385 1634 5605 1648
rect 5302 1620 5317 1632
rect 5299 1618 5321 1620
rect 5326 1618 5356 1632
rect 5417 1630 5570 1634
rect 5399 1618 5591 1630
rect 5634 1618 5664 1632
rect 5670 1618 5683 1648
rect 5698 1630 5728 1648
rect 5771 1618 5784 1648
rect 5814 1618 5827 1648
rect 5842 1630 5872 1648
rect 5916 1632 5929 1648
rect 5965 1634 6185 1648
rect 5882 1620 5897 1632
rect 5879 1618 5901 1620
rect 5906 1618 5936 1632
rect 5997 1630 6150 1634
rect 5979 1618 6171 1630
rect 6214 1618 6244 1632
rect 6250 1618 6263 1648
rect 6278 1630 6308 1648
rect 6351 1618 6364 1648
rect 6394 1618 6407 1648
rect 6422 1630 6452 1648
rect 6496 1632 6509 1648
rect 6545 1634 6765 1648
rect 6462 1620 6477 1632
rect 6459 1618 6481 1620
rect 6486 1618 6516 1632
rect 6577 1630 6730 1634
rect 6559 1618 6751 1630
rect 6794 1618 6824 1632
rect 6830 1618 6843 1648
rect 6858 1630 6888 1648
rect 6931 1618 6944 1648
rect -1 1604 1837 1618
rect 3481 1604 6944 1618
rect 14 1500 27 1604
rect 72 1582 73 1592
rect 88 1582 101 1592
rect 72 1578 101 1582
rect 106 1578 136 1604
rect 154 1590 170 1592
rect 242 1590 295 1604
rect 243 1588 307 1590
rect 350 1588 365 1604
rect 414 1601 444 1604
rect 414 1598 450 1601
rect 380 1590 396 1592
rect 154 1578 169 1582
rect 72 1576 169 1578
rect 197 1576 365 1588
rect 381 1578 396 1582
rect 414 1579 453 1598
rect 472 1592 479 1593
rect 478 1585 479 1592
rect 462 1582 463 1585
rect 478 1582 491 1585
rect 414 1578 444 1579
rect 453 1578 459 1579
rect 462 1578 491 1582
rect 381 1577 491 1578
rect 381 1576 497 1577
rect 56 1568 107 1576
rect 56 1556 81 1568
rect 88 1556 107 1568
rect 138 1568 188 1576
rect 138 1560 154 1568
rect 161 1566 188 1568
rect 197 1566 418 1576
rect 161 1556 418 1566
rect 447 1568 497 1576
rect 447 1559 463 1568
rect 56 1548 107 1556
rect 154 1548 418 1556
rect 444 1556 463 1559
rect 470 1556 497 1568
rect 444 1548 497 1556
rect 72 1540 73 1548
rect 88 1540 101 1548
rect 72 1532 88 1540
rect 69 1525 88 1528
rect 69 1516 91 1525
rect 42 1506 91 1516
rect 42 1500 72 1506
rect 91 1501 96 1506
rect 14 1484 88 1500
rect 106 1492 136 1548
rect 171 1538 379 1548
rect 414 1544 459 1548
rect 462 1547 463 1548
rect 478 1547 491 1548
rect 197 1508 386 1538
rect 212 1505 386 1508
rect 205 1502 386 1505
rect 14 1482 27 1484
rect 42 1482 76 1484
rect 14 1466 88 1482
rect 115 1478 128 1492
rect 143 1478 159 1494
rect 205 1489 216 1502
rect -2 1444 -1 1460
rect 14 1444 27 1466
rect 42 1444 72 1466
rect 115 1462 177 1478
rect 205 1471 216 1487
rect 221 1482 231 1502
rect 241 1482 255 1502
rect 258 1489 267 1502
rect 283 1489 292 1502
rect 221 1471 255 1482
rect 258 1471 267 1487
rect 283 1471 292 1487
rect 299 1482 309 1502
rect 319 1482 333 1502
rect 334 1489 345 1502
rect 299 1471 333 1482
rect 334 1471 345 1487
rect 391 1478 407 1494
rect 414 1492 444 1544
rect 478 1540 479 1547
rect 463 1532 479 1540
rect 450 1500 463 1519
rect 478 1500 508 1516
rect 450 1484 524 1500
rect 450 1482 463 1484
rect 478 1482 512 1484
rect 115 1460 128 1462
rect 143 1460 177 1462
rect 115 1444 177 1460
rect 221 1455 237 1462
rect 299 1455 329 1466
rect 377 1462 423 1478
rect 450 1466 524 1482
rect 377 1460 411 1462
rect 376 1444 423 1460
rect 450 1444 463 1466
rect 478 1444 508 1466
rect 535 1444 536 1460
rect 551 1444 564 1604
rect 594 1500 607 1604
rect 652 1582 653 1592
rect 668 1582 681 1592
rect 652 1578 681 1582
rect 686 1578 716 1604
rect 734 1590 750 1592
rect 822 1590 875 1604
rect 823 1588 887 1590
rect 930 1588 945 1604
rect 994 1601 1024 1604
rect 994 1598 1030 1601
rect 960 1590 976 1592
rect 734 1578 749 1582
rect 652 1576 749 1578
rect 777 1576 945 1588
rect 961 1578 976 1582
rect 994 1579 1033 1598
rect 1052 1592 1059 1593
rect 1058 1585 1059 1592
rect 1042 1582 1043 1585
rect 1058 1582 1071 1585
rect 994 1578 1024 1579
rect 1033 1578 1039 1579
rect 1042 1578 1071 1582
rect 961 1577 1071 1578
rect 961 1576 1077 1577
rect 636 1568 687 1576
rect 636 1556 661 1568
rect 668 1556 687 1568
rect 718 1568 768 1576
rect 718 1560 734 1568
rect 741 1566 768 1568
rect 777 1566 998 1576
rect 741 1556 998 1566
rect 1027 1568 1077 1576
rect 1027 1559 1043 1568
rect 636 1548 687 1556
rect 734 1548 998 1556
rect 1024 1556 1043 1559
rect 1050 1556 1077 1568
rect 1024 1548 1077 1556
rect 652 1540 653 1548
rect 668 1540 681 1548
rect 652 1532 668 1540
rect 649 1525 668 1528
rect 649 1516 671 1525
rect 622 1506 671 1516
rect 622 1500 652 1506
rect 671 1501 676 1506
rect 594 1484 668 1500
rect 686 1492 716 1548
rect 751 1538 959 1548
rect 994 1544 1039 1548
rect 1042 1547 1043 1548
rect 1058 1547 1071 1548
rect 777 1508 966 1538
rect 792 1505 966 1508
rect 785 1502 966 1505
rect 594 1482 607 1484
rect 622 1482 656 1484
rect 594 1466 668 1482
rect 695 1478 708 1492
rect 723 1478 739 1494
rect 785 1489 796 1502
rect 578 1444 579 1460
rect 594 1444 607 1466
rect 622 1444 652 1466
rect 695 1462 757 1478
rect 785 1471 796 1487
rect 801 1482 811 1502
rect 821 1482 835 1502
rect 838 1489 847 1502
rect 863 1489 872 1502
rect 801 1471 835 1482
rect 838 1471 847 1487
rect 863 1471 872 1487
rect 879 1482 889 1502
rect 899 1482 913 1502
rect 914 1489 925 1502
rect 879 1471 913 1482
rect 914 1471 925 1487
rect 971 1478 987 1494
rect 994 1492 1024 1544
rect 1058 1540 1059 1547
rect 1043 1532 1059 1540
rect 1030 1500 1043 1519
rect 1058 1500 1088 1516
rect 1030 1484 1104 1500
rect 1030 1482 1043 1484
rect 1058 1482 1092 1484
rect 695 1460 708 1462
rect 723 1460 757 1462
rect 695 1444 757 1460
rect 801 1455 817 1462
rect 879 1455 909 1466
rect 957 1462 1003 1478
rect 1030 1466 1104 1482
rect 957 1460 991 1462
rect 956 1444 1003 1460
rect 1030 1444 1043 1466
rect 1058 1444 1088 1466
rect 1115 1444 1116 1460
rect 1131 1444 1144 1604
rect 1174 1500 1187 1604
rect 1232 1582 1233 1592
rect 1248 1582 1261 1592
rect 1232 1578 1261 1582
rect 1266 1578 1296 1604
rect 1314 1590 1330 1592
rect 1402 1590 1455 1604
rect 1403 1588 1467 1590
rect 1510 1588 1525 1604
rect 1574 1601 1604 1604
rect 1574 1598 1610 1601
rect 1540 1590 1556 1592
rect 1314 1578 1329 1582
rect 1232 1576 1329 1578
rect 1357 1576 1525 1588
rect 1541 1578 1556 1582
rect 1574 1579 1613 1598
rect 1632 1592 1639 1593
rect 1638 1585 1639 1592
rect 1622 1582 1623 1585
rect 1638 1582 1651 1585
rect 1574 1578 1604 1579
rect 1613 1578 1619 1579
rect 1622 1578 1651 1582
rect 1541 1577 1651 1578
rect 1541 1576 1657 1577
rect 1216 1568 1267 1576
rect 1216 1556 1241 1568
rect 1248 1556 1267 1568
rect 1298 1568 1348 1576
rect 1298 1560 1314 1568
rect 1321 1566 1348 1568
rect 1357 1566 1578 1576
rect 1321 1556 1578 1566
rect 1607 1568 1657 1576
rect 1607 1559 1623 1568
rect 1216 1548 1267 1556
rect 1314 1548 1578 1556
rect 1604 1556 1623 1559
rect 1630 1556 1657 1568
rect 1604 1548 1657 1556
rect 1232 1540 1233 1548
rect 1248 1540 1261 1548
rect 1232 1532 1248 1540
rect 1229 1525 1248 1528
rect 1229 1516 1251 1525
rect 1202 1506 1251 1516
rect 1202 1500 1232 1506
rect 1251 1501 1256 1506
rect 1174 1484 1248 1500
rect 1266 1492 1296 1548
rect 1331 1538 1539 1548
rect 1574 1544 1619 1548
rect 1622 1547 1623 1548
rect 1638 1547 1651 1548
rect 1357 1508 1546 1538
rect 1372 1505 1546 1508
rect 1365 1502 1546 1505
rect 1174 1482 1187 1484
rect 1202 1482 1236 1484
rect 1174 1466 1248 1482
rect 1275 1478 1288 1492
rect 1303 1478 1319 1494
rect 1365 1489 1376 1502
rect 1158 1444 1159 1460
rect 1174 1444 1187 1466
rect 1202 1444 1232 1466
rect 1275 1462 1337 1478
rect 1365 1471 1376 1487
rect 1381 1482 1391 1502
rect 1401 1482 1415 1502
rect 1418 1489 1427 1502
rect 1443 1489 1452 1502
rect 1381 1471 1415 1482
rect 1418 1471 1427 1487
rect 1443 1471 1452 1487
rect 1459 1482 1469 1502
rect 1479 1482 1493 1502
rect 1494 1489 1505 1502
rect 1459 1471 1493 1482
rect 1494 1471 1505 1487
rect 1551 1478 1567 1494
rect 1574 1492 1604 1544
rect 1638 1540 1639 1547
rect 1623 1532 1639 1540
rect 1610 1500 1623 1519
rect 1638 1500 1668 1516
rect 1610 1484 1684 1500
rect 1610 1482 1623 1484
rect 1638 1482 1672 1484
rect 1275 1460 1288 1462
rect 1303 1460 1337 1462
rect 1275 1444 1337 1460
rect 1381 1455 1397 1462
rect 1459 1455 1489 1466
rect 1537 1462 1583 1478
rect 1610 1466 1684 1482
rect 1537 1460 1571 1462
rect 1536 1444 1583 1460
rect 1610 1444 1623 1466
rect 1638 1444 1668 1466
rect 1695 1444 1696 1460
rect 1711 1444 1724 1604
rect 1754 1500 1767 1604
rect 1812 1582 1813 1592
rect 1828 1582 1837 1592
rect 1812 1576 1837 1582
rect 1796 1568 1837 1576
rect 1796 1556 1821 1568
rect 1828 1556 1837 1568
rect 1796 1548 1837 1556
rect 1812 1540 1813 1548
rect 1828 1540 1837 1548
rect 1812 1532 1828 1540
rect 1809 1525 1828 1528
rect 1809 1516 1831 1525
rect 1782 1506 1831 1516
rect 1782 1500 1812 1506
rect 1831 1501 1836 1506
rect 3494 1500 3507 1604
rect 3552 1582 3553 1592
rect 3568 1582 3581 1592
rect 3552 1578 3581 1582
rect 3586 1578 3616 1604
rect 3634 1590 3650 1592
rect 3722 1590 3775 1604
rect 3723 1588 3787 1590
rect 3830 1588 3845 1604
rect 3894 1601 3924 1604
rect 3894 1598 3930 1601
rect 3860 1590 3876 1592
rect 3634 1578 3649 1582
rect 3552 1576 3649 1578
rect 3677 1576 3845 1588
rect 3861 1578 3876 1582
rect 3894 1579 3933 1598
rect 3952 1592 3959 1593
rect 3958 1585 3959 1592
rect 3942 1582 3943 1585
rect 3958 1582 3971 1585
rect 3894 1578 3924 1579
rect 3933 1578 3939 1579
rect 3942 1578 3971 1582
rect 3861 1577 3971 1578
rect 3861 1576 3977 1577
rect 3536 1568 3587 1576
rect 3536 1556 3561 1568
rect 3568 1556 3587 1568
rect 3618 1568 3668 1576
rect 3618 1560 3634 1568
rect 3641 1566 3668 1568
rect 3677 1566 3898 1576
rect 3641 1556 3898 1566
rect 3927 1568 3977 1576
rect 3927 1559 3943 1568
rect 3536 1548 3587 1556
rect 3634 1548 3898 1556
rect 3924 1556 3943 1559
rect 3950 1556 3977 1568
rect 3924 1548 3977 1556
rect 3552 1540 3553 1548
rect 3568 1540 3581 1548
rect 3552 1532 3568 1540
rect 3549 1525 3568 1528
rect 3549 1516 3571 1525
rect 3522 1506 3571 1516
rect 3522 1500 3552 1506
rect 3571 1501 3576 1506
rect 1754 1484 1828 1500
rect 3494 1484 3568 1500
rect 3586 1492 3616 1548
rect 3651 1538 3859 1548
rect 3894 1544 3939 1548
rect 3942 1547 3943 1548
rect 3958 1547 3971 1548
rect 3677 1508 3866 1538
rect 3692 1505 3866 1508
rect 3685 1502 3866 1505
rect 1754 1482 1767 1484
rect 1782 1482 1816 1484
rect 3494 1482 3507 1484
rect 3522 1482 3556 1484
rect 1754 1466 1828 1482
rect 3494 1466 3568 1482
rect 3595 1478 3608 1492
rect 3623 1478 3639 1494
rect 3685 1489 3696 1502
rect 1738 1444 1739 1460
rect 1754 1444 1767 1466
rect 1782 1444 1812 1466
rect 3494 1444 3507 1466
rect 3522 1444 3552 1466
rect 3595 1462 3657 1478
rect 3685 1471 3696 1487
rect 3701 1482 3711 1502
rect 3721 1482 3735 1502
rect 3738 1489 3747 1502
rect 3763 1489 3772 1502
rect 3701 1471 3735 1482
rect 3738 1471 3747 1487
rect 3763 1471 3772 1487
rect 3779 1482 3789 1502
rect 3799 1482 3813 1502
rect 3814 1489 3825 1502
rect 3779 1471 3813 1482
rect 3814 1471 3825 1487
rect 3871 1478 3887 1494
rect 3894 1492 3924 1544
rect 3958 1540 3959 1547
rect 3943 1532 3959 1540
rect 3930 1500 3943 1519
rect 3958 1500 3988 1516
rect 3930 1484 4004 1500
rect 3930 1482 3943 1484
rect 3958 1482 3992 1484
rect 3595 1460 3608 1462
rect 3623 1460 3657 1462
rect 3595 1444 3657 1460
rect 3701 1455 3717 1462
rect 3779 1455 3809 1466
rect 3857 1462 3903 1478
rect 3930 1466 4004 1482
rect 3857 1460 3891 1462
rect 3856 1444 3903 1460
rect 3930 1444 3943 1466
rect 3958 1444 3988 1466
rect 4015 1444 4016 1460
rect 4031 1444 4044 1604
rect 4074 1500 4087 1604
rect 4132 1582 4133 1592
rect 4148 1582 4161 1592
rect 4132 1578 4161 1582
rect 4166 1578 4196 1604
rect 4214 1590 4230 1592
rect 4302 1590 4355 1604
rect 4303 1588 4367 1590
rect 4410 1588 4425 1604
rect 4474 1601 4504 1604
rect 4474 1598 4510 1601
rect 4440 1590 4456 1592
rect 4214 1578 4229 1582
rect 4132 1576 4229 1578
rect 4257 1576 4425 1588
rect 4441 1578 4456 1582
rect 4474 1579 4513 1598
rect 4532 1592 4539 1593
rect 4538 1585 4539 1592
rect 4522 1582 4523 1585
rect 4538 1582 4551 1585
rect 4474 1578 4504 1579
rect 4513 1578 4519 1579
rect 4522 1578 4551 1582
rect 4441 1577 4551 1578
rect 4441 1576 4557 1577
rect 4116 1568 4167 1576
rect 4116 1556 4141 1568
rect 4148 1556 4167 1568
rect 4198 1568 4248 1576
rect 4198 1560 4214 1568
rect 4221 1566 4248 1568
rect 4257 1566 4478 1576
rect 4221 1556 4478 1566
rect 4507 1568 4557 1576
rect 4507 1559 4523 1568
rect 4116 1548 4167 1556
rect 4214 1548 4478 1556
rect 4504 1556 4523 1559
rect 4530 1556 4557 1568
rect 4504 1548 4557 1556
rect 4132 1540 4133 1548
rect 4148 1540 4161 1548
rect 4132 1532 4148 1540
rect 4129 1525 4148 1528
rect 4129 1516 4151 1525
rect 4102 1506 4151 1516
rect 4102 1500 4132 1506
rect 4151 1501 4156 1506
rect 4074 1484 4148 1500
rect 4166 1492 4196 1548
rect 4231 1538 4439 1548
rect 4474 1544 4519 1548
rect 4522 1547 4523 1548
rect 4538 1547 4551 1548
rect 4257 1508 4446 1538
rect 4272 1505 4446 1508
rect 4265 1502 4446 1505
rect 4074 1482 4087 1484
rect 4102 1482 4136 1484
rect 4074 1466 4148 1482
rect 4175 1478 4188 1492
rect 4203 1478 4219 1494
rect 4265 1489 4276 1502
rect 4058 1444 4059 1460
rect 4074 1444 4087 1466
rect 4102 1444 4132 1466
rect 4175 1462 4237 1478
rect 4265 1471 4276 1487
rect 4281 1482 4291 1502
rect 4301 1482 4315 1502
rect 4318 1489 4327 1502
rect 4343 1489 4352 1502
rect 4281 1471 4315 1482
rect 4318 1471 4327 1487
rect 4343 1471 4352 1487
rect 4359 1482 4369 1502
rect 4379 1482 4393 1502
rect 4394 1489 4405 1502
rect 4359 1471 4393 1482
rect 4394 1471 4405 1487
rect 4451 1478 4467 1494
rect 4474 1492 4504 1544
rect 4538 1540 4539 1547
rect 4523 1532 4539 1540
rect 4510 1500 4523 1519
rect 4538 1500 4568 1516
rect 4510 1484 4584 1500
rect 4510 1482 4523 1484
rect 4538 1482 4572 1484
rect 4175 1460 4188 1462
rect 4203 1460 4237 1462
rect 4175 1444 4237 1460
rect 4281 1455 4297 1462
rect 4359 1455 4389 1466
rect 4437 1462 4483 1478
rect 4510 1466 4584 1482
rect 4437 1460 4471 1462
rect 4436 1444 4483 1460
rect 4510 1444 4523 1466
rect 4538 1444 4568 1466
rect 4595 1444 4596 1460
rect 4611 1444 4624 1604
rect 4654 1500 4667 1604
rect 4712 1582 4713 1592
rect 4728 1582 4741 1592
rect 4712 1578 4741 1582
rect 4746 1578 4776 1604
rect 4794 1590 4810 1592
rect 4882 1590 4935 1604
rect 4883 1588 4947 1590
rect 4990 1588 5005 1604
rect 5054 1601 5084 1604
rect 5054 1598 5090 1601
rect 5020 1590 5036 1592
rect 4794 1578 4809 1582
rect 4712 1576 4809 1578
rect 4837 1576 5005 1588
rect 5021 1578 5036 1582
rect 5054 1579 5093 1598
rect 5112 1592 5119 1593
rect 5118 1585 5119 1592
rect 5102 1582 5103 1585
rect 5118 1582 5131 1585
rect 5054 1578 5084 1579
rect 5093 1578 5099 1579
rect 5102 1578 5131 1582
rect 5021 1577 5131 1578
rect 5021 1576 5137 1577
rect 4696 1568 4747 1576
rect 4696 1556 4721 1568
rect 4728 1556 4747 1568
rect 4778 1568 4828 1576
rect 4778 1560 4794 1568
rect 4801 1566 4828 1568
rect 4837 1566 5058 1576
rect 4801 1556 5058 1566
rect 5087 1568 5137 1576
rect 5087 1559 5103 1568
rect 4696 1548 4747 1556
rect 4794 1548 5058 1556
rect 5084 1556 5103 1559
rect 5110 1556 5137 1568
rect 5084 1548 5137 1556
rect 4712 1540 4713 1548
rect 4728 1540 4741 1548
rect 4712 1532 4728 1540
rect 4709 1525 4728 1528
rect 4709 1516 4731 1525
rect 4682 1506 4731 1516
rect 4682 1500 4712 1506
rect 4731 1501 4736 1506
rect 4654 1484 4728 1500
rect 4746 1492 4776 1548
rect 4811 1538 5019 1548
rect 5054 1544 5099 1548
rect 5102 1547 5103 1548
rect 5118 1547 5131 1548
rect 4837 1508 5026 1538
rect 4852 1505 5026 1508
rect 4845 1502 5026 1505
rect 4654 1482 4667 1484
rect 4682 1482 4716 1484
rect 4654 1466 4728 1482
rect 4755 1478 4768 1492
rect 4783 1478 4799 1494
rect 4845 1489 4856 1502
rect 4638 1444 4639 1460
rect 4654 1444 4667 1466
rect 4682 1444 4712 1466
rect 4755 1462 4817 1478
rect 4845 1471 4856 1487
rect 4861 1482 4871 1502
rect 4881 1482 4895 1502
rect 4898 1489 4907 1502
rect 4923 1489 4932 1502
rect 4861 1471 4895 1482
rect 4898 1471 4907 1487
rect 4923 1471 4932 1487
rect 4939 1482 4949 1502
rect 4959 1482 4973 1502
rect 4974 1489 4985 1502
rect 4939 1471 4973 1482
rect 4974 1471 4985 1487
rect 5031 1478 5047 1494
rect 5054 1492 5084 1544
rect 5118 1540 5119 1547
rect 5103 1532 5119 1540
rect 5090 1500 5103 1519
rect 5118 1500 5148 1516
rect 5090 1484 5164 1500
rect 5090 1482 5103 1484
rect 5118 1482 5152 1484
rect 4755 1460 4768 1462
rect 4783 1460 4817 1462
rect 4755 1444 4817 1460
rect 4861 1455 4877 1462
rect 4939 1455 4969 1466
rect 5017 1462 5063 1478
rect 5090 1466 5164 1482
rect 5017 1460 5051 1462
rect 5016 1444 5063 1460
rect 5090 1444 5103 1466
rect 5118 1444 5148 1466
rect 5175 1444 5176 1460
rect 5191 1444 5204 1604
rect 5234 1500 5247 1604
rect 5292 1582 5293 1592
rect 5308 1582 5321 1592
rect 5292 1578 5321 1582
rect 5326 1578 5356 1604
rect 5374 1590 5390 1592
rect 5462 1590 5515 1604
rect 5463 1588 5527 1590
rect 5570 1588 5585 1604
rect 5634 1601 5664 1604
rect 5634 1598 5670 1601
rect 5600 1590 5616 1592
rect 5374 1578 5389 1582
rect 5292 1576 5389 1578
rect 5417 1576 5585 1588
rect 5601 1578 5616 1582
rect 5634 1579 5673 1598
rect 5692 1592 5699 1593
rect 5698 1585 5699 1592
rect 5682 1582 5683 1585
rect 5698 1582 5711 1585
rect 5634 1578 5664 1579
rect 5673 1578 5679 1579
rect 5682 1578 5711 1582
rect 5601 1577 5711 1578
rect 5601 1576 5717 1577
rect 5276 1568 5327 1576
rect 5276 1556 5301 1568
rect 5308 1556 5327 1568
rect 5358 1568 5408 1576
rect 5358 1560 5374 1568
rect 5381 1566 5408 1568
rect 5417 1566 5638 1576
rect 5381 1556 5638 1566
rect 5667 1568 5717 1576
rect 5667 1559 5683 1568
rect 5276 1548 5327 1556
rect 5374 1548 5638 1556
rect 5664 1556 5683 1559
rect 5690 1556 5717 1568
rect 5664 1548 5717 1556
rect 5292 1540 5293 1548
rect 5308 1540 5321 1548
rect 5292 1532 5308 1540
rect 5289 1525 5308 1528
rect 5289 1516 5311 1525
rect 5262 1506 5311 1516
rect 5262 1500 5292 1506
rect 5311 1501 5316 1506
rect 5234 1484 5308 1500
rect 5326 1492 5356 1548
rect 5391 1538 5599 1548
rect 5634 1544 5679 1548
rect 5682 1547 5683 1548
rect 5698 1547 5711 1548
rect 5417 1508 5606 1538
rect 5432 1505 5606 1508
rect 5425 1502 5606 1505
rect 5234 1482 5247 1484
rect 5262 1482 5296 1484
rect 5234 1466 5308 1482
rect 5335 1478 5348 1492
rect 5363 1478 5379 1494
rect 5425 1489 5436 1502
rect 5218 1444 5219 1460
rect 5234 1444 5247 1466
rect 5262 1444 5292 1466
rect 5335 1462 5397 1478
rect 5425 1471 5436 1487
rect 5441 1482 5451 1502
rect 5461 1482 5475 1502
rect 5478 1489 5487 1502
rect 5503 1489 5512 1502
rect 5441 1471 5475 1482
rect 5478 1471 5487 1487
rect 5503 1471 5512 1487
rect 5519 1482 5529 1502
rect 5539 1482 5553 1502
rect 5554 1489 5565 1502
rect 5519 1471 5553 1482
rect 5554 1471 5565 1487
rect 5611 1478 5627 1494
rect 5634 1492 5664 1544
rect 5698 1540 5699 1547
rect 5683 1532 5699 1540
rect 5670 1500 5683 1519
rect 5698 1500 5728 1516
rect 5670 1484 5744 1500
rect 5670 1482 5683 1484
rect 5698 1482 5732 1484
rect 5335 1460 5348 1462
rect 5363 1460 5397 1462
rect 5335 1444 5397 1460
rect 5441 1455 5457 1462
rect 5519 1455 5549 1466
rect 5597 1462 5643 1478
rect 5670 1466 5744 1482
rect 5597 1460 5631 1462
rect 5596 1444 5643 1460
rect 5670 1444 5683 1466
rect 5698 1444 5728 1466
rect 5755 1444 5756 1460
rect 5771 1444 5784 1604
rect 5814 1500 5827 1604
rect 5872 1582 5873 1592
rect 5888 1582 5901 1592
rect 5872 1578 5901 1582
rect 5906 1578 5936 1604
rect 5954 1590 5970 1592
rect 6042 1590 6095 1604
rect 6043 1588 6107 1590
rect 6150 1588 6165 1604
rect 6214 1601 6244 1604
rect 6214 1598 6250 1601
rect 6180 1590 6196 1592
rect 5954 1578 5969 1582
rect 5872 1576 5969 1578
rect 5997 1576 6165 1588
rect 6181 1578 6196 1582
rect 6214 1579 6253 1598
rect 6272 1592 6279 1593
rect 6278 1585 6279 1592
rect 6262 1582 6263 1585
rect 6278 1582 6291 1585
rect 6214 1578 6244 1579
rect 6253 1578 6259 1579
rect 6262 1578 6291 1582
rect 6181 1577 6291 1578
rect 6181 1576 6297 1577
rect 5856 1568 5907 1576
rect 5856 1556 5881 1568
rect 5888 1556 5907 1568
rect 5938 1568 5988 1576
rect 5938 1560 5954 1568
rect 5961 1566 5988 1568
rect 5997 1566 6218 1576
rect 5961 1556 6218 1566
rect 6247 1568 6297 1576
rect 6247 1559 6263 1568
rect 5856 1548 5907 1556
rect 5954 1548 6218 1556
rect 6244 1556 6263 1559
rect 6270 1556 6297 1568
rect 6244 1548 6297 1556
rect 5872 1540 5873 1548
rect 5888 1540 5901 1548
rect 5872 1532 5888 1540
rect 5869 1525 5888 1528
rect 5869 1516 5891 1525
rect 5842 1506 5891 1516
rect 5842 1500 5872 1506
rect 5891 1501 5896 1506
rect 5814 1484 5888 1500
rect 5906 1492 5936 1548
rect 5971 1538 6179 1548
rect 6214 1544 6259 1548
rect 6262 1547 6263 1548
rect 6278 1547 6291 1548
rect 5997 1508 6186 1538
rect 6012 1505 6186 1508
rect 6005 1502 6186 1505
rect 5814 1482 5827 1484
rect 5842 1482 5876 1484
rect 5814 1466 5888 1482
rect 5915 1478 5928 1492
rect 5943 1478 5959 1494
rect 6005 1489 6016 1502
rect 5798 1444 5799 1460
rect 5814 1444 5827 1466
rect 5842 1444 5872 1466
rect 5915 1462 5977 1478
rect 6005 1471 6016 1487
rect 6021 1482 6031 1502
rect 6041 1482 6055 1502
rect 6058 1489 6067 1502
rect 6083 1489 6092 1502
rect 6021 1471 6055 1482
rect 6058 1471 6067 1487
rect 6083 1471 6092 1487
rect 6099 1482 6109 1502
rect 6119 1482 6133 1502
rect 6134 1489 6145 1502
rect 6099 1471 6133 1482
rect 6134 1471 6145 1487
rect 6191 1478 6207 1494
rect 6214 1492 6244 1544
rect 6278 1540 6279 1547
rect 6263 1532 6279 1540
rect 6250 1500 6263 1519
rect 6278 1500 6308 1516
rect 6250 1484 6324 1500
rect 6250 1482 6263 1484
rect 6278 1482 6312 1484
rect 5915 1460 5928 1462
rect 5943 1460 5977 1462
rect 5915 1444 5977 1460
rect 6021 1455 6037 1462
rect 6099 1455 6129 1466
rect 6177 1462 6223 1478
rect 6250 1466 6324 1482
rect 6177 1460 6211 1462
rect 6176 1444 6223 1460
rect 6250 1444 6263 1466
rect 6278 1444 6308 1466
rect 6335 1444 6336 1460
rect 6351 1444 6364 1604
rect 6394 1500 6407 1604
rect 6452 1582 6453 1592
rect 6468 1582 6481 1592
rect 6452 1578 6481 1582
rect 6486 1578 6516 1604
rect 6534 1590 6550 1592
rect 6622 1590 6675 1604
rect 6623 1588 6687 1590
rect 6730 1588 6745 1604
rect 6794 1601 6824 1604
rect 6794 1598 6830 1601
rect 6760 1590 6776 1592
rect 6534 1578 6549 1582
rect 6452 1576 6549 1578
rect 6577 1576 6745 1588
rect 6761 1578 6776 1582
rect 6794 1579 6833 1598
rect 6852 1592 6859 1593
rect 6858 1585 6859 1592
rect 6842 1582 6843 1585
rect 6858 1582 6871 1585
rect 6794 1578 6824 1579
rect 6833 1578 6839 1579
rect 6842 1578 6871 1582
rect 6761 1577 6871 1578
rect 6761 1576 6877 1577
rect 6436 1568 6487 1576
rect 6436 1556 6461 1568
rect 6468 1556 6487 1568
rect 6518 1568 6568 1576
rect 6518 1560 6534 1568
rect 6541 1566 6568 1568
rect 6577 1566 6798 1576
rect 6541 1556 6798 1566
rect 6827 1568 6877 1576
rect 6827 1559 6843 1568
rect 6436 1548 6487 1556
rect 6534 1548 6798 1556
rect 6824 1556 6843 1559
rect 6850 1556 6877 1568
rect 6824 1548 6877 1556
rect 6452 1540 6453 1548
rect 6468 1540 6481 1548
rect 6452 1532 6468 1540
rect 6449 1525 6468 1528
rect 6449 1516 6471 1525
rect 6422 1506 6471 1516
rect 6422 1500 6452 1506
rect 6471 1501 6476 1506
rect 6394 1484 6468 1500
rect 6486 1492 6516 1548
rect 6551 1538 6759 1548
rect 6794 1544 6839 1548
rect 6842 1547 6843 1548
rect 6858 1547 6871 1548
rect 6577 1508 6766 1538
rect 6592 1505 6766 1508
rect 6585 1502 6766 1505
rect 6394 1482 6407 1484
rect 6422 1482 6456 1484
rect 6394 1466 6468 1482
rect 6495 1478 6508 1492
rect 6523 1478 6539 1494
rect 6585 1489 6596 1502
rect 6378 1444 6379 1460
rect 6394 1444 6407 1466
rect 6422 1444 6452 1466
rect 6495 1462 6557 1478
rect 6585 1471 6596 1487
rect 6601 1482 6611 1502
rect 6621 1482 6635 1502
rect 6638 1489 6647 1502
rect 6663 1489 6672 1502
rect 6601 1471 6635 1482
rect 6638 1471 6647 1487
rect 6663 1471 6672 1487
rect 6679 1482 6689 1502
rect 6699 1482 6713 1502
rect 6714 1489 6725 1502
rect 6679 1471 6713 1482
rect 6714 1471 6725 1487
rect 6771 1478 6787 1494
rect 6794 1492 6824 1544
rect 6858 1540 6859 1547
rect 6843 1532 6859 1540
rect 6830 1500 6843 1519
rect 6858 1500 6888 1516
rect 6830 1484 6904 1500
rect 6830 1482 6843 1484
rect 6858 1482 6892 1484
rect 6495 1460 6508 1462
rect 6523 1460 6557 1462
rect 6495 1444 6557 1460
rect 6601 1455 6617 1462
rect 6679 1455 6709 1466
rect 6757 1462 6803 1478
rect 6830 1466 6904 1482
rect 6757 1460 6791 1462
rect 6756 1444 6803 1460
rect 6830 1444 6843 1466
rect 6858 1444 6888 1466
rect 6915 1444 6916 1460
rect 6931 1444 6944 1604
rect -8 1436 33 1444
rect -8 1410 7 1436
rect 14 1410 33 1436
rect 97 1432 159 1444
rect 171 1432 246 1444
rect 304 1432 379 1444
rect 391 1432 422 1444
rect 428 1432 463 1444
rect 97 1430 259 1432
rect -8 1402 33 1410
rect 115 1406 128 1430
rect 143 1428 158 1430
rect -2 1392 -1 1402
rect 14 1392 27 1402
rect 42 1392 72 1406
rect 115 1392 158 1406
rect 182 1403 189 1410
rect 192 1406 259 1430
rect 291 1430 463 1432
rect 261 1408 289 1412
rect 291 1408 371 1430
rect 392 1428 407 1430
rect 261 1406 371 1408
rect 192 1402 371 1406
rect 165 1392 195 1402
rect 197 1392 350 1402
rect 358 1392 388 1402
rect 392 1392 422 1406
rect 450 1392 463 1430
rect 535 1436 570 1444
rect 535 1410 536 1436
rect 543 1410 570 1436
rect 478 1392 508 1406
rect 535 1402 570 1410
rect 572 1436 613 1444
rect 572 1410 587 1436
rect 594 1410 613 1436
rect 677 1432 739 1444
rect 751 1432 826 1444
rect 884 1432 959 1444
rect 971 1432 1002 1444
rect 1008 1432 1043 1444
rect 677 1430 839 1432
rect 572 1402 613 1410
rect 695 1406 708 1430
rect 723 1428 738 1430
rect 535 1392 536 1402
rect 551 1392 564 1402
rect 578 1392 579 1402
rect 594 1392 607 1402
rect 622 1392 652 1406
rect 695 1392 738 1406
rect 762 1403 769 1410
rect 772 1406 839 1430
rect 871 1430 1043 1432
rect 841 1408 869 1412
rect 871 1408 951 1430
rect 972 1428 987 1430
rect 841 1406 951 1408
rect 772 1402 951 1406
rect 745 1392 775 1402
rect 777 1392 930 1402
rect 938 1392 968 1402
rect 972 1392 1002 1406
rect 1030 1392 1043 1430
rect 1115 1436 1150 1444
rect 1115 1410 1116 1436
rect 1123 1410 1150 1436
rect 1058 1392 1088 1406
rect 1115 1402 1150 1410
rect 1152 1436 1193 1444
rect 1152 1410 1167 1436
rect 1174 1410 1193 1436
rect 1257 1432 1319 1444
rect 1331 1432 1406 1444
rect 1464 1432 1539 1444
rect 1551 1432 1582 1444
rect 1588 1432 1623 1444
rect 1257 1430 1419 1432
rect 1152 1402 1193 1410
rect 1275 1406 1288 1430
rect 1303 1428 1318 1430
rect 1115 1392 1116 1402
rect 1131 1392 1144 1402
rect 1158 1392 1159 1402
rect 1174 1392 1187 1402
rect 1202 1392 1232 1406
rect 1275 1392 1318 1406
rect 1342 1403 1349 1410
rect 1352 1406 1419 1430
rect 1451 1430 1623 1432
rect 1421 1408 1449 1412
rect 1451 1408 1531 1430
rect 1552 1428 1567 1430
rect 1421 1406 1531 1408
rect 1352 1402 1531 1406
rect 1325 1392 1355 1402
rect 1357 1392 1510 1402
rect 1518 1392 1548 1402
rect 1552 1392 1582 1406
rect 1610 1392 1623 1430
rect 1695 1436 1730 1444
rect 1695 1410 1696 1436
rect 1703 1410 1730 1436
rect 1638 1392 1668 1406
rect 1695 1402 1730 1410
rect 1732 1436 1773 1444
rect 1732 1410 1747 1436
rect 1754 1410 1773 1436
rect 1732 1402 1773 1410
rect 3481 1436 3513 1444
rect 3481 1410 3487 1436
rect 3494 1410 3513 1436
rect 3577 1432 3639 1444
rect 3651 1432 3726 1444
rect 3784 1432 3859 1444
rect 3871 1432 3902 1444
rect 3908 1432 3943 1444
rect 3577 1430 3739 1432
rect 1695 1392 1696 1402
rect 1711 1392 1724 1402
rect 1738 1392 1739 1402
rect 1754 1392 1767 1402
rect 1782 1392 1812 1406
rect 3481 1402 3513 1410
rect 3595 1406 3608 1430
rect 3623 1428 3638 1430
rect 3494 1392 3507 1402
rect 3522 1392 3552 1406
rect 3595 1392 3638 1406
rect 3662 1403 3669 1410
rect 3672 1406 3739 1430
rect 3771 1430 3943 1432
rect 3741 1408 3769 1412
rect 3771 1408 3851 1430
rect 3872 1428 3887 1430
rect 3741 1406 3851 1408
rect 3672 1402 3851 1406
rect 3645 1392 3675 1402
rect 3677 1392 3830 1402
rect 3838 1392 3868 1402
rect 3872 1392 3902 1406
rect 3930 1392 3943 1430
rect 4015 1436 4050 1444
rect 4015 1410 4016 1436
rect 4023 1410 4050 1436
rect 3958 1392 3988 1406
rect 4015 1402 4050 1410
rect 4052 1436 4093 1444
rect 4052 1410 4067 1436
rect 4074 1410 4093 1436
rect 4157 1432 4219 1444
rect 4231 1432 4306 1444
rect 4364 1432 4439 1444
rect 4451 1432 4482 1444
rect 4488 1432 4523 1444
rect 4157 1430 4319 1432
rect 4052 1402 4093 1410
rect 4175 1406 4188 1430
rect 4203 1428 4218 1430
rect 4015 1392 4016 1402
rect 4031 1392 4044 1402
rect 4058 1392 4059 1402
rect 4074 1392 4087 1402
rect 4102 1392 4132 1406
rect 4175 1392 4218 1406
rect 4242 1403 4249 1410
rect 4252 1406 4319 1430
rect 4351 1430 4523 1432
rect 4321 1408 4349 1412
rect 4351 1408 4431 1430
rect 4452 1428 4467 1430
rect 4321 1406 4431 1408
rect 4252 1402 4431 1406
rect 4225 1392 4255 1402
rect 4257 1392 4410 1402
rect 4418 1392 4448 1402
rect 4452 1392 4482 1406
rect 4510 1392 4523 1430
rect 4595 1436 4630 1444
rect 4595 1410 4596 1436
rect 4603 1410 4630 1436
rect 4538 1392 4568 1406
rect 4595 1402 4630 1410
rect 4632 1436 4673 1444
rect 4632 1410 4647 1436
rect 4654 1410 4673 1436
rect 4737 1432 4799 1444
rect 4811 1432 4886 1444
rect 4944 1432 5019 1444
rect 5031 1432 5062 1444
rect 5068 1432 5103 1444
rect 4737 1430 4899 1432
rect 4632 1402 4673 1410
rect 4755 1406 4768 1430
rect 4783 1428 4798 1430
rect 4595 1392 4596 1402
rect 4611 1392 4624 1402
rect 4638 1392 4639 1402
rect 4654 1392 4667 1402
rect 4682 1392 4712 1406
rect 4755 1392 4798 1406
rect 4822 1403 4829 1410
rect 4832 1406 4899 1430
rect 4931 1430 5103 1432
rect 4901 1408 4929 1412
rect 4931 1408 5011 1430
rect 5032 1428 5047 1430
rect 4901 1406 5011 1408
rect 4832 1402 5011 1406
rect 4805 1392 4835 1402
rect 4837 1392 4990 1402
rect 4998 1392 5028 1402
rect 5032 1392 5062 1406
rect 5090 1392 5103 1430
rect 5175 1436 5210 1444
rect 5175 1410 5176 1436
rect 5183 1410 5210 1436
rect 5118 1392 5148 1406
rect 5175 1402 5210 1410
rect 5212 1436 5253 1444
rect 5212 1410 5227 1436
rect 5234 1410 5253 1436
rect 5317 1432 5379 1444
rect 5391 1432 5466 1444
rect 5524 1432 5599 1444
rect 5611 1432 5642 1444
rect 5648 1432 5683 1444
rect 5317 1430 5479 1432
rect 5212 1402 5253 1410
rect 5335 1406 5348 1430
rect 5363 1428 5378 1430
rect 5175 1392 5176 1402
rect 5191 1392 5204 1402
rect 5218 1392 5219 1402
rect 5234 1392 5247 1402
rect 5262 1392 5292 1406
rect 5335 1392 5378 1406
rect 5402 1403 5409 1410
rect 5412 1406 5479 1430
rect 5511 1430 5683 1432
rect 5481 1408 5509 1412
rect 5511 1408 5591 1430
rect 5612 1428 5627 1430
rect 5481 1406 5591 1408
rect 5412 1402 5591 1406
rect 5385 1392 5415 1402
rect 5417 1392 5570 1402
rect 5578 1392 5608 1402
rect 5612 1392 5642 1406
rect 5670 1392 5683 1430
rect 5755 1436 5790 1444
rect 5755 1410 5756 1436
rect 5763 1410 5790 1436
rect 5698 1392 5728 1406
rect 5755 1402 5790 1410
rect 5792 1436 5833 1444
rect 5792 1410 5807 1436
rect 5814 1410 5833 1436
rect 5897 1432 5959 1444
rect 5971 1432 6046 1444
rect 6104 1432 6179 1444
rect 6191 1432 6222 1444
rect 6228 1432 6263 1444
rect 5897 1430 6059 1432
rect 5792 1402 5833 1410
rect 5915 1406 5928 1430
rect 5943 1428 5958 1430
rect 5755 1392 5756 1402
rect 5771 1392 5784 1402
rect 5798 1392 5799 1402
rect 5814 1392 5827 1402
rect 5842 1392 5872 1406
rect 5915 1392 5958 1406
rect 5982 1403 5989 1410
rect 5992 1406 6059 1430
rect 6091 1430 6263 1432
rect 6061 1408 6089 1412
rect 6091 1408 6171 1430
rect 6192 1428 6207 1430
rect 6061 1406 6171 1408
rect 5992 1402 6171 1406
rect 5965 1392 5995 1402
rect 5997 1392 6150 1402
rect 6158 1392 6188 1402
rect 6192 1392 6222 1406
rect 6250 1392 6263 1430
rect 6335 1436 6370 1444
rect 6335 1410 6336 1436
rect 6343 1410 6370 1436
rect 6278 1392 6308 1406
rect 6335 1402 6370 1410
rect 6372 1436 6413 1444
rect 6372 1410 6387 1436
rect 6394 1410 6413 1436
rect 6477 1432 6539 1444
rect 6551 1432 6626 1444
rect 6684 1432 6759 1444
rect 6771 1432 6802 1444
rect 6808 1432 6843 1444
rect 6477 1430 6639 1432
rect 6372 1402 6413 1410
rect 6495 1406 6508 1430
rect 6523 1428 6538 1430
rect 6335 1392 6336 1402
rect 6351 1392 6364 1402
rect 6378 1392 6379 1402
rect 6394 1392 6407 1402
rect 6422 1392 6452 1406
rect 6495 1392 6538 1406
rect 6562 1403 6569 1410
rect 6572 1406 6639 1430
rect 6671 1430 6843 1432
rect 6641 1408 6669 1412
rect 6671 1408 6751 1430
rect 6772 1428 6787 1430
rect 6641 1406 6751 1408
rect 6572 1402 6751 1406
rect 6545 1392 6575 1402
rect 6577 1392 6730 1402
rect 6738 1392 6768 1402
rect 6772 1392 6802 1406
rect 6830 1392 6843 1430
rect 6915 1436 6950 1444
rect 6915 1410 6916 1436
rect 6923 1410 6950 1436
rect 6858 1392 6888 1406
rect 6915 1402 6950 1410
rect 6915 1392 6916 1402
rect 6931 1392 6944 1402
rect -2 1386 1837 1392
rect -1 1378 1837 1386
rect 3481 1378 6944 1392
rect 14 1348 27 1378
rect 42 1360 72 1378
rect 115 1364 129 1378
rect 165 1364 385 1378
rect 116 1362 129 1364
rect 82 1350 97 1362
rect 79 1348 101 1350
rect 106 1348 136 1362
rect 197 1360 350 1364
rect 179 1348 371 1360
rect 414 1348 444 1362
rect 450 1348 463 1378
rect 478 1360 508 1378
rect 551 1348 564 1378
rect 594 1348 607 1378
rect 622 1360 652 1378
rect 695 1364 709 1378
rect 745 1364 965 1378
rect 696 1362 709 1364
rect 662 1350 677 1362
rect 659 1348 681 1350
rect 686 1348 716 1362
rect 777 1360 930 1364
rect 759 1348 951 1360
rect 994 1348 1024 1362
rect 1030 1348 1043 1378
rect 1058 1360 1088 1378
rect 1131 1348 1144 1378
rect 1174 1348 1187 1378
rect 1202 1360 1232 1378
rect 1275 1364 1289 1378
rect 1325 1364 1545 1378
rect 1276 1362 1289 1364
rect 1242 1350 1257 1362
rect 1239 1348 1261 1350
rect 1266 1348 1296 1362
rect 1357 1360 1510 1364
rect 1339 1348 1531 1360
rect 1574 1348 1604 1362
rect 1610 1348 1623 1378
rect 1638 1360 1668 1378
rect 1711 1348 1724 1378
rect 1754 1348 1767 1378
rect 1782 1360 1812 1378
rect 1822 1350 1837 1362
rect 1819 1348 1837 1350
rect 3494 1348 3507 1378
rect 3522 1360 3552 1378
rect 3595 1364 3609 1378
rect 3645 1364 3865 1378
rect 3596 1362 3609 1364
rect 3562 1350 3577 1362
rect 3559 1348 3581 1350
rect 3586 1348 3616 1362
rect 3677 1360 3830 1364
rect 3659 1348 3851 1360
rect 3894 1348 3924 1362
rect 3930 1348 3943 1378
rect 3958 1360 3988 1378
rect 4031 1348 4044 1378
rect 4074 1348 4087 1378
rect 4102 1360 4132 1378
rect 4175 1364 4189 1378
rect 4225 1364 4445 1378
rect 4176 1362 4189 1364
rect 4142 1350 4157 1362
rect 4139 1348 4161 1350
rect 4166 1348 4196 1362
rect 4257 1360 4410 1364
rect 4239 1348 4431 1360
rect 4474 1348 4504 1362
rect 4510 1348 4523 1378
rect 4538 1360 4568 1378
rect 4611 1348 4624 1378
rect 4654 1348 4667 1378
rect 4682 1360 4712 1378
rect 4755 1364 4769 1378
rect 4805 1364 5025 1378
rect 4756 1362 4769 1364
rect 4722 1350 4737 1362
rect 4719 1348 4741 1350
rect 4746 1348 4776 1362
rect 4837 1360 4990 1364
rect 4819 1348 5011 1360
rect 5054 1348 5084 1362
rect 5090 1348 5103 1378
rect 5118 1360 5148 1378
rect 5191 1348 5204 1378
rect 5234 1348 5247 1378
rect 5262 1360 5292 1378
rect 5335 1364 5349 1378
rect 5385 1364 5605 1378
rect 5336 1362 5349 1364
rect 5302 1350 5317 1362
rect 5299 1348 5321 1350
rect 5326 1348 5356 1362
rect 5417 1360 5570 1364
rect 5399 1348 5591 1360
rect 5634 1348 5664 1362
rect 5670 1348 5683 1378
rect 5698 1360 5728 1378
rect 5771 1348 5784 1378
rect 5814 1348 5827 1378
rect 5842 1360 5872 1378
rect 5915 1364 5929 1378
rect 5965 1364 6185 1378
rect 5916 1362 5929 1364
rect 5882 1350 5897 1362
rect 5879 1348 5901 1350
rect 5906 1348 5936 1362
rect 5997 1360 6150 1364
rect 5979 1348 6171 1360
rect 6214 1348 6244 1362
rect 6250 1348 6263 1378
rect 6278 1360 6308 1378
rect 6351 1348 6364 1378
rect 6394 1348 6407 1378
rect 6422 1360 6452 1378
rect 6495 1364 6509 1378
rect 6545 1364 6765 1378
rect 6496 1362 6509 1364
rect 6462 1350 6477 1362
rect 6459 1348 6481 1350
rect 6486 1348 6516 1362
rect 6577 1360 6730 1364
rect 6559 1348 6751 1360
rect 6794 1348 6824 1362
rect 6830 1348 6843 1378
rect 6858 1360 6888 1378
rect 6931 1348 6944 1378
rect -1 1334 1837 1348
rect 3481 1334 6944 1348
rect 14 1230 27 1334
rect 72 1312 73 1322
rect 88 1312 101 1322
rect 72 1308 101 1312
rect 106 1308 136 1334
rect 154 1320 170 1322
rect 242 1320 295 1334
rect 243 1318 307 1320
rect 350 1318 365 1334
rect 414 1331 444 1334
rect 414 1328 450 1331
rect 380 1320 396 1322
rect 154 1308 169 1312
rect 72 1306 169 1308
rect 197 1306 365 1318
rect 381 1308 396 1312
rect 414 1309 453 1328
rect 472 1322 479 1323
rect 478 1315 479 1322
rect 462 1312 463 1315
rect 478 1312 491 1315
rect 414 1308 444 1309
rect 453 1308 459 1309
rect 462 1308 491 1312
rect 381 1307 491 1308
rect 381 1306 497 1307
rect 56 1298 107 1306
rect 56 1286 81 1298
rect 88 1286 107 1298
rect 138 1298 188 1306
rect 138 1290 154 1298
rect 161 1296 188 1298
rect 197 1296 418 1306
rect 161 1286 418 1296
rect 447 1298 497 1306
rect 447 1289 463 1298
rect 56 1278 107 1286
rect 154 1278 418 1286
rect 444 1286 463 1289
rect 470 1286 497 1298
rect 444 1278 497 1286
rect 72 1270 73 1278
rect 88 1270 101 1278
rect 72 1262 88 1270
rect 69 1255 88 1258
rect 69 1246 91 1255
rect 42 1236 91 1246
rect 42 1230 72 1236
rect 91 1231 96 1236
rect 14 1214 88 1230
rect 106 1222 136 1278
rect 171 1268 379 1278
rect 414 1274 459 1278
rect 462 1277 463 1278
rect 478 1277 491 1278
rect 197 1238 386 1268
rect 212 1235 386 1238
rect 205 1232 386 1235
rect 14 1212 27 1214
rect 42 1212 76 1214
rect 14 1196 88 1212
rect 115 1208 128 1222
rect 143 1208 159 1224
rect 205 1219 216 1232
rect -2 1174 -1 1190
rect 14 1174 27 1196
rect 42 1174 72 1196
rect 115 1192 177 1208
rect 205 1201 216 1217
rect 221 1212 231 1232
rect 241 1212 255 1232
rect 258 1219 267 1232
rect 283 1219 292 1232
rect 221 1201 255 1212
rect 258 1201 267 1217
rect 283 1201 292 1217
rect 299 1212 309 1232
rect 319 1212 333 1232
rect 334 1219 345 1232
rect 299 1201 333 1212
rect 334 1201 345 1217
rect 391 1208 407 1224
rect 414 1222 444 1274
rect 478 1270 479 1277
rect 463 1262 479 1270
rect 450 1230 463 1249
rect 478 1230 508 1246
rect 450 1214 524 1230
rect 450 1212 463 1214
rect 478 1212 512 1214
rect 115 1190 128 1192
rect 143 1190 177 1192
rect 115 1174 177 1190
rect 221 1185 237 1192
rect 299 1185 329 1196
rect 377 1192 423 1208
rect 450 1196 524 1212
rect 377 1190 411 1192
rect 376 1174 423 1190
rect 450 1174 463 1196
rect 478 1174 508 1196
rect 535 1174 536 1190
rect 551 1174 564 1334
rect 594 1230 607 1334
rect 652 1312 653 1322
rect 668 1312 681 1322
rect 652 1308 681 1312
rect 686 1308 716 1334
rect 734 1320 750 1322
rect 822 1320 875 1334
rect 823 1318 887 1320
rect 930 1318 945 1334
rect 994 1331 1024 1334
rect 994 1328 1030 1331
rect 960 1320 976 1322
rect 734 1308 749 1312
rect 652 1306 749 1308
rect 777 1306 945 1318
rect 961 1308 976 1312
rect 994 1309 1033 1328
rect 1052 1322 1059 1323
rect 1058 1315 1059 1322
rect 1042 1312 1043 1315
rect 1058 1312 1071 1315
rect 994 1308 1024 1309
rect 1033 1308 1039 1309
rect 1042 1308 1071 1312
rect 961 1307 1071 1308
rect 961 1306 1077 1307
rect 636 1298 687 1306
rect 636 1286 661 1298
rect 668 1286 687 1298
rect 718 1298 768 1306
rect 718 1290 734 1298
rect 741 1296 768 1298
rect 777 1296 998 1306
rect 741 1286 998 1296
rect 1027 1298 1077 1306
rect 1027 1289 1043 1298
rect 636 1278 687 1286
rect 734 1278 998 1286
rect 1024 1286 1043 1289
rect 1050 1286 1077 1298
rect 1024 1278 1077 1286
rect 652 1270 653 1278
rect 668 1270 681 1278
rect 652 1262 668 1270
rect 649 1255 668 1258
rect 649 1246 671 1255
rect 622 1236 671 1246
rect 622 1230 652 1236
rect 671 1231 676 1236
rect 594 1214 668 1230
rect 686 1222 716 1278
rect 751 1268 959 1278
rect 994 1274 1039 1278
rect 1042 1277 1043 1278
rect 1058 1277 1071 1278
rect 777 1238 966 1268
rect 792 1235 966 1238
rect 785 1232 966 1235
rect 594 1212 607 1214
rect 622 1212 656 1214
rect 594 1196 668 1212
rect 695 1208 708 1222
rect 723 1208 739 1224
rect 785 1219 796 1232
rect 578 1174 579 1190
rect 594 1174 607 1196
rect 622 1174 652 1196
rect 695 1192 757 1208
rect 785 1201 796 1217
rect 801 1212 811 1232
rect 821 1212 835 1232
rect 838 1219 847 1232
rect 863 1219 872 1232
rect 801 1201 835 1212
rect 838 1201 847 1217
rect 863 1201 872 1217
rect 879 1212 889 1232
rect 899 1212 913 1232
rect 914 1219 925 1232
rect 879 1201 913 1212
rect 914 1201 925 1217
rect 971 1208 987 1224
rect 994 1222 1024 1274
rect 1058 1270 1059 1277
rect 1043 1262 1059 1270
rect 1030 1230 1043 1249
rect 1058 1230 1088 1246
rect 1030 1214 1104 1230
rect 1030 1212 1043 1214
rect 1058 1212 1092 1214
rect 695 1190 708 1192
rect 723 1190 757 1192
rect 695 1174 757 1190
rect 801 1185 817 1192
rect 879 1185 909 1196
rect 957 1192 1003 1208
rect 1030 1196 1104 1212
rect 957 1190 991 1192
rect 956 1174 1003 1190
rect 1030 1174 1043 1196
rect 1058 1174 1088 1196
rect 1115 1174 1116 1190
rect 1131 1174 1144 1334
rect 1174 1230 1187 1334
rect 1232 1312 1233 1322
rect 1248 1312 1261 1322
rect 1232 1308 1261 1312
rect 1266 1308 1296 1334
rect 1314 1320 1330 1322
rect 1402 1320 1455 1334
rect 1403 1318 1467 1320
rect 1510 1318 1525 1334
rect 1574 1331 1604 1334
rect 1574 1328 1610 1331
rect 1540 1320 1556 1322
rect 1314 1308 1329 1312
rect 1232 1306 1329 1308
rect 1357 1306 1525 1318
rect 1541 1308 1556 1312
rect 1574 1309 1613 1328
rect 1632 1322 1639 1323
rect 1638 1315 1639 1322
rect 1622 1312 1623 1315
rect 1638 1312 1651 1315
rect 1574 1308 1604 1309
rect 1613 1308 1619 1309
rect 1622 1308 1651 1312
rect 1541 1307 1651 1308
rect 1541 1306 1657 1307
rect 1216 1298 1267 1306
rect 1216 1286 1241 1298
rect 1248 1286 1267 1298
rect 1298 1298 1348 1306
rect 1298 1290 1314 1298
rect 1321 1296 1348 1298
rect 1357 1296 1578 1306
rect 1321 1286 1578 1296
rect 1607 1298 1657 1306
rect 1607 1289 1623 1298
rect 1216 1278 1267 1286
rect 1314 1278 1578 1286
rect 1604 1286 1623 1289
rect 1630 1286 1657 1298
rect 1604 1278 1657 1286
rect 1232 1270 1233 1278
rect 1248 1270 1261 1278
rect 1232 1262 1248 1270
rect 1229 1255 1248 1258
rect 1229 1246 1251 1255
rect 1202 1236 1251 1246
rect 1202 1230 1232 1236
rect 1251 1231 1256 1236
rect 1174 1214 1248 1230
rect 1266 1222 1296 1278
rect 1331 1268 1539 1278
rect 1574 1274 1619 1278
rect 1622 1277 1623 1278
rect 1638 1277 1651 1278
rect 1357 1238 1546 1268
rect 1372 1235 1546 1238
rect 1365 1232 1546 1235
rect 1174 1212 1187 1214
rect 1202 1212 1236 1214
rect 1174 1196 1248 1212
rect 1275 1208 1288 1222
rect 1303 1208 1319 1224
rect 1365 1219 1376 1232
rect 1158 1174 1159 1190
rect 1174 1174 1187 1196
rect 1202 1174 1232 1196
rect 1275 1192 1337 1208
rect 1365 1201 1376 1217
rect 1381 1212 1391 1232
rect 1401 1212 1415 1232
rect 1418 1219 1427 1232
rect 1443 1219 1452 1232
rect 1381 1201 1415 1212
rect 1418 1201 1427 1217
rect 1443 1201 1452 1217
rect 1459 1212 1469 1232
rect 1479 1212 1493 1232
rect 1494 1219 1505 1232
rect 1459 1201 1493 1212
rect 1494 1201 1505 1217
rect 1551 1208 1567 1224
rect 1574 1222 1604 1274
rect 1638 1270 1639 1277
rect 1623 1262 1639 1270
rect 1610 1230 1623 1249
rect 1638 1230 1668 1246
rect 1610 1214 1684 1230
rect 1610 1212 1623 1214
rect 1638 1212 1672 1214
rect 1275 1190 1288 1192
rect 1303 1190 1337 1192
rect 1275 1174 1337 1190
rect 1381 1185 1397 1192
rect 1459 1185 1489 1196
rect 1537 1192 1583 1208
rect 1610 1196 1684 1212
rect 1537 1190 1571 1192
rect 1536 1174 1583 1190
rect 1610 1174 1623 1196
rect 1638 1174 1668 1196
rect 1695 1174 1696 1190
rect 1711 1174 1724 1334
rect 1754 1230 1767 1334
rect 1812 1312 1813 1322
rect 1828 1312 1837 1322
rect 1812 1306 1837 1312
rect 1796 1298 1837 1306
rect 1796 1286 1821 1298
rect 1828 1286 1837 1298
rect 1796 1278 1837 1286
rect 1812 1270 1813 1278
rect 1828 1270 1837 1278
rect 1812 1262 1828 1270
rect 1809 1255 1828 1258
rect 1809 1246 1831 1255
rect 1782 1236 1831 1246
rect 1782 1230 1812 1236
rect 1831 1231 1836 1236
rect 3494 1230 3507 1334
rect 3552 1312 3553 1322
rect 3568 1312 3581 1322
rect 3552 1308 3581 1312
rect 3586 1308 3616 1334
rect 3634 1320 3650 1322
rect 3722 1320 3775 1334
rect 3723 1318 3787 1320
rect 3830 1318 3845 1334
rect 3894 1331 3924 1334
rect 3894 1328 3930 1331
rect 3860 1320 3876 1322
rect 3634 1308 3649 1312
rect 3552 1306 3649 1308
rect 3677 1306 3845 1318
rect 3861 1308 3876 1312
rect 3894 1309 3933 1328
rect 3952 1322 3959 1323
rect 3958 1315 3959 1322
rect 3942 1312 3943 1315
rect 3958 1312 3971 1315
rect 3894 1308 3924 1309
rect 3933 1308 3939 1309
rect 3942 1308 3971 1312
rect 3861 1307 3971 1308
rect 3861 1306 3977 1307
rect 3536 1298 3587 1306
rect 3536 1286 3561 1298
rect 3568 1286 3587 1298
rect 3618 1298 3668 1306
rect 3618 1290 3634 1298
rect 3641 1296 3668 1298
rect 3677 1296 3898 1306
rect 3641 1286 3898 1296
rect 3927 1298 3977 1306
rect 3927 1289 3943 1298
rect 3536 1278 3587 1286
rect 3634 1278 3898 1286
rect 3924 1286 3943 1289
rect 3950 1286 3977 1298
rect 3924 1278 3977 1286
rect 3552 1270 3553 1278
rect 3568 1270 3581 1278
rect 3552 1262 3568 1270
rect 3549 1255 3568 1258
rect 3549 1246 3571 1255
rect 3522 1236 3571 1246
rect 3522 1230 3552 1236
rect 3571 1231 3576 1236
rect 1754 1214 1828 1230
rect 3494 1214 3568 1230
rect 3586 1222 3616 1278
rect 3651 1268 3859 1278
rect 3894 1274 3939 1278
rect 3942 1277 3943 1278
rect 3958 1277 3971 1278
rect 3677 1238 3866 1268
rect 3692 1235 3866 1238
rect 3685 1232 3866 1235
rect 1754 1212 1767 1214
rect 1782 1212 1816 1214
rect 3494 1212 3507 1214
rect 3522 1212 3556 1214
rect 1754 1196 1828 1212
rect 3494 1196 3568 1212
rect 3595 1208 3608 1222
rect 3623 1208 3639 1224
rect 3685 1219 3696 1232
rect 1738 1174 1739 1190
rect 1754 1174 1767 1196
rect 1782 1174 1812 1196
rect 3494 1174 3507 1196
rect 3522 1174 3552 1196
rect 3595 1192 3657 1208
rect 3685 1201 3696 1217
rect 3701 1212 3711 1232
rect 3721 1212 3735 1232
rect 3738 1219 3747 1232
rect 3763 1219 3772 1232
rect 3701 1201 3735 1212
rect 3738 1201 3747 1217
rect 3763 1201 3772 1217
rect 3779 1212 3789 1232
rect 3799 1212 3813 1232
rect 3814 1219 3825 1232
rect 3779 1201 3813 1212
rect 3814 1201 3825 1217
rect 3871 1208 3887 1224
rect 3894 1222 3924 1274
rect 3958 1270 3959 1277
rect 3943 1262 3959 1270
rect 3930 1230 3943 1249
rect 3958 1230 3988 1246
rect 3930 1214 4004 1230
rect 3930 1212 3943 1214
rect 3958 1212 3992 1214
rect 3595 1190 3608 1192
rect 3623 1190 3657 1192
rect 3595 1174 3657 1190
rect 3701 1185 3717 1192
rect 3779 1185 3809 1196
rect 3857 1192 3903 1208
rect 3930 1196 4004 1212
rect 3857 1190 3891 1192
rect 3856 1174 3903 1190
rect 3930 1174 3943 1196
rect 3958 1174 3988 1196
rect 4015 1174 4016 1190
rect 4031 1174 4044 1334
rect 4074 1230 4087 1334
rect 4132 1312 4133 1322
rect 4148 1312 4161 1322
rect 4132 1308 4161 1312
rect 4166 1308 4196 1334
rect 4214 1320 4230 1322
rect 4302 1320 4355 1334
rect 4303 1318 4367 1320
rect 4410 1318 4425 1334
rect 4474 1331 4504 1334
rect 4474 1328 4510 1331
rect 4440 1320 4456 1322
rect 4214 1308 4229 1312
rect 4132 1306 4229 1308
rect 4257 1306 4425 1318
rect 4441 1308 4456 1312
rect 4474 1309 4513 1328
rect 4532 1322 4539 1323
rect 4538 1315 4539 1322
rect 4522 1312 4523 1315
rect 4538 1312 4551 1315
rect 4474 1308 4504 1309
rect 4513 1308 4519 1309
rect 4522 1308 4551 1312
rect 4441 1307 4551 1308
rect 4441 1306 4557 1307
rect 4116 1298 4167 1306
rect 4116 1286 4141 1298
rect 4148 1286 4167 1298
rect 4198 1298 4248 1306
rect 4198 1290 4214 1298
rect 4221 1296 4248 1298
rect 4257 1296 4478 1306
rect 4221 1286 4478 1296
rect 4507 1298 4557 1306
rect 4507 1289 4523 1298
rect 4116 1278 4167 1286
rect 4214 1278 4478 1286
rect 4504 1286 4523 1289
rect 4530 1286 4557 1298
rect 4504 1278 4557 1286
rect 4132 1270 4133 1278
rect 4148 1270 4161 1278
rect 4132 1262 4148 1270
rect 4129 1255 4148 1258
rect 4129 1246 4151 1255
rect 4102 1236 4151 1246
rect 4102 1230 4132 1236
rect 4151 1231 4156 1236
rect 4074 1214 4148 1230
rect 4166 1222 4196 1278
rect 4231 1268 4439 1278
rect 4474 1274 4519 1278
rect 4522 1277 4523 1278
rect 4538 1277 4551 1278
rect 4257 1238 4446 1268
rect 4272 1235 4446 1238
rect 4265 1232 4446 1235
rect 4074 1212 4087 1214
rect 4102 1212 4136 1214
rect 4074 1196 4148 1212
rect 4175 1208 4188 1222
rect 4203 1208 4219 1224
rect 4265 1219 4276 1232
rect 4058 1174 4059 1190
rect 4074 1174 4087 1196
rect 4102 1174 4132 1196
rect 4175 1192 4237 1208
rect 4265 1201 4276 1217
rect 4281 1212 4291 1232
rect 4301 1212 4315 1232
rect 4318 1219 4327 1232
rect 4343 1219 4352 1232
rect 4281 1201 4315 1212
rect 4318 1201 4327 1217
rect 4343 1201 4352 1217
rect 4359 1212 4369 1232
rect 4379 1212 4393 1232
rect 4394 1219 4405 1232
rect 4359 1201 4393 1212
rect 4394 1201 4405 1217
rect 4451 1208 4467 1224
rect 4474 1222 4504 1274
rect 4538 1270 4539 1277
rect 4523 1262 4539 1270
rect 4510 1230 4523 1249
rect 4538 1230 4568 1246
rect 4510 1214 4584 1230
rect 4510 1212 4523 1214
rect 4538 1212 4572 1214
rect 4175 1190 4188 1192
rect 4203 1190 4237 1192
rect 4175 1174 4237 1190
rect 4281 1185 4297 1192
rect 4359 1185 4389 1196
rect 4437 1192 4483 1208
rect 4510 1196 4584 1212
rect 4437 1190 4471 1192
rect 4436 1174 4483 1190
rect 4510 1174 4523 1196
rect 4538 1174 4568 1196
rect 4595 1174 4596 1190
rect 4611 1174 4624 1334
rect 4654 1230 4667 1334
rect 4712 1312 4713 1322
rect 4728 1312 4741 1322
rect 4712 1308 4741 1312
rect 4746 1308 4776 1334
rect 4794 1320 4810 1322
rect 4882 1320 4935 1334
rect 4883 1318 4947 1320
rect 4899 1317 4931 1318
rect 4990 1317 5005 1334
rect 5054 1331 5084 1334
rect 5054 1328 5090 1331
rect 5020 1320 5036 1322
rect 4794 1308 4809 1312
rect 4712 1306 4809 1308
rect 4837 1306 5005 1317
rect 5021 1308 5036 1312
rect 5054 1309 5093 1328
rect 5112 1322 5119 1323
rect 5118 1315 5119 1322
rect 5102 1312 5103 1315
rect 5118 1312 5131 1315
rect 5054 1308 5084 1309
rect 5093 1308 5099 1309
rect 5102 1308 5131 1312
rect 5021 1307 5131 1308
rect 5021 1306 5137 1307
rect 4696 1298 4747 1306
rect 4696 1286 4721 1298
rect 4728 1286 4747 1298
rect 4778 1298 4828 1306
rect 4778 1290 4794 1298
rect 4801 1296 4828 1298
rect 4837 1296 5058 1306
rect 4801 1286 5058 1296
rect 5087 1298 5137 1306
rect 5087 1289 5103 1298
rect 4696 1278 4747 1286
rect 4794 1278 5058 1286
rect 5084 1286 5103 1289
rect 5110 1286 5137 1298
rect 5084 1278 5137 1286
rect 4712 1270 4713 1278
rect 4728 1270 4741 1278
rect 4712 1262 4728 1270
rect 4709 1255 4728 1258
rect 4709 1246 4731 1255
rect 4682 1236 4731 1246
rect 4682 1230 4712 1236
rect 4731 1231 4736 1236
rect 4654 1214 4728 1230
rect 4746 1222 4776 1278
rect 4811 1268 5019 1278
rect 5054 1274 5099 1278
rect 5102 1277 5103 1278
rect 5118 1277 5131 1278
rect 4837 1238 5026 1268
rect 4852 1235 5026 1238
rect 4845 1232 5026 1235
rect 4654 1212 4667 1214
rect 4682 1212 4716 1214
rect 4654 1196 4728 1212
rect 4755 1208 4768 1222
rect 4783 1208 4799 1224
rect 4845 1219 4856 1232
rect 4638 1174 4639 1190
rect 4654 1174 4667 1196
rect 4682 1174 4712 1196
rect 4755 1192 4817 1208
rect 4845 1201 4856 1217
rect 4861 1212 4871 1232
rect 4881 1212 4895 1232
rect 4898 1219 4907 1232
rect 4923 1219 4932 1232
rect 4861 1201 4895 1212
rect 4898 1201 4907 1217
rect 4923 1201 4932 1217
rect 4939 1212 4949 1232
rect 4959 1212 4973 1232
rect 4974 1219 4985 1232
rect 4939 1201 4973 1212
rect 4974 1201 4985 1217
rect 5031 1208 5047 1224
rect 5054 1222 5084 1274
rect 5118 1270 5119 1277
rect 5103 1262 5119 1270
rect 5090 1230 5103 1249
rect 5118 1230 5148 1246
rect 5090 1214 5164 1230
rect 5090 1212 5103 1214
rect 5118 1212 5152 1214
rect 4755 1190 4768 1192
rect 4783 1190 4817 1192
rect 4755 1174 4817 1190
rect 4861 1185 4877 1192
rect 4939 1185 4969 1196
rect 5017 1192 5063 1208
rect 5090 1196 5164 1212
rect 5017 1190 5051 1192
rect 5016 1174 5063 1190
rect 5090 1174 5103 1196
rect 5118 1174 5148 1196
rect 5175 1174 5176 1190
rect 5191 1174 5204 1334
rect 5234 1230 5247 1334
rect 5292 1312 5293 1322
rect 5308 1312 5321 1322
rect 5292 1308 5321 1312
rect 5326 1308 5356 1334
rect 5374 1320 5390 1322
rect 5462 1320 5515 1334
rect 5463 1318 5527 1320
rect 5479 1317 5511 1318
rect 5570 1317 5585 1334
rect 5634 1331 5664 1334
rect 5634 1328 5670 1331
rect 5600 1320 5616 1322
rect 5374 1308 5389 1312
rect 5292 1306 5389 1308
rect 5417 1306 5585 1317
rect 5601 1308 5616 1312
rect 5634 1309 5673 1328
rect 5692 1322 5699 1323
rect 5698 1315 5699 1322
rect 5682 1312 5683 1315
rect 5698 1312 5711 1315
rect 5634 1308 5664 1309
rect 5673 1308 5679 1309
rect 5682 1308 5711 1312
rect 5601 1307 5711 1308
rect 5601 1306 5717 1307
rect 5276 1298 5327 1306
rect 5276 1286 5301 1298
rect 5308 1286 5327 1298
rect 5358 1298 5408 1306
rect 5358 1290 5374 1298
rect 5381 1296 5408 1298
rect 5417 1296 5638 1306
rect 5381 1286 5638 1296
rect 5667 1298 5717 1306
rect 5667 1289 5683 1298
rect 5276 1278 5327 1286
rect 5374 1278 5638 1286
rect 5664 1286 5683 1289
rect 5690 1286 5717 1298
rect 5664 1278 5717 1286
rect 5292 1270 5293 1278
rect 5308 1270 5321 1278
rect 5292 1262 5308 1270
rect 5289 1255 5308 1258
rect 5289 1246 5311 1255
rect 5262 1236 5311 1246
rect 5262 1230 5292 1236
rect 5311 1231 5316 1236
rect 5234 1214 5308 1230
rect 5326 1222 5356 1278
rect 5391 1268 5599 1278
rect 5634 1274 5679 1278
rect 5682 1277 5683 1278
rect 5698 1277 5711 1278
rect 5417 1238 5606 1268
rect 5432 1235 5606 1238
rect 5425 1232 5606 1235
rect 5234 1212 5247 1214
rect 5262 1212 5296 1214
rect 5234 1196 5308 1212
rect 5335 1208 5348 1222
rect 5363 1208 5379 1224
rect 5425 1219 5436 1232
rect 5218 1174 5219 1190
rect 5234 1174 5247 1196
rect 5262 1174 5292 1196
rect 5335 1192 5397 1208
rect 5425 1201 5436 1217
rect 5441 1212 5451 1232
rect 5461 1212 5475 1232
rect 5478 1219 5487 1232
rect 5503 1219 5512 1232
rect 5441 1201 5475 1212
rect 5478 1201 5487 1217
rect 5503 1201 5512 1217
rect 5519 1212 5529 1232
rect 5539 1212 5553 1232
rect 5554 1219 5565 1232
rect 5519 1201 5553 1212
rect 5554 1201 5565 1217
rect 5611 1208 5627 1224
rect 5634 1222 5664 1274
rect 5698 1270 5699 1277
rect 5683 1262 5699 1270
rect 5670 1230 5683 1249
rect 5698 1230 5728 1246
rect 5670 1214 5744 1230
rect 5670 1212 5683 1214
rect 5698 1212 5732 1214
rect 5335 1190 5348 1192
rect 5363 1190 5397 1192
rect 5335 1174 5397 1190
rect 5441 1185 5457 1192
rect 5519 1185 5549 1196
rect 5597 1192 5643 1208
rect 5670 1196 5744 1212
rect 5597 1190 5631 1192
rect 5596 1174 5643 1190
rect 5670 1174 5683 1196
rect 5698 1174 5728 1196
rect 5755 1174 5756 1190
rect 5771 1174 5784 1334
rect 5814 1230 5827 1334
rect 5872 1312 5873 1322
rect 5888 1312 5901 1322
rect 5872 1308 5901 1312
rect 5906 1308 5936 1334
rect 5954 1320 5970 1322
rect 6042 1320 6095 1334
rect 6043 1318 6107 1320
rect 6059 1317 6091 1318
rect 6150 1317 6165 1334
rect 6214 1331 6244 1334
rect 6214 1328 6250 1331
rect 6180 1320 6196 1322
rect 5954 1308 5969 1312
rect 5872 1306 5969 1308
rect 5997 1306 6165 1317
rect 6181 1308 6196 1312
rect 6214 1309 6253 1328
rect 6272 1322 6279 1323
rect 6278 1315 6279 1322
rect 6262 1312 6263 1315
rect 6278 1312 6291 1315
rect 6214 1308 6244 1309
rect 6253 1308 6259 1309
rect 6262 1308 6291 1312
rect 6181 1307 6291 1308
rect 6181 1306 6297 1307
rect 5856 1298 5907 1306
rect 5856 1286 5881 1298
rect 5888 1286 5907 1298
rect 5938 1298 5988 1306
rect 5938 1290 5954 1298
rect 5961 1296 5988 1298
rect 5997 1296 6218 1306
rect 5961 1286 6218 1296
rect 6247 1298 6297 1306
rect 6247 1289 6263 1298
rect 5856 1278 5907 1286
rect 5954 1278 6218 1286
rect 6244 1286 6263 1289
rect 6270 1286 6297 1298
rect 6244 1278 6297 1286
rect 5872 1270 5873 1278
rect 5888 1270 5901 1278
rect 5872 1262 5888 1270
rect 5869 1255 5888 1258
rect 5869 1246 5891 1255
rect 5842 1236 5891 1246
rect 5842 1230 5872 1236
rect 5891 1231 5896 1236
rect 5814 1214 5888 1230
rect 5906 1222 5936 1278
rect 5971 1268 6179 1278
rect 6214 1274 6259 1278
rect 6262 1277 6263 1278
rect 6278 1277 6291 1278
rect 5997 1238 6186 1268
rect 6012 1235 6186 1238
rect 6005 1232 6186 1235
rect 5814 1212 5827 1214
rect 5842 1212 5876 1214
rect 5814 1196 5888 1212
rect 5915 1208 5928 1222
rect 5943 1208 5959 1224
rect 6005 1219 6016 1232
rect 5798 1174 5799 1190
rect 5814 1174 5827 1196
rect 5842 1174 5872 1196
rect 5915 1192 5977 1208
rect 6005 1201 6016 1217
rect 6021 1212 6031 1232
rect 6041 1212 6055 1232
rect 6058 1219 6067 1232
rect 6083 1219 6092 1232
rect 6021 1201 6055 1212
rect 6058 1201 6067 1217
rect 6083 1201 6092 1217
rect 6099 1212 6109 1232
rect 6119 1212 6133 1232
rect 6134 1219 6145 1232
rect 6099 1201 6133 1212
rect 6134 1201 6145 1217
rect 6191 1208 6207 1224
rect 6214 1222 6244 1274
rect 6278 1270 6279 1277
rect 6263 1262 6279 1270
rect 6250 1230 6263 1249
rect 6278 1230 6308 1246
rect 6250 1214 6324 1230
rect 6250 1212 6263 1214
rect 6278 1212 6312 1214
rect 5915 1190 5928 1192
rect 5943 1190 5977 1192
rect 5915 1174 5977 1190
rect 6021 1185 6037 1192
rect 6099 1185 6129 1196
rect 6177 1192 6223 1208
rect 6250 1196 6324 1212
rect 6177 1190 6211 1192
rect 6176 1174 6223 1190
rect 6250 1174 6263 1196
rect 6278 1174 6308 1196
rect 6335 1174 6336 1190
rect 6351 1174 6364 1334
rect 6394 1230 6407 1334
rect 6452 1312 6453 1322
rect 6468 1312 6481 1322
rect 6452 1308 6481 1312
rect 6486 1308 6516 1334
rect 6534 1320 6550 1322
rect 6622 1320 6675 1334
rect 6623 1318 6687 1320
rect 6639 1317 6671 1318
rect 6730 1317 6745 1334
rect 6794 1331 6824 1334
rect 6794 1328 6830 1331
rect 6760 1320 6776 1322
rect 6534 1308 6549 1312
rect 6452 1306 6549 1308
rect 6577 1306 6745 1317
rect 6761 1308 6776 1312
rect 6794 1309 6833 1328
rect 6852 1322 6859 1323
rect 6858 1315 6859 1322
rect 6842 1312 6843 1315
rect 6858 1312 6871 1315
rect 6794 1308 6824 1309
rect 6833 1308 6839 1309
rect 6842 1308 6871 1312
rect 6761 1307 6871 1308
rect 6761 1306 6877 1307
rect 6436 1298 6487 1306
rect 6436 1286 6461 1298
rect 6468 1286 6487 1298
rect 6518 1298 6568 1306
rect 6518 1290 6534 1298
rect 6541 1296 6568 1298
rect 6577 1296 6798 1306
rect 6541 1286 6798 1296
rect 6827 1298 6877 1306
rect 6827 1289 6843 1298
rect 6436 1278 6487 1286
rect 6534 1278 6798 1286
rect 6824 1286 6843 1289
rect 6850 1286 6877 1298
rect 6824 1278 6877 1286
rect 6452 1270 6453 1278
rect 6468 1270 6481 1278
rect 6452 1262 6468 1270
rect 6449 1255 6468 1258
rect 6449 1246 6471 1255
rect 6422 1236 6471 1246
rect 6422 1230 6452 1236
rect 6471 1231 6476 1236
rect 6394 1214 6468 1230
rect 6486 1222 6516 1278
rect 6551 1268 6759 1278
rect 6794 1274 6839 1278
rect 6842 1277 6843 1278
rect 6858 1277 6871 1278
rect 6577 1238 6766 1268
rect 6592 1235 6766 1238
rect 6585 1232 6766 1235
rect 6394 1212 6407 1214
rect 6422 1212 6456 1214
rect 6394 1196 6468 1212
rect 6495 1208 6508 1222
rect 6523 1208 6539 1224
rect 6585 1219 6596 1232
rect 6378 1174 6379 1190
rect 6394 1174 6407 1196
rect 6422 1174 6452 1196
rect 6495 1192 6557 1208
rect 6585 1201 6596 1217
rect 6601 1212 6611 1232
rect 6621 1212 6635 1232
rect 6638 1219 6647 1232
rect 6663 1219 6672 1232
rect 6601 1201 6635 1212
rect 6638 1201 6647 1217
rect 6663 1201 6672 1217
rect 6679 1212 6689 1232
rect 6699 1212 6713 1232
rect 6714 1219 6725 1232
rect 6679 1201 6713 1212
rect 6714 1201 6725 1217
rect 6771 1208 6787 1224
rect 6794 1222 6824 1274
rect 6858 1270 6859 1277
rect 6843 1262 6859 1270
rect 6830 1230 6843 1249
rect 6858 1230 6888 1246
rect 6830 1214 6904 1230
rect 6830 1212 6843 1214
rect 6858 1212 6892 1214
rect 6495 1190 6508 1192
rect 6523 1190 6557 1192
rect 6495 1174 6557 1190
rect 6601 1185 6617 1192
rect 6679 1185 6709 1196
rect 6757 1192 6803 1208
rect 6830 1196 6904 1212
rect 6757 1190 6791 1192
rect 6756 1174 6803 1190
rect 6830 1174 6843 1196
rect 6858 1174 6888 1196
rect 6915 1174 6916 1190
rect 6931 1174 6944 1334
rect -8 1166 33 1174
rect -8 1140 7 1166
rect 14 1140 33 1166
rect 97 1162 159 1174
rect 171 1162 246 1174
rect 304 1162 379 1174
rect 391 1162 422 1174
rect 428 1162 463 1174
rect 97 1160 259 1162
rect -8 1132 33 1140
rect 115 1136 128 1160
rect 143 1158 158 1160
rect -2 1122 -1 1132
rect 14 1122 27 1132
rect 42 1122 72 1136
rect 115 1122 158 1136
rect 182 1133 189 1140
rect 192 1136 259 1160
rect 291 1160 463 1162
rect 261 1138 289 1142
rect 291 1138 371 1160
rect 392 1158 407 1160
rect 261 1136 371 1138
rect 192 1132 371 1136
rect 165 1122 195 1132
rect 197 1122 350 1132
rect 358 1122 388 1132
rect 392 1122 422 1136
rect 450 1122 463 1160
rect 535 1166 570 1174
rect 535 1140 536 1166
rect 543 1140 570 1166
rect 478 1122 508 1136
rect 535 1132 570 1140
rect 572 1166 613 1174
rect 572 1140 587 1166
rect 594 1140 613 1166
rect 677 1162 739 1174
rect 751 1162 826 1174
rect 884 1162 959 1174
rect 971 1162 1002 1174
rect 1008 1162 1043 1174
rect 677 1160 839 1162
rect 572 1132 613 1140
rect 695 1136 708 1160
rect 723 1158 738 1160
rect 535 1122 536 1132
rect 551 1122 564 1132
rect 578 1122 579 1132
rect 594 1122 607 1132
rect 622 1122 652 1136
rect 695 1122 738 1136
rect 762 1133 769 1140
rect 772 1136 839 1160
rect 871 1160 1043 1162
rect 841 1138 869 1142
rect 871 1138 951 1160
rect 972 1158 987 1160
rect 841 1136 951 1138
rect 772 1132 951 1136
rect 745 1122 775 1132
rect 777 1122 930 1132
rect 938 1122 968 1132
rect 972 1122 1002 1136
rect 1030 1122 1043 1160
rect 1115 1166 1150 1174
rect 1115 1140 1116 1166
rect 1123 1140 1150 1166
rect 1058 1122 1088 1136
rect 1115 1132 1150 1140
rect 1152 1166 1193 1174
rect 1152 1140 1167 1166
rect 1174 1140 1193 1166
rect 1257 1162 1319 1174
rect 1331 1162 1406 1174
rect 1464 1162 1539 1174
rect 1551 1162 1582 1174
rect 1588 1162 1623 1174
rect 1257 1160 1419 1162
rect 1152 1132 1193 1140
rect 1275 1136 1288 1160
rect 1303 1158 1318 1160
rect 1115 1122 1116 1132
rect 1131 1122 1144 1132
rect 1158 1122 1159 1132
rect 1174 1122 1187 1132
rect 1202 1122 1232 1136
rect 1275 1122 1318 1136
rect 1342 1133 1349 1140
rect 1352 1136 1419 1160
rect 1451 1160 1623 1162
rect 1421 1138 1449 1142
rect 1451 1138 1531 1160
rect 1552 1158 1567 1160
rect 1421 1136 1531 1138
rect 1352 1132 1531 1136
rect 1325 1122 1355 1132
rect 1357 1122 1510 1132
rect 1518 1122 1548 1132
rect 1552 1122 1582 1136
rect 1610 1122 1623 1160
rect 1695 1166 1730 1174
rect 1695 1140 1696 1166
rect 1703 1140 1730 1166
rect 1638 1122 1668 1136
rect 1695 1132 1730 1140
rect 1732 1166 1773 1174
rect 1732 1140 1747 1166
rect 1754 1140 1773 1166
rect 1732 1132 1773 1140
rect 3481 1166 3513 1174
rect 3481 1140 3487 1166
rect 3494 1140 3513 1166
rect 3577 1162 3639 1174
rect 3651 1162 3726 1174
rect 3784 1162 3859 1174
rect 3871 1162 3902 1174
rect 3908 1162 3943 1174
rect 3577 1160 3739 1162
rect 1695 1122 1696 1132
rect 1711 1122 1724 1132
rect 1738 1122 1739 1132
rect 1754 1122 1767 1132
rect 1782 1122 1812 1136
rect 3481 1132 3513 1140
rect 3595 1136 3608 1160
rect 3623 1158 3638 1160
rect 3494 1122 3507 1132
rect 3522 1122 3552 1136
rect 3595 1122 3638 1136
rect 3662 1133 3669 1140
rect 3672 1136 3739 1160
rect 3771 1160 3943 1162
rect 3741 1138 3769 1142
rect 3771 1138 3851 1160
rect 3872 1158 3887 1160
rect 3741 1136 3851 1138
rect 3672 1132 3851 1136
rect 3645 1122 3675 1132
rect 3677 1122 3830 1132
rect 3838 1122 3868 1132
rect 3872 1122 3902 1136
rect 3930 1122 3943 1160
rect 4015 1166 4050 1174
rect 4015 1140 4016 1166
rect 4023 1140 4050 1166
rect 3958 1122 3988 1136
rect 4015 1132 4050 1140
rect 4052 1166 4093 1174
rect 4052 1140 4067 1166
rect 4074 1140 4093 1166
rect 4157 1162 4219 1174
rect 4231 1162 4306 1174
rect 4364 1162 4439 1174
rect 4451 1162 4482 1174
rect 4488 1162 4523 1174
rect 4157 1160 4319 1162
rect 4052 1132 4093 1140
rect 4175 1136 4188 1160
rect 4203 1158 4218 1160
rect 4015 1122 4016 1132
rect 4031 1122 4044 1132
rect 4058 1122 4059 1132
rect 4074 1122 4087 1132
rect 4102 1122 4132 1136
rect 4175 1122 4218 1136
rect 4242 1133 4249 1140
rect 4252 1136 4319 1160
rect 4351 1160 4523 1162
rect 4321 1138 4349 1142
rect 4351 1138 4431 1160
rect 4452 1158 4467 1160
rect 4321 1136 4431 1138
rect 4252 1132 4431 1136
rect 4225 1122 4255 1132
rect 4257 1122 4410 1132
rect 4418 1122 4448 1132
rect 4452 1122 4482 1136
rect 4510 1122 4523 1160
rect 4595 1166 4630 1174
rect 4595 1140 4596 1166
rect 4603 1140 4630 1166
rect 4538 1122 4568 1136
rect 4595 1132 4630 1140
rect 4632 1166 4673 1174
rect 4632 1140 4647 1166
rect 4654 1140 4673 1166
rect 4737 1162 4799 1174
rect 4811 1162 4886 1174
rect 4944 1162 5019 1174
rect 5031 1162 5062 1174
rect 5068 1162 5103 1174
rect 4737 1160 4899 1162
rect 4755 1141 4768 1160
rect 4783 1158 4798 1160
rect 4632 1132 4673 1140
rect 4756 1135 4768 1141
rect 4595 1122 4596 1132
rect 4611 1122 4624 1132
rect 4638 1122 4639 1132
rect 4654 1122 4667 1132
rect 4682 1122 4712 1135
rect 4756 1122 4798 1135
rect 4822 1133 4829 1140
rect 4832 1135 4899 1160
rect 4931 1160 5103 1162
rect 4901 1138 4929 1142
rect 4931 1138 5011 1160
rect 5032 1158 5047 1160
rect 4901 1136 5011 1138
rect 4901 1135 4929 1136
rect 4931 1135 5011 1136
rect 4832 1132 5011 1135
rect 4805 1131 4813 1132
rect 4832 1131 4835 1132
rect 4805 1124 4835 1131
rect 4837 1124 4990 1132
rect 5017 1131 5028 1132
rect 4998 1124 5028 1131
rect 4805 1122 5028 1124
rect 5032 1122 5062 1135
rect 5090 1122 5103 1160
rect 5175 1166 5210 1174
rect 5175 1140 5176 1166
rect 5183 1140 5210 1166
rect 5118 1122 5148 1135
rect 5175 1132 5210 1140
rect 5212 1166 5253 1174
rect 5212 1140 5227 1166
rect 5234 1140 5253 1166
rect 5317 1162 5379 1174
rect 5391 1162 5466 1174
rect 5524 1162 5599 1174
rect 5611 1162 5642 1174
rect 5648 1162 5683 1174
rect 5317 1160 5479 1162
rect 5335 1141 5348 1160
rect 5363 1158 5378 1160
rect 5212 1132 5253 1140
rect 5336 1135 5348 1141
rect 5175 1122 5176 1132
rect 5191 1122 5204 1132
rect 5218 1122 5219 1132
rect 5234 1122 5247 1132
rect 5262 1122 5292 1135
rect 5336 1122 5378 1135
rect 5402 1133 5409 1140
rect 5412 1135 5479 1160
rect 5511 1160 5683 1162
rect 5481 1138 5509 1142
rect 5511 1138 5591 1160
rect 5612 1158 5627 1160
rect 5481 1136 5591 1138
rect 5481 1135 5509 1136
rect 5511 1135 5591 1136
rect 5412 1132 5591 1135
rect 5385 1131 5393 1132
rect 5412 1131 5415 1132
rect 5385 1124 5415 1131
rect 5417 1124 5570 1132
rect 5597 1131 5608 1132
rect 5578 1124 5608 1131
rect 5385 1122 5608 1124
rect 5612 1122 5642 1135
rect 5670 1122 5683 1160
rect 5755 1166 5790 1174
rect 5755 1140 5756 1166
rect 5763 1140 5790 1166
rect 5698 1122 5728 1135
rect 5755 1132 5790 1140
rect 5792 1166 5833 1174
rect 5792 1140 5807 1166
rect 5814 1140 5833 1166
rect 5897 1162 5959 1174
rect 5971 1162 6046 1174
rect 6104 1162 6179 1174
rect 6191 1162 6222 1174
rect 6228 1162 6263 1174
rect 5897 1160 6059 1162
rect 5915 1141 5928 1160
rect 5943 1158 5958 1160
rect 5792 1132 5833 1140
rect 5916 1135 5928 1141
rect 5755 1122 5756 1132
rect 5771 1122 5784 1132
rect 5798 1122 5799 1132
rect 5814 1122 5827 1132
rect 5842 1122 5872 1135
rect 5916 1122 5958 1135
rect 5982 1133 5989 1140
rect 5992 1135 6059 1160
rect 6091 1160 6263 1162
rect 6061 1138 6089 1142
rect 6091 1138 6171 1160
rect 6192 1158 6207 1160
rect 6061 1136 6171 1138
rect 6061 1135 6089 1136
rect 6091 1135 6171 1136
rect 5992 1132 6171 1135
rect 5965 1131 5973 1132
rect 5992 1131 5995 1132
rect 5965 1124 5995 1131
rect 5997 1124 6150 1132
rect 6177 1131 6188 1132
rect 6158 1124 6188 1131
rect 5965 1122 6188 1124
rect 6192 1122 6222 1135
rect 6250 1122 6263 1160
rect 6335 1166 6370 1174
rect 6335 1140 6336 1166
rect 6343 1140 6370 1166
rect 6278 1122 6308 1135
rect 6335 1132 6370 1140
rect 6372 1166 6413 1174
rect 6372 1140 6387 1166
rect 6394 1140 6413 1166
rect 6477 1162 6539 1174
rect 6551 1162 6626 1174
rect 6684 1162 6759 1174
rect 6771 1162 6802 1174
rect 6808 1162 6843 1174
rect 6477 1160 6639 1162
rect 6495 1141 6508 1160
rect 6523 1158 6538 1160
rect 6372 1132 6413 1140
rect 6496 1135 6508 1141
rect 6335 1122 6336 1132
rect 6351 1122 6364 1132
rect 6378 1122 6379 1132
rect 6394 1122 6407 1132
rect 6422 1122 6452 1135
rect 6496 1122 6538 1135
rect 6562 1133 6569 1140
rect 6572 1135 6639 1160
rect 6671 1160 6843 1162
rect 6641 1138 6669 1142
rect 6671 1138 6751 1160
rect 6772 1158 6787 1160
rect 6641 1136 6751 1138
rect 6641 1135 6669 1136
rect 6671 1135 6751 1136
rect 6572 1132 6751 1135
rect 6545 1131 6553 1132
rect 6572 1131 6575 1132
rect 6545 1124 6575 1131
rect 6577 1124 6730 1132
rect 6757 1131 6768 1132
rect 6738 1124 6768 1131
rect 6545 1122 6768 1124
rect 6772 1122 6802 1135
rect 6830 1122 6843 1160
rect 6915 1166 6950 1174
rect 6915 1140 6916 1166
rect 6923 1140 6950 1166
rect 6858 1122 6888 1135
rect 6915 1132 6950 1140
rect 6915 1122 6916 1132
rect 6931 1122 6944 1132
rect -2 1116 1837 1122
rect -1 1108 1837 1116
rect 3481 1108 6944 1122
rect 14 1078 27 1108
rect 42 1090 72 1108
rect 115 1094 129 1108
rect 165 1094 385 1108
rect 116 1092 129 1094
rect 82 1080 97 1092
rect 79 1078 101 1080
rect 106 1078 136 1092
rect 197 1090 350 1094
rect 179 1078 371 1090
rect 414 1078 444 1092
rect 450 1078 463 1108
rect 478 1090 508 1108
rect 551 1078 564 1108
rect 594 1078 607 1108
rect 622 1090 652 1108
rect 695 1094 709 1108
rect 745 1094 965 1108
rect 696 1092 709 1094
rect 662 1080 677 1092
rect 659 1078 681 1080
rect 686 1078 716 1092
rect 777 1090 930 1094
rect 759 1078 951 1090
rect 994 1078 1024 1092
rect 1030 1078 1043 1108
rect 1058 1090 1088 1108
rect 1131 1078 1144 1108
rect 1174 1078 1187 1108
rect 1202 1090 1232 1108
rect 1275 1094 1289 1108
rect 1325 1094 1545 1108
rect 1276 1092 1289 1094
rect 1242 1080 1257 1092
rect 1239 1078 1261 1080
rect 1266 1078 1296 1092
rect 1357 1090 1510 1094
rect 1339 1078 1531 1090
rect 1574 1078 1604 1092
rect 1610 1078 1623 1108
rect 1638 1090 1668 1108
rect 1711 1078 1724 1108
rect 1754 1078 1767 1108
rect 1782 1090 1812 1108
rect 1822 1080 1837 1092
rect 1819 1078 1837 1080
rect 3494 1078 3507 1108
rect 3522 1090 3552 1108
rect 3595 1094 3609 1108
rect 3645 1094 3865 1108
rect 3596 1092 3609 1094
rect 3562 1080 3577 1092
rect 3559 1078 3581 1080
rect 3586 1078 3616 1092
rect 3677 1090 3830 1094
rect 3659 1078 3851 1090
rect 3894 1078 3924 1092
rect 3930 1078 3943 1108
rect 3958 1090 3988 1108
rect 4031 1078 4044 1108
rect 4074 1078 4087 1108
rect 4102 1090 4132 1108
rect 4175 1094 4189 1108
rect 4225 1094 4445 1108
rect 4176 1092 4189 1094
rect 4142 1080 4157 1092
rect 4139 1078 4161 1080
rect 4166 1078 4196 1092
rect 4257 1090 4410 1094
rect 4239 1078 4431 1090
rect 4474 1078 4504 1092
rect 4510 1078 4523 1108
rect 4538 1090 4568 1108
rect 4611 1078 4624 1108
rect -1 1064 1837 1078
rect 3481 1077 4624 1078
rect 4654 1077 4667 1108
rect 4682 1090 4712 1108
rect 4756 1091 4769 1108
rect 4805 1094 5025 1108
rect 4722 1079 4737 1091
rect 4719 1077 4741 1079
rect 4746 1077 4776 1091
rect 4837 1089 4990 1094
rect 4819 1077 5011 1089
rect 5054 1077 5084 1091
rect 5090 1077 5103 1108
rect 5118 1090 5148 1108
rect 5191 1077 5204 1108
rect 5234 1077 5247 1108
rect 5262 1090 5292 1108
rect 5336 1091 5349 1108
rect 5385 1094 5605 1108
rect 5302 1079 5317 1091
rect 5299 1077 5321 1079
rect 5326 1077 5356 1091
rect 5417 1089 5570 1094
rect 5399 1077 5591 1089
rect 5634 1077 5664 1091
rect 5670 1077 5683 1108
rect 5698 1090 5728 1108
rect 5771 1077 5784 1108
rect 5814 1077 5827 1108
rect 5842 1090 5872 1108
rect 5916 1091 5929 1108
rect 5965 1094 6185 1108
rect 5882 1079 5897 1091
rect 5879 1077 5901 1079
rect 5906 1077 5936 1091
rect 5997 1089 6150 1094
rect 5979 1077 6171 1089
rect 6214 1077 6244 1091
rect 6250 1077 6263 1108
rect 6278 1090 6308 1108
rect 6351 1077 6364 1108
rect 6394 1077 6407 1108
rect 6422 1090 6452 1108
rect 6496 1091 6509 1108
rect 6545 1094 6765 1108
rect 6462 1079 6477 1091
rect 6459 1077 6481 1079
rect 6486 1077 6516 1091
rect 6577 1089 6730 1094
rect 6559 1077 6751 1089
rect 6794 1077 6824 1091
rect 6830 1077 6843 1108
rect 6858 1090 6888 1108
rect 6931 1077 6944 1108
rect 3481 1064 6944 1077
rect 14 960 27 1064
rect 72 1042 73 1052
rect 88 1042 101 1052
rect 72 1038 101 1042
rect 106 1038 136 1064
rect 154 1050 170 1052
rect 242 1050 295 1064
rect 243 1048 307 1050
rect 350 1048 365 1064
rect 414 1061 444 1064
rect 414 1058 450 1061
rect 380 1050 396 1052
rect 154 1038 169 1042
rect 72 1036 169 1038
rect 197 1036 365 1048
rect 381 1038 396 1042
rect 414 1039 453 1058
rect 472 1052 479 1053
rect 478 1045 479 1052
rect 462 1042 463 1045
rect 478 1042 491 1045
rect 414 1038 444 1039
rect 453 1038 459 1039
rect 462 1038 491 1042
rect 381 1037 491 1038
rect 381 1036 497 1037
rect 56 1028 107 1036
rect 56 1016 81 1028
rect 88 1016 107 1028
rect 138 1028 188 1036
rect 138 1020 154 1028
rect 161 1026 188 1028
rect 197 1026 418 1036
rect 161 1016 418 1026
rect 447 1028 497 1036
rect 447 1019 463 1028
rect 56 1008 107 1016
rect 154 1008 418 1016
rect 444 1016 463 1019
rect 470 1016 497 1028
rect 444 1008 497 1016
rect 72 1000 73 1008
rect 88 1000 101 1008
rect 72 992 88 1000
rect 69 985 88 988
rect 69 976 91 985
rect 42 966 91 976
rect 42 960 72 966
rect 91 961 96 966
rect 14 944 88 960
rect 106 952 136 1008
rect 171 998 379 1008
rect 414 1004 459 1008
rect 462 1007 463 1008
rect 478 1007 491 1008
rect 197 968 386 998
rect 212 965 386 968
rect 205 962 386 965
rect 14 942 27 944
rect 42 942 76 944
rect 14 926 88 942
rect 115 938 128 952
rect 143 938 159 954
rect 205 949 216 962
rect -2 904 -1 920
rect 14 904 27 926
rect 42 904 72 926
rect 115 922 177 938
rect 205 931 216 947
rect 221 942 231 962
rect 241 942 255 962
rect 258 949 267 962
rect 283 949 292 962
rect 221 931 255 942
rect 258 931 267 947
rect 283 931 292 947
rect 299 942 309 962
rect 319 942 333 962
rect 334 949 345 962
rect 299 931 333 942
rect 334 931 345 947
rect 391 938 407 954
rect 414 952 444 1004
rect 478 1000 479 1007
rect 463 992 479 1000
rect 450 960 463 979
rect 478 960 508 976
rect 450 944 524 960
rect 450 942 463 944
rect 478 942 512 944
rect 115 920 128 922
rect 143 920 177 922
rect 115 904 177 920
rect 221 915 237 922
rect 299 915 329 926
rect 377 922 423 938
rect 450 926 524 942
rect 377 920 411 922
rect 376 904 423 920
rect 450 904 463 926
rect 478 904 508 926
rect 535 904 536 920
rect 551 904 564 1064
rect 594 960 607 1064
rect 652 1042 653 1052
rect 668 1042 681 1052
rect 652 1038 681 1042
rect 686 1038 716 1064
rect 734 1050 750 1052
rect 822 1050 875 1064
rect 823 1048 887 1050
rect 930 1048 945 1064
rect 994 1061 1024 1064
rect 994 1058 1030 1061
rect 960 1050 976 1052
rect 734 1038 749 1042
rect 652 1036 749 1038
rect 777 1036 945 1048
rect 961 1038 976 1042
rect 994 1039 1033 1058
rect 1052 1052 1059 1053
rect 1058 1045 1059 1052
rect 1042 1042 1043 1045
rect 1058 1042 1071 1045
rect 994 1038 1024 1039
rect 1033 1038 1039 1039
rect 1042 1038 1071 1042
rect 961 1037 1071 1038
rect 961 1036 1077 1037
rect 636 1028 687 1036
rect 636 1016 661 1028
rect 668 1016 687 1028
rect 718 1028 768 1036
rect 718 1020 734 1028
rect 741 1026 768 1028
rect 777 1026 998 1036
rect 741 1016 998 1026
rect 1027 1028 1077 1036
rect 1027 1019 1043 1028
rect 636 1008 687 1016
rect 734 1008 998 1016
rect 1024 1016 1043 1019
rect 1050 1016 1077 1028
rect 1024 1008 1077 1016
rect 652 1000 653 1008
rect 668 1000 681 1008
rect 652 992 668 1000
rect 649 985 668 988
rect 649 976 671 985
rect 622 966 671 976
rect 622 960 652 966
rect 671 961 676 966
rect 594 944 668 960
rect 686 952 716 1008
rect 751 998 959 1008
rect 994 1004 1039 1008
rect 1042 1007 1043 1008
rect 1058 1007 1071 1008
rect 777 968 966 998
rect 792 965 966 968
rect 785 962 966 965
rect 594 942 607 944
rect 622 942 656 944
rect 594 926 668 942
rect 695 938 708 952
rect 723 938 739 954
rect 785 949 796 962
rect 578 904 579 920
rect 594 904 607 926
rect 622 904 652 926
rect 695 922 757 938
rect 785 931 796 947
rect 801 942 811 962
rect 821 942 835 962
rect 838 949 847 962
rect 863 949 872 962
rect 801 931 835 942
rect 838 931 847 947
rect 863 931 872 947
rect 879 942 889 962
rect 899 942 913 962
rect 914 949 925 962
rect 879 931 913 942
rect 914 931 925 947
rect 971 938 987 954
rect 994 952 1024 1004
rect 1058 1000 1059 1007
rect 1043 992 1059 1000
rect 1030 960 1043 979
rect 1058 960 1088 976
rect 1030 944 1104 960
rect 1030 942 1043 944
rect 1058 942 1092 944
rect 695 920 708 922
rect 723 920 757 922
rect 695 904 757 920
rect 801 915 817 922
rect 879 915 909 926
rect 957 922 1003 938
rect 1030 926 1104 942
rect 957 920 991 922
rect 956 904 1003 920
rect 1030 904 1043 926
rect 1058 904 1088 926
rect 1115 904 1116 920
rect 1131 904 1144 1064
rect 1174 960 1187 1064
rect 1232 1042 1233 1052
rect 1248 1042 1261 1052
rect 1232 1038 1261 1042
rect 1266 1038 1296 1064
rect 1314 1050 1330 1052
rect 1402 1050 1455 1064
rect 1403 1048 1467 1050
rect 1510 1048 1525 1064
rect 1574 1061 1604 1064
rect 1574 1058 1610 1061
rect 1540 1050 1556 1052
rect 1314 1038 1329 1042
rect 1232 1036 1329 1038
rect 1357 1036 1525 1048
rect 1541 1038 1556 1042
rect 1574 1039 1613 1058
rect 1632 1052 1639 1053
rect 1638 1045 1639 1052
rect 1622 1042 1623 1045
rect 1638 1042 1651 1045
rect 1574 1038 1604 1039
rect 1613 1038 1619 1039
rect 1622 1038 1651 1042
rect 1541 1037 1651 1038
rect 1541 1036 1657 1037
rect 1216 1028 1267 1036
rect 1216 1016 1241 1028
rect 1248 1016 1267 1028
rect 1298 1028 1348 1036
rect 1298 1020 1314 1028
rect 1321 1026 1348 1028
rect 1357 1026 1578 1036
rect 1321 1016 1578 1026
rect 1607 1028 1657 1036
rect 1607 1019 1623 1028
rect 1216 1008 1267 1016
rect 1314 1008 1578 1016
rect 1604 1016 1623 1019
rect 1630 1016 1657 1028
rect 1604 1008 1657 1016
rect 1232 1000 1233 1008
rect 1248 1000 1261 1008
rect 1232 992 1248 1000
rect 1229 985 1248 988
rect 1229 976 1251 985
rect 1202 966 1251 976
rect 1202 960 1232 966
rect 1251 961 1256 966
rect 1174 944 1248 960
rect 1266 952 1296 1008
rect 1331 998 1539 1008
rect 1574 1004 1619 1008
rect 1622 1007 1623 1008
rect 1638 1007 1651 1008
rect 1357 968 1546 998
rect 1372 965 1546 968
rect 1365 962 1546 965
rect 1174 942 1187 944
rect 1202 942 1236 944
rect 1174 926 1248 942
rect 1275 938 1288 952
rect 1303 938 1319 954
rect 1365 949 1376 962
rect 1158 904 1159 920
rect 1174 904 1187 926
rect 1202 904 1232 926
rect 1275 922 1337 938
rect 1365 931 1376 947
rect 1381 942 1391 962
rect 1401 942 1415 962
rect 1418 949 1427 962
rect 1443 949 1452 962
rect 1381 931 1415 942
rect 1418 931 1427 947
rect 1443 931 1452 947
rect 1459 942 1469 962
rect 1479 942 1493 962
rect 1494 949 1505 962
rect 1459 931 1493 942
rect 1494 931 1505 947
rect 1551 938 1567 954
rect 1574 952 1604 1004
rect 1638 1000 1639 1007
rect 1623 992 1639 1000
rect 1610 960 1623 979
rect 1638 960 1668 976
rect 1610 944 1684 960
rect 1610 942 1623 944
rect 1638 942 1672 944
rect 1275 920 1288 922
rect 1303 920 1337 922
rect 1275 904 1337 920
rect 1381 915 1397 922
rect 1459 915 1489 926
rect 1537 922 1583 938
rect 1610 926 1684 942
rect 1537 920 1571 922
rect 1536 904 1583 920
rect 1610 904 1623 926
rect 1638 904 1668 926
rect 1695 904 1696 920
rect 1711 904 1724 1064
rect 1754 960 1767 1064
rect 1812 1042 1813 1052
rect 1828 1042 1837 1052
rect 1812 1036 1837 1042
rect 1796 1028 1837 1036
rect 1796 1016 1821 1028
rect 1828 1016 1837 1028
rect 1796 1008 1837 1016
rect 1812 1000 1813 1008
rect 1828 1000 1837 1008
rect 1812 992 1828 1000
rect 1809 985 1828 988
rect 1809 976 1831 985
rect 1782 966 1831 976
rect 1782 960 1812 966
rect 1831 961 1836 966
rect 3494 960 3507 1064
rect 3552 1042 3553 1052
rect 3568 1042 3581 1052
rect 3552 1038 3581 1042
rect 3586 1038 3616 1064
rect 3634 1050 3650 1052
rect 3722 1050 3775 1064
rect 3723 1048 3787 1050
rect 3830 1048 3845 1064
rect 3894 1061 3924 1064
rect 3894 1058 3930 1061
rect 3860 1050 3876 1052
rect 3634 1038 3649 1042
rect 3552 1036 3649 1038
rect 3677 1036 3845 1048
rect 3861 1038 3876 1042
rect 3894 1039 3933 1058
rect 3952 1052 3959 1053
rect 3958 1045 3959 1052
rect 3942 1042 3943 1045
rect 3958 1042 3971 1045
rect 3894 1038 3924 1039
rect 3933 1038 3939 1039
rect 3942 1038 3971 1042
rect 3861 1037 3971 1038
rect 3861 1036 3977 1037
rect 3536 1028 3587 1036
rect 3536 1016 3561 1028
rect 3568 1016 3587 1028
rect 3618 1028 3668 1036
rect 3618 1020 3634 1028
rect 3641 1026 3668 1028
rect 3677 1026 3898 1036
rect 3641 1016 3898 1026
rect 3927 1028 3977 1036
rect 3927 1019 3943 1028
rect 3536 1008 3587 1016
rect 3634 1008 3898 1016
rect 3924 1016 3943 1019
rect 3950 1016 3977 1028
rect 3924 1008 3977 1016
rect 3552 1000 3553 1008
rect 3568 1000 3581 1008
rect 3552 992 3568 1000
rect 3549 985 3568 988
rect 3549 976 3571 985
rect 3522 966 3571 976
rect 3522 960 3552 966
rect 3571 961 3576 966
rect 1754 944 1828 960
rect 3494 944 3568 960
rect 3586 952 3616 1008
rect 3651 998 3859 1008
rect 3894 1004 3939 1008
rect 3942 1007 3943 1008
rect 3958 1007 3971 1008
rect 3677 968 3866 998
rect 3692 965 3866 968
rect 3685 962 3866 965
rect 1754 942 1767 944
rect 1782 942 1816 944
rect 3494 942 3507 944
rect 3522 942 3556 944
rect 1754 926 1828 942
rect 3494 926 3568 942
rect 3595 938 3608 952
rect 3623 938 3639 954
rect 3685 949 3696 962
rect 1738 904 1739 920
rect 1754 904 1767 926
rect 1782 904 1812 926
rect 3494 914 3507 926
rect 3522 914 3552 926
rect 3595 922 3657 938
rect 3685 931 3696 947
rect 3701 942 3711 962
rect 3721 942 3735 962
rect 3738 949 3747 962
rect 3763 949 3772 962
rect 3701 931 3735 942
rect 3738 931 3747 947
rect 3763 931 3772 947
rect 3779 942 3789 962
rect 3799 942 3813 962
rect 3814 949 3825 962
rect 3779 931 3813 942
rect 3814 931 3825 947
rect 3871 938 3887 954
rect 3894 952 3924 1004
rect 3958 1000 3959 1007
rect 3943 992 3959 1000
rect 3930 960 3943 979
rect 3958 960 3988 976
rect 3930 944 4004 960
rect 3930 942 3943 944
rect 3958 942 3992 944
rect 3595 920 3608 922
rect 3623 920 3657 922
rect 3595 914 3657 920
rect 3701 915 3717 922
rect 3779 915 3809 926
rect 3857 922 3903 938
rect 3930 926 4004 942
rect 3857 920 3891 922
rect 3857 914 3903 920
rect 3930 914 3943 926
rect 3958 914 3988 926
rect 4031 914 4044 1064
rect 4074 960 4087 1064
rect 4132 1042 4133 1052
rect 4148 1042 4161 1052
rect 4132 1038 4161 1042
rect 4166 1038 4196 1064
rect 4214 1050 4230 1052
rect 4302 1050 4355 1064
rect 4303 1048 4367 1050
rect 4410 1048 4425 1064
rect 4474 1061 4504 1064
rect 4611 1063 6944 1064
rect 4474 1058 4510 1061
rect 4440 1050 4456 1052
rect 4214 1038 4229 1042
rect 4132 1036 4229 1038
rect 4257 1036 4425 1048
rect 4441 1038 4456 1042
rect 4474 1039 4513 1058
rect 4532 1052 4539 1053
rect 4538 1045 4539 1052
rect 4522 1042 4523 1045
rect 4538 1042 4551 1045
rect 4474 1038 4504 1039
rect 4513 1038 4519 1039
rect 4522 1038 4551 1042
rect 4441 1037 4551 1038
rect 4441 1036 4557 1037
rect 4116 1028 4167 1036
rect 4116 1016 4141 1028
rect 4148 1016 4167 1028
rect 4198 1028 4248 1036
rect 4198 1020 4214 1028
rect 4221 1026 4248 1028
rect 4257 1026 4478 1036
rect 4221 1016 4478 1026
rect 4507 1028 4557 1036
rect 4507 1019 4523 1028
rect 4116 1008 4167 1016
rect 4214 1008 4478 1016
rect 4504 1016 4523 1019
rect 4530 1016 4557 1028
rect 4504 1008 4557 1016
rect 4132 1000 4133 1008
rect 4148 1000 4161 1008
rect 4132 992 4148 1000
rect 4129 985 4148 988
rect 4129 976 4151 985
rect 4102 966 4151 976
rect 4102 960 4132 966
rect 4151 961 4156 966
rect 4074 944 4148 960
rect 4166 952 4196 1008
rect 4231 998 4439 1008
rect 4474 1004 4519 1008
rect 4522 1007 4523 1008
rect 4538 1007 4551 1008
rect 4257 968 4446 998
rect 4272 965 4446 968
rect 4265 962 4446 965
rect 4074 942 4087 944
rect 4102 942 4136 944
rect 4074 926 4148 942
rect 4175 938 4188 952
rect 4203 938 4219 954
rect 4265 949 4276 962
rect 4074 914 4087 926
rect 4102 914 4132 926
rect 4175 922 4237 938
rect 4265 931 4276 947
rect 4281 942 4291 962
rect 4301 942 4315 962
rect 4318 949 4327 962
rect 4343 949 4352 962
rect 4281 931 4315 942
rect 4318 931 4327 947
rect 4343 931 4352 947
rect 4359 942 4369 962
rect 4379 942 4393 962
rect 4394 949 4405 962
rect 4359 931 4393 942
rect 4394 931 4405 947
rect 4451 938 4467 954
rect 4474 952 4504 1004
rect 4538 1000 4539 1007
rect 4523 992 4539 1000
rect 4510 960 4523 979
rect 4538 960 4568 976
rect 4510 944 4584 960
rect 4510 942 4523 944
rect 4538 942 4572 944
rect 4175 920 4188 922
rect 4203 920 4237 922
rect 4175 914 4237 920
rect 4281 915 4297 922
rect 4359 915 4389 926
rect 4437 922 4483 938
rect 4510 926 4584 942
rect 4437 920 4471 922
rect 4437 914 4483 920
rect 4510 914 4523 926
rect 4538 914 4568 926
rect 4611 914 4624 1063
rect 4654 959 4667 1063
rect 4712 1041 4713 1051
rect 4728 1041 4741 1051
rect 4712 1037 4741 1041
rect 4746 1037 4776 1063
rect 4794 1049 4810 1051
rect 4882 1049 4935 1063
rect 4883 1047 4947 1049
rect 4990 1047 5005 1063
rect 5054 1060 5084 1063
rect 5054 1057 5090 1060
rect 5020 1049 5036 1051
rect 4794 1037 4809 1041
rect 4712 1035 4809 1037
rect 4837 1035 5005 1047
rect 5021 1037 5036 1041
rect 5054 1038 5093 1057
rect 5112 1051 5119 1052
rect 5118 1044 5119 1051
rect 5102 1041 5103 1044
rect 5118 1041 5131 1044
rect 5054 1037 5084 1038
rect 5093 1037 5099 1038
rect 5102 1037 5131 1041
rect 5021 1036 5131 1037
rect 5021 1035 5137 1036
rect 4696 1027 4747 1035
rect 4696 1015 4721 1027
rect 4728 1015 4747 1027
rect 4778 1027 4828 1035
rect 4778 1019 4794 1027
rect 4801 1025 4828 1027
rect 4837 1025 5058 1035
rect 4801 1015 5058 1025
rect 5087 1027 5137 1035
rect 5087 1018 5103 1027
rect 4696 1007 4747 1015
rect 4794 1007 5058 1015
rect 5084 1015 5103 1018
rect 5110 1015 5137 1027
rect 5084 1007 5137 1015
rect 4712 999 4713 1007
rect 4728 999 4741 1007
rect 4712 991 4728 999
rect 4709 984 4728 987
rect 4709 975 4731 984
rect 4682 965 4731 975
rect 4682 959 4712 965
rect 4731 960 4736 965
rect 4654 943 4728 959
rect 4746 951 4776 1007
rect 4811 997 5019 1007
rect 5054 1003 5099 1007
rect 5102 1006 5103 1007
rect 5118 1006 5131 1007
rect 4837 967 5026 997
rect 4852 964 5026 967
rect 4845 961 5026 964
rect 4654 941 4667 943
rect 4682 941 4716 943
rect 4654 925 4728 941
rect 4755 937 4768 951
rect 4783 937 4799 953
rect 4845 948 4856 961
rect 4654 914 4667 925
rect 4682 914 4712 925
rect 4755 921 4817 937
rect 4845 930 4856 946
rect 4861 941 4871 961
rect 4881 941 4895 961
rect 4898 948 4907 961
rect 4923 948 4932 961
rect 4861 930 4895 941
rect 4898 930 4907 946
rect 4923 930 4932 946
rect 4939 941 4949 961
rect 4959 941 4973 961
rect 4974 948 4985 961
rect 4939 930 4973 941
rect 4974 930 4985 946
rect 5031 937 5047 953
rect 5054 951 5084 1003
rect 5118 999 5119 1006
rect 5103 991 5119 999
rect 5090 959 5103 978
rect 5118 959 5148 975
rect 5090 943 5164 959
rect 5090 941 5103 943
rect 5118 941 5152 943
rect 4755 919 4768 921
rect 4783 919 4817 921
rect 4755 914 4817 919
rect 4861 914 4877 921
rect 4939 914 4969 925
rect 5017 921 5063 937
rect 5090 925 5164 941
rect 5017 919 5051 921
rect 5017 914 5063 919
rect 5090 914 5103 925
rect 5118 914 5148 925
rect 5191 914 5204 1063
rect 5234 959 5247 1063
rect 5292 1041 5293 1051
rect 5308 1041 5321 1051
rect 5292 1037 5321 1041
rect 5326 1037 5356 1063
rect 5374 1049 5390 1051
rect 5462 1049 5515 1063
rect 5463 1047 5527 1049
rect 5570 1047 5585 1063
rect 5634 1060 5664 1063
rect 5634 1057 5670 1060
rect 5600 1049 5616 1051
rect 5374 1037 5389 1041
rect 5292 1035 5389 1037
rect 5417 1035 5585 1047
rect 5601 1037 5616 1041
rect 5634 1038 5673 1057
rect 5692 1051 5699 1052
rect 5698 1044 5699 1051
rect 5682 1041 5683 1044
rect 5698 1041 5711 1044
rect 5634 1037 5664 1038
rect 5673 1037 5679 1038
rect 5682 1037 5711 1041
rect 5601 1036 5711 1037
rect 5601 1035 5717 1036
rect 5276 1027 5327 1035
rect 5276 1015 5301 1027
rect 5308 1015 5327 1027
rect 5358 1027 5408 1035
rect 5358 1019 5374 1027
rect 5381 1025 5408 1027
rect 5417 1025 5638 1035
rect 5381 1015 5638 1025
rect 5667 1027 5717 1035
rect 5667 1018 5683 1027
rect 5276 1007 5327 1015
rect 5374 1007 5638 1015
rect 5664 1015 5683 1018
rect 5690 1015 5717 1027
rect 5664 1007 5717 1015
rect 5292 999 5293 1007
rect 5308 999 5321 1007
rect 5292 991 5308 999
rect 5289 984 5308 987
rect 5289 975 5311 984
rect 5262 965 5311 975
rect 5262 959 5292 965
rect 5311 960 5316 965
rect 5234 943 5308 959
rect 5326 951 5356 1007
rect 5391 997 5599 1007
rect 5634 1003 5679 1007
rect 5682 1006 5683 1007
rect 5698 1006 5711 1007
rect 5417 967 5606 997
rect 5432 964 5606 967
rect 5425 961 5606 964
rect 5234 941 5247 943
rect 5262 941 5296 943
rect 5234 925 5308 941
rect 5335 937 5348 951
rect 5363 937 5379 953
rect 5425 948 5436 961
rect 5234 914 5247 925
rect 5262 914 5292 925
rect 5335 921 5397 937
rect 5425 930 5436 946
rect 5441 941 5451 961
rect 5461 941 5475 961
rect 5478 948 5487 961
rect 5503 948 5512 961
rect 5441 930 5475 941
rect 5478 930 5487 946
rect 5503 930 5512 946
rect 5519 941 5529 961
rect 5539 941 5553 961
rect 5554 948 5565 961
rect 5519 930 5553 941
rect 5554 930 5565 946
rect 5611 937 5627 953
rect 5634 951 5664 1003
rect 5698 999 5699 1006
rect 5683 991 5699 999
rect 5670 959 5683 978
rect 5698 959 5728 975
rect 5670 943 5744 959
rect 5670 941 5683 943
rect 5698 941 5732 943
rect 5335 919 5348 921
rect 5363 919 5397 921
rect 5335 914 5397 919
rect 5441 914 5457 921
rect 5519 914 5549 925
rect 5597 921 5643 937
rect 5670 925 5744 941
rect 5597 919 5631 921
rect 5597 914 5643 919
rect 5670 914 5683 925
rect 5698 914 5728 925
rect 5771 914 5784 1063
rect 5814 959 5827 1063
rect 5872 1041 5873 1051
rect 5888 1041 5901 1051
rect 5872 1037 5901 1041
rect 5906 1037 5936 1063
rect 5954 1049 5970 1051
rect 6042 1049 6095 1063
rect 6043 1047 6107 1049
rect 6150 1047 6165 1063
rect 6214 1060 6244 1063
rect 6214 1057 6250 1060
rect 6180 1049 6196 1051
rect 5954 1037 5969 1041
rect 5872 1035 5969 1037
rect 5997 1035 6165 1047
rect 6181 1037 6196 1041
rect 6214 1038 6253 1057
rect 6272 1051 6279 1052
rect 6278 1044 6279 1051
rect 6262 1041 6263 1044
rect 6278 1041 6291 1044
rect 6214 1037 6244 1038
rect 6253 1037 6259 1038
rect 6262 1037 6291 1041
rect 6181 1036 6291 1037
rect 6181 1035 6297 1036
rect 5856 1027 5907 1035
rect 5856 1015 5881 1027
rect 5888 1015 5907 1027
rect 5938 1027 5988 1035
rect 5938 1019 5954 1027
rect 5961 1025 5988 1027
rect 5997 1025 6218 1035
rect 5961 1015 6218 1025
rect 6247 1027 6297 1035
rect 6247 1018 6263 1027
rect 5856 1007 5907 1015
rect 5954 1007 6218 1015
rect 6244 1015 6263 1018
rect 6270 1015 6297 1027
rect 6244 1007 6297 1015
rect 5872 999 5873 1007
rect 5888 999 5901 1007
rect 5872 991 5888 999
rect 5869 984 5888 987
rect 5869 975 5891 984
rect 5842 965 5891 975
rect 5842 959 5872 965
rect 5891 960 5896 965
rect 5814 943 5888 959
rect 5906 951 5936 1007
rect 5971 997 6179 1007
rect 6214 1003 6259 1007
rect 6262 1006 6263 1007
rect 6278 1006 6291 1007
rect 5997 967 6186 997
rect 6012 964 6186 967
rect 6005 961 6186 964
rect 5814 941 5827 943
rect 5842 941 5876 943
rect 5814 925 5888 941
rect 5915 937 5928 951
rect 5943 937 5959 953
rect 6005 948 6016 961
rect 5814 914 5827 925
rect 5842 914 5872 925
rect 5915 921 5977 937
rect 6005 930 6016 946
rect 6021 941 6031 961
rect 6041 941 6055 961
rect 6058 948 6067 961
rect 6083 948 6092 961
rect 6021 930 6055 941
rect 6058 930 6067 946
rect 6083 930 6092 946
rect 6099 941 6109 961
rect 6119 941 6133 961
rect 6134 948 6145 961
rect 6099 930 6133 941
rect 6134 930 6145 946
rect 6191 937 6207 953
rect 6214 951 6244 1003
rect 6278 999 6279 1006
rect 6263 991 6279 999
rect 6250 959 6263 978
rect 6278 959 6308 975
rect 6250 943 6324 959
rect 6250 941 6263 943
rect 6278 941 6312 943
rect 5915 919 5928 921
rect 5943 919 5977 921
rect 5915 914 5977 919
rect 6021 914 6037 921
rect 6099 914 6129 925
rect 6177 921 6223 937
rect 6250 925 6324 941
rect 6177 919 6211 921
rect 6177 914 6223 919
rect 6250 914 6263 925
rect 6278 914 6308 925
rect 6351 914 6364 1063
rect 6394 959 6407 1063
rect 6452 1041 6453 1051
rect 6468 1041 6481 1051
rect 6452 1037 6481 1041
rect 6486 1037 6516 1063
rect 6534 1049 6550 1051
rect 6622 1049 6675 1063
rect 6623 1047 6687 1049
rect 6730 1047 6745 1063
rect 6794 1060 6824 1063
rect 6794 1057 6830 1060
rect 6760 1049 6776 1051
rect 6534 1037 6549 1041
rect 6452 1035 6549 1037
rect 6577 1035 6745 1047
rect 6761 1037 6776 1041
rect 6794 1038 6833 1057
rect 6852 1051 6859 1052
rect 6858 1044 6859 1051
rect 6842 1041 6843 1044
rect 6858 1041 6871 1044
rect 6794 1037 6824 1038
rect 6833 1037 6839 1038
rect 6842 1037 6871 1041
rect 6761 1036 6871 1037
rect 6761 1035 6877 1036
rect 6436 1027 6487 1035
rect 6436 1015 6461 1027
rect 6468 1015 6487 1027
rect 6518 1027 6568 1035
rect 6518 1019 6534 1027
rect 6541 1025 6568 1027
rect 6577 1025 6798 1035
rect 6541 1015 6798 1025
rect 6827 1027 6877 1035
rect 6827 1018 6843 1027
rect 6436 1007 6487 1015
rect 6534 1007 6798 1015
rect 6824 1015 6843 1018
rect 6850 1015 6877 1027
rect 6824 1007 6877 1015
rect 6452 999 6453 1007
rect 6468 999 6481 1007
rect 6452 991 6468 999
rect 6449 984 6468 987
rect 6449 975 6471 984
rect 6422 965 6471 975
rect 6422 959 6452 965
rect 6471 960 6476 965
rect 6394 943 6468 959
rect 6486 951 6516 1007
rect 6551 997 6759 1007
rect 6794 1003 6839 1007
rect 6842 1006 6843 1007
rect 6858 1006 6871 1007
rect 6577 967 6766 997
rect 6592 964 6766 967
rect 6585 961 6766 964
rect 6394 941 6407 943
rect 6422 941 6456 943
rect 6394 925 6468 941
rect 6495 937 6508 951
rect 6523 937 6539 953
rect 6585 948 6596 961
rect 6394 914 6407 925
rect 6422 914 6452 925
rect 6495 921 6557 937
rect 6585 930 6596 946
rect 6601 941 6611 961
rect 6621 941 6635 961
rect 6638 948 6647 961
rect 6663 948 6672 961
rect 6601 930 6635 941
rect 6638 930 6647 946
rect 6663 930 6672 946
rect 6679 941 6689 961
rect 6699 941 6713 961
rect 6714 948 6725 961
rect 6679 930 6713 941
rect 6714 930 6725 946
rect 6771 937 6787 953
rect 6794 951 6824 1003
rect 6858 999 6859 1006
rect 6843 991 6859 999
rect 6830 959 6843 978
rect 6858 959 6888 975
rect 6830 943 6904 959
rect 6830 941 6843 943
rect 6858 941 6892 943
rect 6495 919 6508 921
rect 6523 919 6557 921
rect 6495 914 6557 919
rect 6601 914 6617 921
rect 6679 914 6709 925
rect 6757 921 6803 937
rect 6830 925 6904 941
rect 6757 919 6791 921
rect 6757 914 6803 919
rect 6830 914 6843 925
rect 6858 914 6888 925
rect 6931 914 6944 1063
rect -8 896 33 904
rect -8 870 7 896
rect 14 870 33 896
rect 97 892 159 904
rect 171 892 246 904
rect 304 892 379 904
rect 391 892 422 904
rect 428 892 463 904
rect 97 890 259 892
rect -8 862 33 870
rect 115 866 128 890
rect 143 888 158 890
rect -2 852 -1 862
rect 14 852 27 862
rect 42 852 72 866
rect 115 852 158 866
rect 182 863 189 870
rect 192 866 259 890
rect 291 890 463 892
rect 261 868 289 872
rect 291 868 371 890
rect 392 888 407 890
rect 261 866 371 868
rect 192 862 371 866
rect 165 852 195 862
rect 197 852 350 862
rect 358 852 388 862
rect 392 852 422 866
rect 450 852 463 890
rect 535 896 570 904
rect 535 870 536 896
rect 543 870 570 896
rect 478 852 508 866
rect 535 862 570 870
rect 572 896 613 904
rect 572 870 587 896
rect 594 870 613 896
rect 677 892 739 904
rect 751 892 826 904
rect 884 892 959 904
rect 971 892 1002 904
rect 1008 892 1043 904
rect 677 890 839 892
rect 572 862 613 870
rect 695 866 708 890
rect 723 888 738 890
rect 535 852 536 862
rect 551 852 564 862
rect 578 852 579 862
rect 594 852 607 862
rect 622 852 652 866
rect 695 852 738 866
rect 762 863 769 870
rect 772 866 839 890
rect 871 890 1043 892
rect 841 868 869 872
rect 871 868 951 890
rect 972 888 987 890
rect 841 866 951 868
rect 772 862 951 866
rect 745 852 775 862
rect 777 852 930 862
rect 938 852 968 862
rect 972 852 1002 866
rect 1030 852 1043 890
rect 1115 896 1150 904
rect 1115 870 1116 896
rect 1123 870 1150 896
rect 1058 852 1088 866
rect 1115 862 1150 870
rect 1152 896 1193 904
rect 1152 870 1167 896
rect 1174 870 1193 896
rect 1257 892 1319 904
rect 1331 892 1406 904
rect 1464 892 1539 904
rect 1551 892 1582 904
rect 1588 892 1623 904
rect 1257 890 1419 892
rect 1152 862 1193 870
rect 1275 866 1288 890
rect 1303 888 1318 890
rect 1115 852 1116 862
rect 1131 852 1144 862
rect 1158 852 1159 862
rect 1174 852 1187 862
rect 1202 852 1232 866
rect 1275 852 1318 866
rect 1342 863 1349 870
rect 1352 866 1419 890
rect 1451 890 1623 892
rect 1421 868 1449 872
rect 1451 868 1531 890
rect 1552 888 1567 890
rect 1421 866 1531 868
rect 1352 862 1531 866
rect 1325 852 1355 862
rect 1357 852 1510 862
rect 1518 852 1548 862
rect 1552 852 1582 866
rect 1610 852 1623 890
rect 1695 896 1730 904
rect 1695 870 1696 896
rect 1703 870 1730 896
rect 1638 852 1668 866
rect 1695 862 1730 870
rect 1732 896 1773 904
rect 1732 870 1747 896
rect 1754 870 1773 896
rect 1732 862 1773 870
rect 1695 852 1696 862
rect 1711 852 1724 862
rect 1738 852 1739 862
rect 1754 852 1767 862
rect 1782 852 1812 866
rect -2 846 1837 852
rect -1 838 1837 846
rect 14 808 27 838
rect 42 820 72 838
rect 115 824 129 838
rect 165 824 385 838
rect 116 822 129 824
rect 82 810 97 822
rect 79 808 101 810
rect 106 808 136 822
rect 197 820 350 824
rect 179 808 371 820
rect 414 808 444 822
rect 450 808 463 838
rect 478 820 508 838
rect 551 808 564 838
rect 594 808 607 838
rect 622 820 652 838
rect 695 824 709 838
rect 745 824 965 838
rect 696 822 709 824
rect 662 810 677 822
rect 659 808 681 810
rect 686 808 716 822
rect 777 820 930 824
rect 759 808 951 820
rect 994 808 1024 822
rect 1030 808 1043 838
rect 1058 820 1088 838
rect 1131 808 1144 838
rect 1174 808 1187 838
rect 1202 820 1232 838
rect 1275 824 1289 838
rect 1325 824 1545 838
rect 1276 822 1289 824
rect 1242 810 1257 822
rect 1239 808 1261 810
rect 1266 808 1296 822
rect 1357 820 1510 824
rect 1339 808 1531 820
rect 1574 808 1604 822
rect 1610 808 1623 838
rect 1638 820 1668 838
rect 1711 808 1724 838
rect 1754 808 1767 838
rect 1782 820 1812 838
rect 1822 810 1837 822
rect 1819 808 1837 810
rect -1 794 1837 808
rect 14 690 27 794
rect 72 772 73 782
rect 88 772 101 782
rect 72 768 101 772
rect 106 768 136 794
rect 154 780 170 782
rect 242 780 295 794
rect 243 778 307 780
rect 350 778 365 794
rect 414 791 444 794
rect 414 788 450 791
rect 380 780 396 782
rect 154 768 169 772
rect 72 766 169 768
rect 197 766 365 778
rect 381 768 396 772
rect 414 769 453 788
rect 472 782 479 783
rect 478 775 479 782
rect 462 772 463 775
rect 478 772 491 775
rect 414 768 444 769
rect 453 768 459 769
rect 462 768 491 772
rect 381 767 491 768
rect 381 766 497 767
rect 56 758 107 766
rect 56 746 81 758
rect 88 746 107 758
rect 138 758 188 766
rect 138 750 154 758
rect 161 756 188 758
rect 197 756 418 766
rect 161 746 418 756
rect 447 758 497 766
rect 447 749 463 758
rect 56 738 107 746
rect 154 738 418 746
rect 444 746 463 749
rect 470 746 497 758
rect 444 738 497 746
rect 72 730 73 738
rect 88 730 101 738
rect 72 722 88 730
rect 69 715 88 718
rect 69 706 91 715
rect 42 696 91 706
rect 42 690 72 696
rect 91 691 96 696
rect 14 674 88 690
rect 106 682 136 738
rect 171 728 379 738
rect 414 734 459 738
rect 462 737 463 738
rect 478 737 491 738
rect 197 698 386 728
rect 212 695 386 698
rect 205 692 386 695
rect 14 672 27 674
rect 42 672 76 674
rect 14 656 88 672
rect 115 668 128 682
rect 143 668 159 684
rect 205 679 216 692
rect -2 634 -1 650
rect 14 634 27 656
rect 42 634 72 656
rect 115 652 177 668
rect 205 661 216 677
rect 221 672 231 692
rect 241 672 255 692
rect 258 679 267 692
rect 283 679 292 692
rect 221 661 255 672
rect 258 661 267 677
rect 283 661 292 677
rect 299 672 309 692
rect 319 672 333 692
rect 334 679 345 692
rect 299 661 333 672
rect 334 661 345 677
rect 391 668 407 684
rect 414 682 444 734
rect 478 730 479 737
rect 463 722 479 730
rect 450 690 463 709
rect 478 690 508 706
rect 450 674 524 690
rect 450 672 463 674
rect 478 672 512 674
rect 115 650 128 652
rect 143 650 177 652
rect 115 634 177 650
rect 221 645 237 652
rect 299 645 329 656
rect 377 652 423 668
rect 450 656 524 672
rect 377 650 411 652
rect 376 634 423 650
rect 450 634 463 656
rect 478 634 508 656
rect 535 634 536 650
rect 551 634 564 794
rect 594 690 607 794
rect 652 772 653 782
rect 668 772 681 782
rect 652 768 681 772
rect 686 768 716 794
rect 734 780 750 782
rect 822 780 875 794
rect 823 778 887 780
rect 930 778 945 794
rect 994 791 1024 794
rect 994 788 1030 791
rect 960 780 976 782
rect 734 768 749 772
rect 652 766 749 768
rect 777 766 945 778
rect 961 768 976 772
rect 994 769 1033 788
rect 1052 782 1059 783
rect 1058 775 1059 782
rect 1042 772 1043 775
rect 1058 772 1071 775
rect 994 768 1024 769
rect 1033 768 1039 769
rect 1042 768 1071 772
rect 961 767 1071 768
rect 961 766 1077 767
rect 636 758 687 766
rect 636 746 661 758
rect 668 746 687 758
rect 718 758 768 766
rect 718 750 734 758
rect 741 756 768 758
rect 777 756 998 766
rect 741 746 998 756
rect 1027 758 1077 766
rect 1027 749 1043 758
rect 636 738 687 746
rect 734 738 998 746
rect 1024 746 1043 749
rect 1050 746 1077 758
rect 1024 738 1077 746
rect 652 730 653 738
rect 668 730 681 738
rect 652 722 668 730
rect 649 715 668 718
rect 649 706 671 715
rect 622 696 671 706
rect 622 690 652 696
rect 671 691 676 696
rect 594 674 668 690
rect 686 682 716 738
rect 751 728 959 738
rect 994 734 1039 738
rect 1042 737 1043 738
rect 1058 737 1071 738
rect 777 698 966 728
rect 792 695 966 698
rect 785 692 966 695
rect 594 672 607 674
rect 622 672 656 674
rect 594 656 668 672
rect 695 668 708 682
rect 723 668 739 684
rect 785 679 796 692
rect 578 634 579 650
rect 594 634 607 656
rect 622 634 652 656
rect 695 652 757 668
rect 785 661 796 677
rect 801 672 811 692
rect 821 672 835 692
rect 838 679 847 692
rect 863 679 872 692
rect 801 661 835 672
rect 838 661 847 677
rect 863 661 872 677
rect 879 672 889 692
rect 899 672 913 692
rect 914 679 925 692
rect 879 661 913 672
rect 914 661 925 677
rect 971 668 987 684
rect 994 682 1024 734
rect 1058 730 1059 737
rect 1043 722 1059 730
rect 1030 690 1043 709
rect 1058 690 1088 706
rect 1030 674 1104 690
rect 1030 672 1043 674
rect 1058 672 1092 674
rect 695 650 708 652
rect 723 650 757 652
rect 695 634 757 650
rect 801 645 817 652
rect 879 645 909 656
rect 957 652 1003 668
rect 1030 656 1104 672
rect 957 650 991 652
rect 956 634 1003 650
rect 1030 634 1043 656
rect 1058 634 1088 656
rect 1115 634 1116 650
rect 1131 634 1144 794
rect 1174 690 1187 794
rect 1232 772 1233 782
rect 1248 772 1261 782
rect 1232 768 1261 772
rect 1266 768 1296 794
rect 1314 780 1330 782
rect 1402 780 1455 794
rect 1403 778 1467 780
rect 1510 778 1525 794
rect 1574 791 1604 794
rect 1574 788 1610 791
rect 1540 780 1556 782
rect 1314 768 1329 772
rect 1232 766 1329 768
rect 1357 766 1525 778
rect 1541 768 1556 772
rect 1574 769 1613 788
rect 1632 782 1639 783
rect 1638 775 1639 782
rect 1622 772 1623 775
rect 1638 772 1651 775
rect 1574 768 1604 769
rect 1613 768 1619 769
rect 1622 768 1651 772
rect 1541 767 1651 768
rect 1541 766 1657 767
rect 1216 758 1267 766
rect 1216 746 1241 758
rect 1248 746 1267 758
rect 1298 758 1348 766
rect 1298 750 1314 758
rect 1321 756 1348 758
rect 1357 756 1578 766
rect 1321 746 1578 756
rect 1607 758 1657 766
rect 1607 749 1623 758
rect 1216 738 1267 746
rect 1314 738 1578 746
rect 1604 746 1623 749
rect 1630 746 1657 758
rect 1604 738 1657 746
rect 1232 730 1233 738
rect 1248 730 1261 738
rect 1232 722 1248 730
rect 1229 715 1248 718
rect 1229 706 1251 715
rect 1202 696 1251 706
rect 1202 690 1232 696
rect 1251 691 1256 696
rect 1174 674 1248 690
rect 1266 682 1296 738
rect 1331 728 1539 738
rect 1574 734 1619 738
rect 1622 737 1623 738
rect 1638 737 1651 738
rect 1357 698 1546 728
rect 1372 695 1546 698
rect 1365 692 1546 695
rect 1174 672 1187 674
rect 1202 672 1236 674
rect 1174 656 1248 672
rect 1275 668 1288 682
rect 1303 668 1319 684
rect 1365 679 1376 692
rect 1158 634 1159 650
rect 1174 634 1187 656
rect 1202 634 1232 656
rect 1275 652 1337 668
rect 1365 661 1376 677
rect 1381 672 1391 692
rect 1401 672 1415 692
rect 1418 679 1427 692
rect 1443 679 1452 692
rect 1381 661 1415 672
rect 1418 661 1427 677
rect 1443 661 1452 677
rect 1459 672 1469 692
rect 1479 672 1493 692
rect 1494 679 1505 692
rect 1459 661 1493 672
rect 1494 661 1505 677
rect 1551 668 1567 684
rect 1574 682 1604 734
rect 1638 730 1639 737
rect 1623 722 1639 730
rect 1610 690 1623 709
rect 1638 690 1668 706
rect 1610 674 1684 690
rect 1610 672 1623 674
rect 1638 672 1672 674
rect 1275 650 1288 652
rect 1303 650 1337 652
rect 1275 634 1337 650
rect 1381 645 1397 652
rect 1459 645 1489 656
rect 1537 652 1583 668
rect 1610 656 1684 672
rect 1537 650 1571 652
rect 1536 634 1583 650
rect 1610 634 1623 656
rect 1638 634 1668 656
rect 1695 634 1696 650
rect 1711 634 1724 794
rect 1754 690 1767 794
rect 1812 772 1813 782
rect 1828 772 1837 782
rect 1812 766 1837 772
rect 1796 758 1837 766
rect 1796 746 1821 758
rect 1828 746 1837 758
rect 1796 738 1837 746
rect 1812 730 1813 738
rect 1828 730 1837 738
rect 1812 722 1828 730
rect 1809 715 1828 718
rect 1809 706 1831 715
rect 1782 696 1831 706
rect 1782 690 1812 696
rect 1831 691 1836 696
rect 1754 674 1828 690
rect 1754 672 1767 674
rect 1782 672 1816 674
rect 1754 656 1828 672
rect 1738 634 1739 650
rect 1754 634 1767 656
rect 1782 634 1812 656
rect -8 626 33 634
rect -8 600 7 626
rect 14 600 33 626
rect 97 622 159 634
rect 171 622 246 634
rect 304 622 379 634
rect 391 622 422 634
rect 428 622 463 634
rect 97 620 259 622
rect -8 592 33 600
rect 115 596 128 620
rect 143 618 158 620
rect -2 582 -1 592
rect 14 582 27 592
rect 42 582 72 596
rect 115 582 158 596
rect 182 593 189 600
rect 192 596 259 620
rect 291 620 463 622
rect 261 598 289 602
rect 291 598 371 620
rect 392 618 407 620
rect 261 596 371 598
rect 192 592 371 596
rect 165 582 195 592
rect 197 582 350 592
rect 358 582 388 592
rect 392 582 422 596
rect 450 582 463 620
rect 535 626 570 634
rect 535 600 536 626
rect 543 600 570 626
rect 478 582 508 596
rect 535 592 570 600
rect 572 626 613 634
rect 572 600 587 626
rect 594 600 613 626
rect 677 622 739 634
rect 751 622 826 634
rect 884 622 959 634
rect 971 622 1002 634
rect 1008 622 1043 634
rect 677 620 839 622
rect 572 592 613 600
rect 695 596 708 620
rect 723 618 738 620
rect 535 582 536 592
rect 551 582 564 592
rect 578 582 579 592
rect 594 582 607 592
rect 622 582 652 596
rect 695 582 738 596
rect 762 593 769 600
rect 772 596 839 620
rect 871 620 1043 622
rect 841 598 869 602
rect 871 598 951 620
rect 972 618 987 620
rect 841 596 951 598
rect 772 592 951 596
rect 745 582 775 592
rect 777 582 930 592
rect 938 582 968 592
rect 972 582 1002 596
rect 1030 582 1043 620
rect 1115 626 1150 634
rect 1115 600 1116 626
rect 1123 600 1150 626
rect 1058 582 1088 596
rect 1115 592 1150 600
rect 1152 626 1193 634
rect 1152 600 1167 626
rect 1174 600 1193 626
rect 1257 622 1319 634
rect 1331 622 1406 634
rect 1464 622 1539 634
rect 1551 622 1582 634
rect 1588 622 1623 634
rect 1257 620 1419 622
rect 1275 611 1288 620
rect 1303 618 1318 620
rect 1352 611 1419 620
rect 1451 620 1623 622
rect 1451 611 1531 620
rect 1552 618 1567 620
rect 1610 611 1623 620
rect 1695 626 1730 634
rect 1695 611 1696 626
rect 1703 611 1730 626
rect 1732 626 1773 634
rect 1732 611 1747 626
rect 1754 611 1773 626
rect 1152 592 1193 600
rect 1115 582 1116 592
rect 1131 582 1144 592
rect 1158 582 1159 592
rect 1174 582 1187 592
rect 1202 582 1232 596
rect -2 576 1261 582
rect -1 568 1261 576
rect 14 538 27 568
rect 42 550 72 568
rect 115 554 129 568
rect 165 554 385 568
rect 116 552 129 554
rect 82 540 97 552
rect 79 538 101 540
rect 106 538 136 552
rect 197 550 350 554
rect 179 538 371 550
rect 414 538 444 552
rect 450 538 463 568
rect 478 550 508 568
rect 551 538 564 568
rect 594 538 607 568
rect 622 550 652 568
rect 695 554 709 568
rect 745 554 965 568
rect 696 552 709 554
rect 662 540 677 552
rect 659 538 681 540
rect 686 538 716 552
rect 777 550 930 554
rect 759 538 951 550
rect 994 538 1024 552
rect 1030 538 1043 568
rect 1058 550 1088 568
rect 1131 538 1144 568
rect 1174 538 1187 568
rect 1202 550 1232 568
rect 1242 540 1257 552
rect 1239 538 1261 540
rect -1 524 1261 538
rect 14 420 27 524
rect 72 502 73 512
rect 88 502 101 512
rect 72 498 101 502
rect 106 498 136 524
rect 154 510 170 512
rect 242 510 295 524
rect 243 508 307 510
rect 350 508 365 524
rect 414 521 444 524
rect 414 518 450 521
rect 380 510 396 512
rect 154 498 169 502
rect 72 496 169 498
rect 197 496 365 508
rect 381 498 396 502
rect 414 499 453 518
rect 472 512 479 513
rect 478 505 479 512
rect 462 502 463 505
rect 478 502 491 505
rect 414 498 444 499
rect 453 498 459 499
rect 462 498 491 502
rect 381 497 491 498
rect 381 496 497 497
rect 56 488 107 496
rect 56 476 81 488
rect 88 476 107 488
rect 138 488 188 496
rect 138 480 154 488
rect 161 486 188 488
rect 197 486 418 496
rect 161 476 418 486
rect 447 488 497 496
rect 447 479 463 488
rect 56 468 107 476
rect 154 468 418 476
rect 444 476 463 479
rect 470 476 497 488
rect 444 468 497 476
rect 72 460 73 468
rect 88 460 101 468
rect 72 452 88 460
rect 69 445 88 448
rect 69 436 91 445
rect 42 426 91 436
rect 42 420 72 426
rect 91 421 96 426
rect 14 404 88 420
rect 106 412 136 468
rect 171 458 379 468
rect 414 464 459 468
rect 462 467 463 468
rect 478 467 491 468
rect 197 428 386 458
rect 212 425 386 428
rect 205 422 386 425
rect 14 402 27 404
rect 42 402 76 404
rect 14 386 88 402
rect 115 398 128 412
rect 143 398 159 414
rect 205 409 216 422
rect -2 364 -1 380
rect 14 364 27 386
rect 42 364 72 386
rect 115 382 177 398
rect 205 391 216 407
rect 221 402 231 422
rect 241 402 255 422
rect 258 409 267 422
rect 283 409 292 422
rect 221 391 255 402
rect 258 391 267 407
rect 283 391 292 407
rect 299 402 309 422
rect 319 402 333 422
rect 334 409 345 422
rect 299 391 333 402
rect 334 391 345 407
rect 391 398 407 414
rect 414 412 444 464
rect 478 460 479 467
rect 463 452 479 460
rect 450 420 463 439
rect 478 420 508 436
rect 450 404 524 420
rect 450 402 463 404
rect 478 402 512 404
rect 115 380 128 382
rect 143 380 177 382
rect 115 364 177 380
rect 221 375 237 382
rect 299 375 329 386
rect 377 382 423 398
rect 450 386 524 402
rect 377 380 411 382
rect 376 364 423 380
rect 450 364 463 386
rect 478 364 508 386
rect 535 364 536 380
rect 551 364 564 524
rect 594 420 607 524
rect 652 502 653 512
rect 668 502 681 512
rect 652 498 681 502
rect 686 498 716 524
rect 734 510 750 512
rect 822 510 875 524
rect 823 508 887 510
rect 930 508 945 524
rect 994 521 1024 524
rect 994 518 1030 521
rect 960 510 976 512
rect 734 498 749 502
rect 652 496 749 498
rect 777 496 945 508
rect 961 498 976 502
rect 994 499 1033 518
rect 1052 512 1059 513
rect 1058 505 1059 512
rect 1042 502 1043 505
rect 1058 502 1071 505
rect 994 498 1024 499
rect 1033 498 1039 499
rect 1042 498 1071 502
rect 961 497 1071 498
rect 961 496 1077 497
rect 636 488 687 496
rect 636 476 661 488
rect 668 476 687 488
rect 718 488 768 496
rect 718 480 734 488
rect 741 486 768 488
rect 777 486 998 496
rect 741 476 998 486
rect 1027 488 1077 496
rect 1027 479 1043 488
rect 636 468 687 476
rect 734 468 998 476
rect 1024 476 1043 479
rect 1050 476 1077 488
rect 1024 468 1077 476
rect 652 460 653 468
rect 668 460 681 468
rect 652 452 668 460
rect 649 445 668 448
rect 649 436 671 445
rect 622 426 671 436
rect 622 420 652 426
rect 671 421 676 426
rect 594 404 668 420
rect 686 412 716 468
rect 751 458 959 468
rect 994 464 1039 468
rect 1042 467 1043 468
rect 1058 467 1071 468
rect 777 428 966 458
rect 792 425 966 428
rect 785 422 966 425
rect 594 402 607 404
rect 622 402 656 404
rect 594 386 668 402
rect 695 398 708 412
rect 723 398 739 414
rect 785 409 796 422
rect 578 364 579 380
rect 594 364 607 386
rect 622 364 652 386
rect 695 382 757 398
rect 785 391 796 407
rect 801 402 811 422
rect 821 402 835 422
rect 838 409 847 422
rect 863 409 872 422
rect 801 391 835 402
rect 838 391 847 407
rect 863 391 872 407
rect 879 402 889 422
rect 899 402 913 422
rect 914 409 925 422
rect 879 391 913 402
rect 914 391 925 407
rect 971 398 987 414
rect 994 412 1024 464
rect 1058 460 1059 467
rect 1043 452 1059 460
rect 1030 420 1043 439
rect 1058 420 1088 436
rect 1030 404 1104 420
rect 1030 402 1043 404
rect 1058 402 1092 404
rect 695 380 708 382
rect 723 380 757 382
rect 695 364 757 380
rect 801 375 817 382
rect 879 375 909 386
rect 957 382 1003 398
rect 1030 386 1104 402
rect 957 380 991 382
rect 956 364 1003 380
rect 1030 364 1043 386
rect 1058 364 1088 386
rect 1115 364 1116 380
rect 1131 364 1144 524
rect 1174 420 1187 524
rect 1232 502 1233 512
rect 1248 502 1261 512
rect 1232 496 1261 502
rect 1216 488 1261 496
rect 1216 476 1241 488
rect 1248 476 1261 488
rect 1216 468 1261 476
rect 1232 460 1233 468
rect 1248 460 1261 468
rect 1232 452 1248 460
rect 1229 445 1248 448
rect 1229 436 1251 445
rect 1202 426 1251 436
rect 1202 420 1232 426
rect 1251 421 1256 426
rect 1174 404 1248 420
rect 1174 402 1187 404
rect 1202 402 1236 404
rect 1174 386 1248 402
rect 1158 364 1159 380
rect 1174 364 1187 386
rect 1202 364 1232 386
rect -8 356 33 364
rect -8 330 7 356
rect 14 330 33 356
rect 97 352 159 364
rect 171 352 246 364
rect 304 352 379 364
rect 391 352 422 364
rect 428 352 463 364
rect 97 350 259 352
rect -8 322 33 330
rect 115 326 128 350
rect 143 348 158 350
rect -2 312 -1 322
rect 14 312 27 322
rect 42 312 72 326
rect 115 312 158 326
rect 182 323 189 330
rect 192 326 259 350
rect 291 350 463 352
rect 261 328 289 332
rect 291 328 371 350
rect 392 348 407 350
rect 261 326 371 328
rect 192 322 371 326
rect 165 312 195 322
rect 197 312 350 322
rect 358 312 388 322
rect 392 312 422 326
rect 450 312 463 350
rect 535 356 570 364
rect 535 330 536 356
rect 543 330 570 356
rect 478 312 508 326
rect 535 322 570 330
rect 572 356 613 364
rect 572 330 587 356
rect 594 330 613 356
rect 677 352 739 364
rect 751 352 826 364
rect 884 352 959 364
rect 971 352 1002 364
rect 1008 352 1043 364
rect 677 350 839 352
rect 572 322 613 330
rect 695 326 708 350
rect 723 348 738 350
rect 535 312 536 322
rect 551 312 564 322
rect 578 312 579 322
rect 594 312 607 322
rect 622 312 652 326
rect 695 312 738 326
rect 762 323 769 330
rect 772 326 839 350
rect 871 350 1043 352
rect 841 328 869 332
rect 871 328 951 350
rect 972 348 987 350
rect 841 326 951 328
rect 772 322 951 326
rect 745 312 775 322
rect 777 312 930 322
rect 938 312 968 322
rect 972 312 1002 326
rect 1030 312 1043 350
rect 1115 356 1150 364
rect 1115 330 1116 356
rect 1123 330 1150 356
rect 1058 312 1088 326
rect 1115 322 1150 330
rect 1152 356 1193 364
rect 1152 330 1167 356
rect 1174 330 1193 356
rect 1257 350 1261 364
rect 1152 322 1193 330
rect 1115 312 1116 322
rect 1131 312 1144 322
rect 1158 312 1159 322
rect 1174 312 1187 322
rect 1202 312 1232 326
rect -2 306 1261 312
rect -1 298 1261 306
rect 14 268 27 298
rect 42 280 72 298
rect 115 284 129 298
rect 165 284 385 298
rect 116 282 129 284
rect 82 270 97 282
rect 79 268 101 270
rect 106 268 136 282
rect 197 280 350 284
rect 179 268 371 280
rect 414 268 444 282
rect 450 268 463 298
rect 478 280 508 298
rect 551 268 564 298
rect 594 268 607 298
rect 622 280 652 298
rect 695 284 709 298
rect 745 284 965 298
rect 696 282 709 284
rect 662 270 677 282
rect 659 268 681 270
rect 686 268 716 282
rect 777 280 930 284
rect 759 268 951 280
rect 994 268 1024 282
rect 1030 268 1043 298
rect 1058 280 1088 298
rect 1131 268 1144 298
rect 1174 268 1187 298
rect 1202 280 1232 298
rect 1242 270 1257 282
rect 1239 268 1261 270
rect -1 254 1261 268
rect 14 150 27 254
rect 72 232 73 242
rect 88 232 101 242
rect 72 228 101 232
rect 106 228 136 254
rect 154 240 170 242
rect 242 240 295 254
rect 243 238 307 240
rect 350 238 365 254
rect 414 251 444 254
rect 414 248 450 251
rect 380 240 396 242
rect 154 228 169 232
rect 72 226 169 228
rect 197 226 365 238
rect 381 228 396 232
rect 414 229 453 248
rect 472 242 479 243
rect 478 235 479 242
rect 462 232 463 235
rect 478 232 491 235
rect 414 228 444 229
rect 453 228 459 229
rect 462 228 491 232
rect 381 227 491 228
rect 381 226 497 227
rect 56 218 107 226
rect 56 206 81 218
rect 88 206 107 218
rect 138 218 188 226
rect 138 210 154 218
rect 161 216 188 218
rect 197 216 418 226
rect 161 206 418 216
rect 447 218 497 226
rect 447 209 463 218
rect 56 198 107 206
rect 154 198 418 206
rect 444 206 463 209
rect 470 206 497 218
rect 444 198 497 206
rect 72 190 73 198
rect 88 190 101 198
rect 72 182 88 190
rect 69 175 88 178
rect 69 166 91 175
rect 42 156 91 166
rect 42 150 72 156
rect 91 151 96 156
rect 14 134 88 150
rect 106 142 136 198
rect 171 188 379 198
rect 414 194 459 198
rect 462 197 463 198
rect 478 197 491 198
rect 197 158 386 188
rect 212 155 386 158
rect 205 152 386 155
rect 14 132 27 134
rect 42 132 76 134
rect 14 116 88 132
rect 115 128 128 142
rect 143 128 159 144
rect 205 139 216 152
rect -2 94 -1 110
rect 14 94 27 116
rect 42 94 72 116
rect 115 112 177 128
rect 205 121 216 137
rect 221 132 231 152
rect 241 132 255 152
rect 258 139 267 152
rect 283 139 292 152
rect 221 121 255 132
rect 258 121 267 137
rect 283 121 292 137
rect 299 132 309 152
rect 319 132 333 152
rect 334 139 345 152
rect 299 121 333 132
rect 334 121 345 137
rect 391 128 407 144
rect 414 142 444 194
rect 478 190 479 197
rect 463 182 479 190
rect 450 150 463 169
rect 478 150 508 166
rect 450 134 524 150
rect 450 132 463 134
rect 478 132 512 134
rect 115 110 128 112
rect 143 110 177 112
rect 115 94 177 110
rect 221 105 237 112
rect 299 105 329 116
rect 377 112 423 128
rect 450 116 524 132
rect 377 110 411 112
rect 376 94 423 110
rect 450 94 463 116
rect 478 94 508 116
rect 535 94 536 110
rect 551 94 564 254
rect 594 150 607 254
rect 652 232 653 242
rect 668 232 681 242
rect 652 228 681 232
rect 686 228 716 254
rect 734 240 750 242
rect 822 240 875 254
rect 823 238 887 240
rect 930 238 945 254
rect 994 251 1024 254
rect 994 248 1030 251
rect 960 240 976 242
rect 734 228 749 232
rect 652 226 749 228
rect 777 226 945 238
rect 961 228 976 232
rect 994 229 1033 248
rect 1052 242 1059 243
rect 1058 235 1059 242
rect 1042 232 1043 235
rect 1058 232 1071 235
rect 994 228 1024 229
rect 1033 228 1039 229
rect 1042 228 1071 232
rect 961 227 1071 228
rect 961 226 1077 227
rect 636 218 687 226
rect 636 206 661 218
rect 668 206 687 218
rect 718 218 768 226
rect 718 210 734 218
rect 741 216 768 218
rect 777 216 998 226
rect 741 206 998 216
rect 1027 218 1077 226
rect 1027 209 1043 218
rect 636 198 687 206
rect 734 198 998 206
rect 1024 206 1043 209
rect 1050 206 1077 218
rect 1024 198 1077 206
rect 652 190 653 198
rect 668 190 681 198
rect 652 182 668 190
rect 649 175 668 178
rect 649 166 671 175
rect 622 156 671 166
rect 622 150 652 156
rect 671 151 676 156
rect 594 134 668 150
rect 686 142 716 198
rect 751 188 959 198
rect 994 194 1039 198
rect 1042 197 1043 198
rect 1058 197 1071 198
rect 777 158 966 188
rect 792 155 966 158
rect 785 152 966 155
rect 594 132 607 134
rect 622 132 656 134
rect 594 116 668 132
rect 695 128 708 142
rect 723 128 739 144
rect 785 139 796 152
rect 578 94 579 110
rect 594 94 607 116
rect 622 94 652 116
rect 695 112 757 128
rect 785 121 796 137
rect 801 132 811 152
rect 821 132 835 152
rect 838 139 847 152
rect 863 139 872 152
rect 801 121 835 132
rect 838 121 847 137
rect 863 121 872 137
rect 879 132 889 152
rect 899 132 913 152
rect 914 139 925 152
rect 879 121 913 132
rect 914 121 925 137
rect 971 128 987 144
rect 994 142 1024 194
rect 1058 190 1059 197
rect 1043 182 1059 190
rect 1030 150 1043 169
rect 1058 150 1088 166
rect 1030 134 1104 150
rect 1030 132 1043 134
rect 1058 132 1092 134
rect 695 110 708 112
rect 723 110 757 112
rect 695 94 757 110
rect 801 105 817 112
rect 879 105 909 116
rect 957 112 1003 128
rect 1030 116 1104 132
rect 957 110 991 112
rect 956 94 1003 110
rect 1030 94 1043 116
rect 1058 94 1088 116
rect 1115 94 1116 110
rect 1131 94 1144 254
rect 1174 150 1187 254
rect 1232 232 1233 242
rect 1248 232 1261 242
rect 1232 226 1261 232
rect 1216 218 1261 226
rect 1216 206 1241 218
rect 1248 206 1261 218
rect 1216 198 1261 206
rect 1232 190 1233 198
rect 1248 190 1261 198
rect 1232 182 1248 190
rect 1229 175 1248 178
rect 1229 166 1251 175
rect 1202 156 1251 166
rect 1202 150 1232 156
rect 1251 151 1256 156
rect 1174 134 1248 150
rect 1174 132 1187 134
rect 1202 132 1236 134
rect 1174 116 1248 132
rect 1158 94 1159 110
rect 1174 94 1187 116
rect 1202 94 1232 116
rect -8 86 33 94
rect -8 60 7 86
rect 14 60 33 86
rect 97 82 159 94
rect 171 82 246 94
rect 304 82 379 94
rect 391 82 422 94
rect 428 82 463 94
rect 97 80 259 82
rect -8 52 33 60
rect 115 56 128 80
rect 143 78 158 80
rect -2 42 -1 52
rect 14 42 27 52
rect 42 42 72 56
rect 115 42 158 56
rect 182 53 189 60
rect 192 56 259 80
rect 291 80 463 82
rect 261 58 289 62
rect 291 58 371 80
rect 392 78 407 80
rect 261 56 371 58
rect 192 52 371 56
rect 165 42 195 52
rect 197 42 350 52
rect 358 42 388 52
rect 392 42 422 56
rect 450 42 463 80
rect 535 86 570 94
rect 535 60 536 86
rect 543 60 570 86
rect 478 42 508 56
rect 535 52 570 60
rect 572 86 613 94
rect 572 60 587 86
rect 594 60 613 86
rect 677 82 739 94
rect 751 82 826 94
rect 884 82 959 94
rect 971 82 1002 94
rect 1008 82 1043 94
rect 677 80 839 82
rect 572 52 613 60
rect 695 56 708 80
rect 723 78 738 80
rect 535 42 536 52
rect 551 42 564 52
rect 578 42 579 52
rect 594 42 607 52
rect 622 42 652 56
rect 695 42 738 56
rect 762 53 769 60
rect 772 56 839 80
rect 871 80 1043 82
rect 841 58 869 62
rect 871 58 951 80
rect 972 78 987 80
rect 841 56 951 58
rect 772 52 951 56
rect 745 42 775 52
rect 777 42 930 52
rect 938 42 968 52
rect 972 42 1002 56
rect 1030 42 1043 80
rect 1115 86 1150 94
rect 1115 60 1116 86
rect 1123 60 1150 86
rect 1058 42 1088 56
rect 1115 52 1150 60
rect 1152 86 1193 94
rect 1152 60 1167 86
rect 1174 60 1193 86
rect 1257 80 1261 94
rect 1152 52 1193 60
rect 1115 42 1116 52
rect 1131 42 1144 52
rect 1158 42 1159 52
rect 1174 42 1187 52
rect 1202 42 1232 56
rect -2 36 1261 42
rect -1 28 1261 36
rect 14 -2 27 28
rect 42 10 72 28
rect 115 14 129 28
rect 165 14 385 28
rect 116 12 129 14
rect 82 0 97 12
rect 79 -2 101 0
rect 106 -2 136 12
rect 197 10 350 14
rect 179 -2 371 10
rect 414 -2 444 12
rect 450 -2 463 28
rect 478 10 508 28
rect 551 -2 564 28
rect 594 -2 607 28
rect 622 10 652 28
rect 695 14 709 28
rect 745 14 965 28
rect 696 12 709 14
rect 662 0 677 12
rect 659 -2 681 0
rect 686 -2 716 12
rect 777 10 930 14
rect 759 -2 951 10
rect 994 -2 1024 12
rect 1030 -2 1043 28
rect 1058 10 1088 28
rect 1131 -2 1144 28
rect 1174 -2 1187 28
rect 1202 10 1232 28
rect 1242 0 1257 12
rect 1239 -2 1261 0
rect -1 -16 1261 -2
rect 14 -120 27 -16
rect 72 -38 73 -28
rect 88 -38 101 -28
rect 72 -42 101 -38
rect 106 -42 136 -16
rect 154 -30 170 -28
rect 242 -30 295 -16
rect 243 -32 307 -30
rect 350 -32 365 -16
rect 414 -19 444 -16
rect 414 -22 450 -19
rect 380 -30 396 -28
rect 154 -42 169 -38
rect 72 -44 169 -42
rect 197 -44 365 -32
rect 381 -42 396 -38
rect 414 -41 453 -22
rect 472 -28 479 -27
rect 478 -35 479 -28
rect 462 -38 463 -35
rect 478 -38 491 -35
rect 414 -42 444 -41
rect 453 -42 459 -41
rect 462 -42 491 -38
rect 381 -43 491 -42
rect 381 -44 497 -43
rect 56 -52 107 -44
rect 56 -64 81 -52
rect 88 -64 107 -52
rect 138 -52 188 -44
rect 138 -60 154 -52
rect 161 -54 188 -52
rect 197 -54 418 -44
rect 161 -64 418 -54
rect 447 -52 497 -44
rect 447 -61 463 -52
rect 56 -72 107 -64
rect 154 -72 418 -64
rect 444 -64 463 -61
rect 470 -64 497 -52
rect 444 -72 497 -64
rect 72 -80 73 -72
rect 88 -80 101 -72
rect 72 -88 88 -80
rect 69 -95 88 -92
rect 69 -104 91 -95
rect 42 -114 91 -104
rect 42 -120 72 -114
rect 91 -119 96 -114
rect 14 -136 88 -120
rect 106 -128 136 -72
rect 171 -82 379 -72
rect 414 -76 459 -72
rect 462 -73 463 -72
rect 478 -73 491 -72
rect 197 -112 386 -82
rect 212 -115 386 -112
rect 205 -118 386 -115
rect 14 -138 27 -136
rect 42 -138 76 -136
rect 14 -154 88 -138
rect 115 -142 128 -128
rect 143 -142 159 -126
rect 205 -131 216 -118
rect -2 -176 -1 -160
rect 14 -176 27 -154
rect 42 -176 72 -154
rect 115 -158 177 -142
rect 205 -149 216 -133
rect 221 -138 231 -118
rect 241 -138 255 -118
rect 258 -131 267 -118
rect 283 -131 292 -118
rect 221 -149 255 -138
rect 258 -149 267 -133
rect 283 -149 292 -133
rect 299 -138 309 -118
rect 319 -138 333 -118
rect 334 -131 345 -118
rect 299 -149 333 -138
rect 334 -149 345 -133
rect 391 -142 407 -126
rect 414 -128 444 -76
rect 478 -80 479 -73
rect 463 -88 479 -80
rect 450 -120 463 -101
rect 478 -120 508 -104
rect 450 -136 524 -120
rect 450 -138 463 -136
rect 478 -138 512 -136
rect 115 -160 128 -158
rect 143 -160 177 -158
rect 115 -176 177 -160
rect 221 -165 237 -158
rect 299 -165 329 -154
rect 377 -158 423 -142
rect 450 -154 524 -138
rect 377 -160 411 -158
rect 376 -176 423 -160
rect 450 -176 463 -154
rect 478 -176 508 -154
rect 535 -176 536 -160
rect 551 -176 564 -16
rect 594 -120 607 -16
rect 652 -38 653 -28
rect 668 -38 681 -28
rect 652 -42 681 -38
rect 686 -42 716 -16
rect 734 -30 750 -28
rect 822 -30 875 -16
rect 823 -32 887 -30
rect 930 -32 945 -16
rect 994 -19 1024 -16
rect 994 -22 1030 -19
rect 960 -30 976 -28
rect 734 -42 749 -38
rect 652 -44 749 -42
rect 777 -44 945 -32
rect 961 -42 976 -38
rect 994 -41 1033 -22
rect 1052 -28 1059 -27
rect 1058 -35 1059 -28
rect 1042 -38 1043 -35
rect 1058 -38 1071 -35
rect 994 -42 1024 -41
rect 1033 -42 1039 -41
rect 1042 -42 1071 -38
rect 961 -43 1071 -42
rect 961 -44 1077 -43
rect 636 -52 687 -44
rect 636 -64 661 -52
rect 668 -64 687 -52
rect 718 -52 768 -44
rect 718 -60 734 -52
rect 741 -54 768 -52
rect 777 -54 998 -44
rect 741 -64 998 -54
rect 1027 -52 1077 -44
rect 1027 -61 1043 -52
rect 636 -72 687 -64
rect 734 -72 998 -64
rect 1024 -64 1043 -61
rect 1050 -64 1077 -52
rect 1024 -72 1077 -64
rect 652 -80 653 -72
rect 668 -80 681 -72
rect 652 -88 668 -80
rect 649 -95 668 -92
rect 649 -104 671 -95
rect 622 -114 671 -104
rect 622 -120 652 -114
rect 671 -119 676 -114
rect 594 -136 668 -120
rect 686 -128 716 -72
rect 751 -82 959 -72
rect 994 -76 1039 -72
rect 1042 -73 1043 -72
rect 1058 -73 1071 -72
rect 777 -112 966 -82
rect 792 -115 966 -112
rect 785 -118 966 -115
rect 594 -138 607 -136
rect 622 -138 656 -136
rect 594 -154 668 -138
rect 695 -142 708 -128
rect 723 -142 739 -126
rect 785 -131 796 -118
rect 578 -176 579 -160
rect 594 -176 607 -154
rect 622 -176 652 -154
rect 695 -158 757 -142
rect 785 -149 796 -133
rect 801 -138 811 -118
rect 821 -138 835 -118
rect 838 -131 847 -118
rect 863 -131 872 -118
rect 801 -149 835 -138
rect 838 -149 847 -133
rect 863 -149 872 -133
rect 879 -138 889 -118
rect 899 -138 913 -118
rect 914 -131 925 -118
rect 879 -149 913 -138
rect 914 -149 925 -133
rect 971 -142 987 -126
rect 994 -128 1024 -76
rect 1058 -80 1059 -73
rect 1043 -88 1059 -80
rect 1030 -120 1043 -101
rect 1058 -120 1088 -104
rect 1030 -136 1104 -120
rect 1030 -138 1043 -136
rect 1058 -138 1092 -136
rect 695 -160 708 -158
rect 723 -160 757 -158
rect 695 -176 757 -160
rect 801 -165 817 -158
rect 879 -165 909 -154
rect 957 -158 1003 -142
rect 1030 -154 1104 -138
rect 957 -160 991 -158
rect 956 -176 1003 -160
rect 1030 -176 1043 -154
rect 1058 -176 1088 -154
rect 1115 -176 1116 -160
rect 1131 -176 1144 -16
rect 1174 -120 1187 -16
rect 1232 -38 1233 -28
rect 1248 -38 1261 -28
rect 1232 -44 1261 -38
rect 1216 -52 1261 -44
rect 1216 -64 1241 -52
rect 1248 -64 1261 -52
rect 1216 -72 1261 -64
rect 1232 -80 1233 -72
rect 1248 -80 1261 -72
rect 1232 -88 1248 -80
rect 1229 -95 1248 -92
rect 1229 -104 1251 -95
rect 1202 -114 1251 -104
rect 1202 -120 1232 -114
rect 1251 -119 1256 -114
rect 1174 -136 1248 -120
rect 1174 -138 1187 -136
rect 1202 -138 1236 -136
rect 1174 -154 1248 -138
rect 1158 -176 1159 -160
rect 1174 -176 1187 -154
rect 1202 -176 1232 -154
rect -8 -184 33 -176
rect -8 -210 7 -184
rect 14 -210 33 -184
rect 97 -188 159 -176
rect 171 -188 246 -176
rect 304 -188 379 -176
rect 391 -188 422 -176
rect 428 -188 463 -176
rect 97 -190 259 -188
rect -8 -218 33 -210
rect 115 -214 128 -190
rect 143 -192 158 -190
rect -2 -228 -1 -218
rect 14 -228 27 -218
rect 42 -228 72 -214
rect 115 -228 158 -214
rect 182 -217 189 -210
rect 192 -214 259 -190
rect 291 -190 463 -188
rect 261 -212 289 -208
rect 291 -212 371 -190
rect 392 -192 407 -190
rect 261 -214 371 -212
rect 192 -218 371 -214
rect 165 -228 195 -218
rect 197 -228 350 -218
rect 358 -228 388 -218
rect 392 -228 422 -214
rect 450 -228 463 -190
rect 535 -184 570 -176
rect 535 -210 536 -184
rect 543 -210 570 -184
rect 478 -228 508 -214
rect 535 -218 570 -210
rect 572 -184 613 -176
rect 572 -210 587 -184
rect 594 -210 613 -184
rect 677 -188 739 -176
rect 751 -188 826 -176
rect 884 -188 959 -176
rect 971 -188 1002 -176
rect 1008 -188 1043 -176
rect 677 -190 839 -188
rect 572 -218 613 -210
rect 695 -214 708 -190
rect 723 -192 738 -190
rect 535 -228 536 -218
rect 551 -228 564 -218
rect 578 -228 579 -218
rect 594 -228 607 -218
rect 622 -228 652 -214
rect 695 -228 738 -214
rect 762 -217 769 -210
rect 772 -214 839 -190
rect 871 -190 1043 -188
rect 841 -212 869 -208
rect 871 -212 951 -190
rect 972 -192 987 -190
rect 841 -214 951 -212
rect 772 -218 951 -214
rect 745 -228 775 -218
rect 777 -228 930 -218
rect 938 -228 968 -218
rect 972 -228 1002 -214
rect 1030 -228 1043 -190
rect 1115 -184 1150 -176
rect 1115 -210 1116 -184
rect 1123 -210 1150 -184
rect 1058 -228 1088 -214
rect 1115 -218 1150 -210
rect 1152 -184 1193 -176
rect 1152 -210 1167 -184
rect 1174 -210 1193 -184
rect 1257 -190 1261 -176
rect 1152 -218 1193 -210
rect 1115 -228 1116 -218
rect 1131 -228 1144 -218
rect 1158 -228 1159 -218
rect 1174 -228 1187 -218
rect 1202 -228 1232 -214
rect -2 -234 1261 -228
rect -1 -242 1261 -234
rect 14 -272 27 -242
rect 42 -260 72 -242
rect 115 -256 129 -242
rect 165 -256 385 -242
rect 116 -258 129 -256
rect 82 -270 97 -258
rect 79 -272 101 -270
rect 106 -272 136 -258
rect 197 -260 350 -256
rect 179 -272 371 -260
rect 414 -272 444 -258
rect 450 -272 463 -242
rect 478 -260 508 -242
rect 551 -272 564 -242
rect 594 -272 607 -242
rect 622 -260 652 -242
rect 695 -256 709 -242
rect 745 -256 965 -242
rect 696 -258 709 -256
rect 662 -270 677 -258
rect 659 -272 681 -270
rect 686 -272 716 -258
rect 777 -260 930 -256
rect 759 -272 951 -260
rect 994 -272 1024 -258
rect 1030 -272 1043 -242
rect 1058 -260 1088 -242
rect 1131 -272 1144 -242
rect 1174 -272 1187 -242
rect 1202 -260 1232 -242
rect 1242 -270 1257 -258
rect 1239 -272 1261 -270
rect -1 -286 1261 -272
rect 14 -390 27 -286
rect 72 -308 73 -298
rect 88 -308 101 -298
rect 72 -312 101 -308
rect 106 -312 136 -286
rect 154 -300 170 -298
rect 242 -300 295 -286
rect 243 -302 307 -300
rect 350 -302 365 -286
rect 414 -289 444 -286
rect 414 -292 450 -289
rect 380 -300 396 -298
rect 154 -312 169 -308
rect 72 -314 169 -312
rect 197 -314 365 -302
rect 381 -312 396 -308
rect 414 -311 453 -292
rect 472 -298 479 -297
rect 478 -305 479 -298
rect 462 -308 463 -305
rect 478 -308 491 -305
rect 414 -312 444 -311
rect 453 -312 459 -311
rect 462 -312 491 -308
rect 381 -313 491 -312
rect 381 -314 497 -313
rect 56 -322 107 -314
rect 56 -334 81 -322
rect 88 -334 107 -322
rect 138 -322 188 -314
rect 138 -330 154 -322
rect 161 -324 188 -322
rect 197 -324 418 -314
rect 161 -334 418 -324
rect 447 -322 497 -314
rect 447 -331 463 -322
rect 56 -342 107 -334
rect 154 -342 418 -334
rect 444 -334 463 -331
rect 470 -334 497 -322
rect 444 -342 497 -334
rect 72 -350 73 -342
rect 88 -350 101 -342
rect 72 -358 88 -350
rect 69 -365 88 -362
rect 69 -374 91 -365
rect 42 -384 91 -374
rect 42 -390 72 -384
rect 91 -389 96 -384
rect 14 -406 88 -390
rect 106 -398 136 -342
rect 171 -352 379 -342
rect 414 -346 459 -342
rect 462 -343 463 -342
rect 478 -343 491 -342
rect 197 -382 386 -352
rect 212 -385 386 -382
rect 205 -388 386 -385
rect 14 -408 27 -406
rect 42 -408 76 -406
rect 14 -424 88 -408
rect 115 -412 128 -398
rect 143 -412 159 -396
rect 205 -401 216 -388
rect -2 -446 -1 -430
rect 14 -446 27 -424
rect 42 -446 72 -424
rect 115 -428 177 -412
rect 205 -419 216 -403
rect 221 -408 231 -388
rect 241 -408 255 -388
rect 258 -401 267 -388
rect 283 -401 292 -388
rect 221 -419 255 -408
rect 258 -419 267 -403
rect 283 -419 292 -403
rect 299 -408 309 -388
rect 319 -408 333 -388
rect 334 -401 345 -388
rect 299 -419 333 -408
rect 334 -419 345 -403
rect 391 -412 407 -396
rect 414 -398 444 -346
rect 478 -350 479 -343
rect 463 -358 479 -350
rect 450 -390 463 -371
rect 478 -390 508 -374
rect 450 -406 524 -390
rect 450 -408 463 -406
rect 478 -408 512 -406
rect 115 -430 128 -428
rect 143 -430 177 -428
rect 115 -446 177 -430
rect 221 -435 237 -428
rect 299 -435 329 -424
rect 377 -428 423 -412
rect 450 -424 524 -408
rect 377 -430 411 -428
rect 376 -446 423 -430
rect 450 -446 463 -424
rect 478 -446 508 -424
rect 535 -446 536 -430
rect 551 -446 564 -286
rect 594 -390 607 -286
rect 652 -308 653 -298
rect 668 -308 681 -298
rect 652 -312 681 -308
rect 686 -312 716 -286
rect 734 -300 750 -298
rect 822 -300 875 -286
rect 823 -302 887 -300
rect 930 -302 945 -286
rect 994 -289 1024 -286
rect 994 -292 1030 -289
rect 960 -300 976 -298
rect 734 -312 749 -308
rect 652 -314 749 -312
rect 777 -314 945 -302
rect 961 -312 976 -308
rect 994 -311 1033 -292
rect 1052 -298 1059 -297
rect 1058 -305 1059 -298
rect 1042 -308 1043 -305
rect 1058 -308 1071 -305
rect 994 -312 1024 -311
rect 1033 -312 1039 -311
rect 1042 -312 1071 -308
rect 961 -313 1071 -312
rect 961 -314 1077 -313
rect 636 -322 687 -314
rect 636 -334 661 -322
rect 668 -334 687 -322
rect 718 -322 768 -314
rect 718 -330 734 -322
rect 741 -324 768 -322
rect 777 -324 998 -314
rect 741 -334 998 -324
rect 1027 -322 1077 -314
rect 1027 -331 1043 -322
rect 636 -342 687 -334
rect 734 -342 998 -334
rect 1024 -334 1043 -331
rect 1050 -334 1077 -322
rect 1024 -342 1077 -334
rect 652 -350 653 -342
rect 668 -350 681 -342
rect 652 -358 668 -350
rect 649 -365 668 -362
rect 649 -374 671 -365
rect 622 -384 671 -374
rect 622 -390 652 -384
rect 671 -389 676 -384
rect 594 -406 668 -390
rect 686 -398 716 -342
rect 751 -352 959 -342
rect 994 -346 1039 -342
rect 1042 -343 1043 -342
rect 1058 -343 1071 -342
rect 777 -382 966 -352
rect 792 -385 966 -382
rect 785 -388 966 -385
rect 594 -408 607 -406
rect 622 -408 656 -406
rect 594 -424 668 -408
rect 695 -412 708 -398
rect 723 -412 739 -396
rect 785 -401 796 -388
rect 578 -446 579 -430
rect 594 -446 607 -424
rect 622 -446 652 -424
rect 695 -428 757 -412
rect 785 -419 796 -403
rect 801 -408 811 -388
rect 821 -408 835 -388
rect 838 -401 847 -388
rect 863 -401 872 -388
rect 801 -419 835 -408
rect 838 -419 847 -403
rect 863 -419 872 -403
rect 879 -408 889 -388
rect 899 -408 913 -388
rect 914 -401 925 -388
rect 879 -419 913 -408
rect 914 -419 925 -403
rect 971 -412 987 -396
rect 994 -398 1024 -346
rect 1058 -350 1059 -343
rect 1043 -358 1059 -350
rect 1030 -390 1043 -371
rect 1058 -390 1088 -374
rect 1030 -406 1104 -390
rect 1030 -408 1043 -406
rect 1058 -408 1092 -406
rect 695 -430 708 -428
rect 723 -430 757 -428
rect 695 -446 757 -430
rect 801 -435 817 -428
rect 879 -435 909 -424
rect 957 -428 1003 -412
rect 1030 -424 1104 -408
rect 957 -430 991 -428
rect 956 -446 1003 -430
rect 1030 -446 1043 -424
rect 1058 -446 1088 -424
rect 1115 -446 1116 -430
rect 1131 -446 1144 -286
rect 1174 -390 1187 -286
rect 1232 -308 1233 -298
rect 1248 -308 1261 -298
rect 1232 -314 1261 -308
rect 1216 -322 1261 -314
rect 1216 -334 1241 -322
rect 1248 -334 1261 -322
rect 1216 -342 1261 -334
rect 1232 -350 1233 -342
rect 1248 -350 1261 -342
rect 1232 -358 1248 -350
rect 1229 -365 1248 -362
rect 1229 -374 1251 -365
rect 1202 -384 1251 -374
rect 1202 -390 1232 -384
rect 1251 -389 1256 -384
rect 1174 -406 1248 -390
rect 1174 -408 1187 -406
rect 1202 -408 1236 -406
rect 1174 -424 1248 -408
rect 1158 -446 1159 -430
rect 1174 -446 1187 -424
rect 1202 -446 1232 -424
rect -8 -454 33 -446
rect -8 -480 7 -454
rect 14 -480 33 -454
rect 97 -458 159 -446
rect 171 -458 246 -446
rect 304 -458 379 -446
rect 391 -458 422 -446
rect 428 -458 463 -446
rect 97 -460 259 -458
rect -8 -488 33 -480
rect 115 -484 128 -460
rect 143 -462 158 -460
rect -2 -498 -1 -488
rect 14 -498 27 -488
rect 42 -498 72 -484
rect 115 -498 158 -484
rect 182 -487 189 -480
rect 192 -484 259 -460
rect 291 -460 463 -458
rect 261 -482 289 -478
rect 291 -482 371 -460
rect 392 -462 407 -460
rect 261 -484 371 -482
rect 192 -488 371 -484
rect 165 -498 195 -488
rect 197 -498 350 -488
rect 358 -498 388 -488
rect 392 -498 422 -484
rect 450 -498 463 -460
rect 535 -454 570 -446
rect 535 -480 536 -454
rect 543 -480 570 -454
rect 478 -498 508 -484
rect 535 -488 570 -480
rect 572 -454 613 -446
rect 572 -480 587 -454
rect 594 -480 613 -454
rect 677 -458 739 -446
rect 751 -458 826 -446
rect 884 -458 959 -446
rect 971 -458 1002 -446
rect 1008 -458 1043 -446
rect 677 -460 839 -458
rect 572 -488 613 -480
rect 695 -484 708 -460
rect 723 -462 738 -460
rect 535 -498 536 -488
rect 551 -498 564 -488
rect 578 -498 579 -488
rect 594 -498 607 -488
rect 622 -498 652 -484
rect 695 -498 738 -484
rect 762 -487 769 -480
rect 772 -484 839 -460
rect 871 -460 1043 -458
rect 841 -482 869 -478
rect 871 -482 951 -460
rect 972 -462 987 -460
rect 841 -484 951 -482
rect 772 -488 951 -484
rect 745 -498 775 -488
rect 777 -498 930 -488
rect 938 -498 968 -488
rect 972 -498 1002 -484
rect 1030 -498 1043 -460
rect 1115 -454 1150 -446
rect 1115 -480 1116 -454
rect 1123 -480 1150 -454
rect 1058 -498 1088 -484
rect 1115 -488 1150 -480
rect 1152 -454 1193 -446
rect 1152 -480 1167 -454
rect 1174 -480 1193 -454
rect 1257 -460 1261 -446
rect 1152 -488 1193 -480
rect 1115 -498 1116 -488
rect 1131 -498 1144 -488
rect 1158 -498 1159 -488
rect 1174 -498 1187 -488
rect 1202 -498 1232 -484
rect -2 -504 1261 -498
rect -1 -512 1261 -504
rect 14 -542 27 -512
rect 42 -530 72 -512
rect 115 -526 129 -512
rect 165 -526 385 -512
rect 116 -528 129 -526
rect 82 -540 97 -528
rect 79 -542 101 -540
rect 106 -542 136 -528
rect 197 -530 350 -526
rect 179 -542 371 -530
rect 414 -542 444 -528
rect 450 -542 463 -512
rect 478 -530 508 -512
rect 551 -542 564 -512
rect 594 -542 607 -512
rect 622 -530 652 -512
rect 695 -526 709 -512
rect 745 -526 965 -512
rect 696 -528 709 -526
rect 662 -540 677 -528
rect 659 -542 681 -540
rect 686 -542 716 -528
rect 777 -530 930 -526
rect 759 -542 951 -530
rect 994 -542 1024 -528
rect 1030 -542 1043 -512
rect 1058 -530 1088 -512
rect 1131 -542 1144 -512
rect 1174 -542 1187 -512
rect 1202 -530 1232 -512
rect 1242 -540 1257 -528
rect 1239 -542 1261 -540
rect -1 -556 1261 -542
rect 14 -660 27 -556
rect 72 -578 73 -568
rect 88 -578 101 -568
rect 72 -582 101 -578
rect 106 -582 136 -556
rect 154 -570 170 -568
rect 242 -570 295 -556
rect 243 -572 307 -570
rect 350 -572 365 -556
rect 414 -559 444 -556
rect 414 -562 450 -559
rect 380 -570 396 -568
rect 154 -582 169 -578
rect 72 -584 169 -582
rect 197 -584 365 -572
rect 381 -582 396 -578
rect 414 -581 453 -562
rect 472 -568 479 -567
rect 478 -575 479 -568
rect 462 -578 463 -575
rect 478 -578 491 -575
rect 414 -582 444 -581
rect 453 -582 459 -581
rect 462 -582 491 -578
rect 381 -583 491 -582
rect 381 -584 497 -583
rect 56 -592 107 -584
rect 56 -604 81 -592
rect 88 -604 107 -592
rect 138 -592 188 -584
rect 138 -600 154 -592
rect 161 -594 188 -592
rect 197 -594 418 -584
rect 161 -604 418 -594
rect 447 -592 497 -584
rect 447 -601 463 -592
rect 56 -612 107 -604
rect 154 -612 418 -604
rect 444 -604 463 -601
rect 470 -604 497 -592
rect 444 -612 497 -604
rect 72 -620 73 -612
rect 88 -620 101 -612
rect 72 -628 88 -620
rect 69 -635 88 -632
rect 69 -644 91 -635
rect 42 -654 91 -644
rect 42 -660 72 -654
rect 91 -659 96 -654
rect 14 -676 88 -660
rect 106 -668 136 -612
rect 171 -622 379 -612
rect 414 -616 459 -612
rect 462 -613 463 -612
rect 478 -613 491 -612
rect 197 -652 386 -622
rect 212 -655 386 -652
rect 205 -658 386 -655
rect 14 -678 27 -676
rect 42 -678 76 -676
rect 14 -694 88 -678
rect 115 -682 128 -668
rect 143 -682 159 -666
rect 205 -671 216 -658
rect -2 -716 -1 -700
rect 14 -716 27 -694
rect 42 -716 72 -694
rect 115 -698 177 -682
rect 205 -689 216 -673
rect 221 -678 231 -658
rect 241 -678 255 -658
rect 258 -671 267 -658
rect 283 -671 292 -658
rect 221 -689 255 -678
rect 258 -689 267 -673
rect 283 -689 292 -673
rect 299 -678 309 -658
rect 319 -678 333 -658
rect 334 -671 345 -658
rect 299 -689 333 -678
rect 334 -689 345 -673
rect 391 -682 407 -666
rect 414 -668 444 -616
rect 478 -620 479 -613
rect 463 -628 479 -620
rect 450 -660 463 -641
rect 478 -660 508 -644
rect 450 -676 524 -660
rect 450 -678 463 -676
rect 478 -678 512 -676
rect 115 -700 128 -698
rect 143 -700 177 -698
rect 115 -716 177 -700
rect 221 -705 237 -698
rect 299 -705 329 -694
rect 377 -698 423 -682
rect 450 -694 524 -678
rect 377 -700 411 -698
rect 376 -716 423 -700
rect 450 -716 463 -694
rect 478 -716 508 -694
rect 535 -716 536 -700
rect 551 -716 564 -556
rect 594 -660 607 -556
rect 652 -578 653 -568
rect 668 -578 681 -568
rect 652 -582 681 -578
rect 686 -582 716 -556
rect 734 -570 750 -568
rect 822 -570 875 -556
rect 823 -572 887 -570
rect 930 -572 945 -556
rect 994 -559 1024 -556
rect 994 -562 1030 -559
rect 960 -570 976 -568
rect 734 -582 749 -578
rect 652 -584 749 -582
rect 777 -584 945 -572
rect 961 -582 976 -578
rect 994 -581 1033 -562
rect 1052 -568 1059 -567
rect 1058 -575 1059 -568
rect 1042 -578 1043 -575
rect 1058 -578 1071 -575
rect 994 -582 1024 -581
rect 1033 -582 1039 -581
rect 1042 -582 1071 -578
rect 961 -583 1071 -582
rect 961 -584 1077 -583
rect 636 -592 687 -584
rect 636 -604 661 -592
rect 668 -604 687 -592
rect 718 -592 768 -584
rect 718 -600 734 -592
rect 741 -594 768 -592
rect 777 -594 998 -584
rect 741 -604 998 -594
rect 1027 -592 1077 -584
rect 1027 -601 1043 -592
rect 636 -612 687 -604
rect 734 -612 998 -604
rect 1024 -604 1043 -601
rect 1050 -604 1077 -592
rect 1024 -612 1077 -604
rect 652 -620 653 -612
rect 668 -620 681 -612
rect 652 -628 668 -620
rect 649 -635 668 -632
rect 649 -644 671 -635
rect 622 -654 671 -644
rect 622 -660 652 -654
rect 671 -659 676 -654
rect 594 -676 668 -660
rect 686 -668 716 -612
rect 751 -622 959 -612
rect 994 -616 1039 -612
rect 1042 -613 1043 -612
rect 1058 -613 1071 -612
rect 777 -652 966 -622
rect 792 -655 966 -652
rect 785 -658 966 -655
rect 594 -678 607 -676
rect 622 -678 656 -676
rect 594 -694 668 -678
rect 695 -682 708 -668
rect 723 -682 739 -666
rect 785 -671 796 -658
rect 578 -716 579 -700
rect 594 -716 607 -694
rect 622 -716 652 -694
rect 695 -698 757 -682
rect 785 -689 796 -673
rect 801 -678 811 -658
rect 821 -678 835 -658
rect 838 -671 847 -658
rect 863 -671 872 -658
rect 801 -689 835 -678
rect 838 -689 847 -673
rect 863 -689 872 -673
rect 879 -678 889 -658
rect 899 -678 913 -658
rect 914 -671 925 -658
rect 879 -689 913 -678
rect 914 -689 925 -673
rect 971 -682 987 -666
rect 994 -668 1024 -616
rect 1058 -620 1059 -613
rect 1043 -628 1059 -620
rect 1030 -660 1043 -641
rect 1058 -660 1088 -644
rect 1030 -676 1104 -660
rect 1030 -678 1043 -676
rect 1058 -678 1092 -676
rect 695 -700 708 -698
rect 723 -700 757 -698
rect 695 -716 757 -700
rect 801 -705 817 -698
rect 879 -705 909 -694
rect 957 -698 1003 -682
rect 1030 -694 1104 -678
rect 957 -700 991 -698
rect 956 -716 1003 -700
rect 1030 -716 1043 -694
rect 1058 -716 1088 -694
rect 1115 -716 1116 -700
rect 1131 -716 1144 -556
rect 1174 -660 1187 -556
rect 1232 -578 1233 -568
rect 1248 -578 1261 -568
rect 1232 -584 1261 -578
rect 1216 -592 1261 -584
rect 1216 -604 1241 -592
rect 1248 -604 1261 -592
rect 1216 -612 1261 -604
rect 1232 -620 1233 -612
rect 1248 -620 1261 -612
rect 1232 -628 1248 -620
rect 1229 -635 1248 -632
rect 1229 -644 1251 -635
rect 1202 -654 1251 -644
rect 1202 -660 1232 -654
rect 1251 -659 1256 -654
rect 1174 -676 1248 -660
rect 1174 -678 1187 -676
rect 1202 -678 1236 -676
rect 1174 -694 1248 -678
rect 1158 -716 1159 -700
rect 1174 -716 1187 -694
rect 1202 -716 1232 -694
rect -8 -724 33 -716
rect -8 -750 7 -724
rect 14 -750 33 -724
rect 97 -728 159 -716
rect 171 -728 246 -716
rect 304 -728 379 -716
rect 391 -728 422 -716
rect 428 -728 463 -716
rect 97 -730 259 -728
rect -8 -758 33 -750
rect 115 -754 128 -730
rect 143 -732 158 -730
rect -2 -768 -1 -758
rect 14 -768 27 -758
rect 42 -768 72 -754
rect 115 -768 158 -754
rect 182 -757 189 -750
rect 192 -754 259 -730
rect 291 -730 463 -728
rect 261 -752 289 -748
rect 291 -752 371 -730
rect 392 -732 407 -730
rect 261 -754 371 -752
rect 192 -758 371 -754
rect 165 -768 195 -758
rect 197 -768 350 -758
rect 358 -768 388 -758
rect 392 -768 422 -754
rect 450 -768 463 -730
rect 535 -724 570 -716
rect 535 -750 536 -724
rect 543 -750 570 -724
rect 478 -768 508 -754
rect 535 -758 570 -750
rect 572 -724 613 -716
rect 572 -750 587 -724
rect 594 -750 613 -724
rect 677 -728 739 -716
rect 751 -728 826 -716
rect 884 -728 959 -716
rect 971 -728 1002 -716
rect 1008 -728 1043 -716
rect 677 -730 839 -728
rect 572 -758 613 -750
rect 695 -754 708 -730
rect 723 -732 738 -730
rect 535 -768 536 -758
rect 551 -768 564 -758
rect 578 -768 579 -758
rect 594 -768 607 -758
rect 622 -768 652 -754
rect 695 -768 738 -754
rect 762 -757 769 -750
rect 772 -754 839 -730
rect 871 -730 1043 -728
rect 841 -752 869 -748
rect 871 -752 951 -730
rect 972 -732 987 -730
rect 841 -754 951 -752
rect 772 -758 951 -754
rect 745 -768 775 -758
rect 777 -768 930 -758
rect 938 -768 968 -758
rect 972 -768 1002 -754
rect 1030 -768 1043 -730
rect 1115 -724 1150 -716
rect 1115 -750 1116 -724
rect 1123 -750 1150 -724
rect 1058 -768 1088 -754
rect 1115 -758 1150 -750
rect 1152 -724 1193 -716
rect 1152 -750 1167 -724
rect 1174 -750 1193 -724
rect 1257 -730 1261 -716
rect 1152 -758 1193 -750
rect 1115 -768 1116 -758
rect 1131 -768 1144 -758
rect 1158 -768 1159 -758
rect 1174 -768 1187 -758
rect 1202 -768 1232 -754
rect -2 -774 1261 -768
rect -1 -782 1261 -774
rect 14 -812 27 -782
rect 42 -800 72 -782
rect 115 -796 129 -782
rect 165 -796 385 -782
rect 116 -798 129 -796
rect 82 -810 97 -798
rect 79 -812 101 -810
rect 106 -812 136 -798
rect 197 -800 350 -796
rect 179 -812 371 -800
rect 414 -812 444 -798
rect 450 -812 463 -782
rect 478 -800 508 -782
rect 551 -812 564 -782
rect 594 -812 607 -782
rect 622 -800 652 -782
rect 695 -796 709 -782
rect 745 -796 965 -782
rect 696 -798 709 -796
rect 662 -810 677 -798
rect 659 -812 681 -810
rect 686 -812 716 -798
rect 777 -800 930 -796
rect 759 -812 951 -800
rect 994 -812 1024 -798
rect 1030 -812 1043 -782
rect 1058 -800 1088 -782
rect 1131 -812 1144 -782
rect 1174 -812 1187 -782
rect 1202 -800 1232 -782
rect 1242 -810 1257 -798
rect 1239 -812 1261 -810
rect -1 -826 1261 -812
rect 14 -930 27 -826
rect 72 -848 73 -838
rect 88 -848 101 -838
rect 72 -852 101 -848
rect 106 -852 136 -826
rect 154 -840 170 -838
rect 242 -840 295 -826
rect 243 -842 307 -840
rect 350 -842 365 -826
rect 414 -829 444 -826
rect 414 -832 450 -829
rect 380 -840 396 -838
rect 154 -852 169 -848
rect 72 -854 169 -852
rect 197 -854 365 -842
rect 381 -852 396 -848
rect 414 -851 453 -832
rect 472 -838 479 -837
rect 478 -845 479 -838
rect 462 -848 463 -845
rect 478 -848 491 -845
rect 414 -852 444 -851
rect 453 -852 459 -851
rect 462 -852 491 -848
rect 381 -853 491 -852
rect 381 -854 497 -853
rect 56 -862 107 -854
rect 56 -874 81 -862
rect 88 -874 107 -862
rect 138 -862 188 -854
rect 138 -870 154 -862
rect 161 -864 188 -862
rect 197 -864 418 -854
rect 161 -874 418 -864
rect 447 -862 497 -854
rect 447 -871 463 -862
rect 56 -882 107 -874
rect 154 -882 418 -874
rect 444 -874 463 -871
rect 470 -874 497 -862
rect 444 -882 497 -874
rect 72 -890 73 -882
rect 88 -890 101 -882
rect 72 -898 88 -890
rect 69 -905 88 -902
rect 69 -914 91 -905
rect 42 -924 91 -914
rect 42 -930 72 -924
rect 91 -929 96 -924
rect 14 -946 88 -930
rect 106 -938 136 -882
rect 171 -892 379 -882
rect 414 -886 459 -882
rect 462 -883 463 -882
rect 478 -883 491 -882
rect 197 -922 386 -892
rect 212 -925 386 -922
rect 205 -928 386 -925
rect 14 -948 27 -946
rect 42 -948 76 -946
rect 14 -964 88 -948
rect 115 -952 128 -938
rect 143 -952 159 -936
rect 205 -941 216 -928
rect -2 -986 -1 -970
rect 14 -986 27 -964
rect 42 -986 72 -964
rect 115 -968 177 -952
rect 205 -959 216 -943
rect 221 -948 231 -928
rect 241 -948 255 -928
rect 258 -941 267 -928
rect 283 -941 292 -928
rect 221 -959 255 -948
rect 258 -959 267 -943
rect 283 -959 292 -943
rect 299 -948 309 -928
rect 319 -948 333 -928
rect 334 -941 345 -928
rect 299 -959 333 -948
rect 334 -959 345 -943
rect 391 -952 407 -936
rect 414 -938 444 -886
rect 478 -890 479 -883
rect 463 -898 479 -890
rect 450 -930 463 -911
rect 478 -930 508 -914
rect 450 -946 524 -930
rect 450 -948 463 -946
rect 478 -948 512 -946
rect 115 -970 128 -968
rect 143 -970 177 -968
rect 115 -986 177 -970
rect 221 -975 237 -968
rect 299 -975 329 -964
rect 377 -968 423 -952
rect 450 -964 524 -948
rect 377 -970 411 -968
rect 376 -986 423 -970
rect 450 -986 463 -964
rect 478 -986 508 -964
rect 535 -986 536 -970
rect 551 -986 564 -826
rect 594 -930 607 -826
rect 652 -848 653 -838
rect 668 -848 681 -838
rect 652 -852 681 -848
rect 686 -852 716 -826
rect 734 -840 750 -838
rect 822 -840 875 -826
rect 823 -842 887 -840
rect 930 -842 945 -826
rect 994 -829 1024 -826
rect 994 -832 1030 -829
rect 960 -840 976 -838
rect 734 -852 749 -848
rect 652 -854 749 -852
rect 777 -854 945 -842
rect 961 -852 976 -848
rect 994 -851 1033 -832
rect 1052 -838 1059 -837
rect 1058 -845 1059 -838
rect 1042 -848 1043 -845
rect 1058 -848 1071 -845
rect 994 -852 1024 -851
rect 1033 -852 1039 -851
rect 1042 -852 1071 -848
rect 961 -853 1071 -852
rect 961 -854 1077 -853
rect 636 -862 687 -854
rect 636 -874 661 -862
rect 668 -874 687 -862
rect 718 -862 768 -854
rect 718 -870 734 -862
rect 741 -864 768 -862
rect 777 -864 998 -854
rect 741 -874 998 -864
rect 1027 -862 1077 -854
rect 1027 -871 1043 -862
rect 636 -882 687 -874
rect 734 -882 998 -874
rect 1024 -874 1043 -871
rect 1050 -874 1077 -862
rect 1024 -882 1077 -874
rect 652 -890 653 -882
rect 668 -890 681 -882
rect 652 -898 668 -890
rect 649 -905 668 -902
rect 649 -914 671 -905
rect 622 -924 671 -914
rect 622 -930 652 -924
rect 671 -929 676 -924
rect 594 -946 668 -930
rect 686 -938 716 -882
rect 751 -892 959 -882
rect 994 -886 1039 -882
rect 1042 -883 1043 -882
rect 1058 -883 1071 -882
rect 777 -922 966 -892
rect 792 -925 966 -922
rect 785 -928 966 -925
rect 594 -948 607 -946
rect 622 -948 656 -946
rect 594 -964 668 -948
rect 695 -952 708 -938
rect 723 -952 739 -936
rect 785 -941 796 -928
rect 578 -986 579 -970
rect 594 -986 607 -964
rect 622 -986 652 -964
rect 695 -968 757 -952
rect 785 -959 796 -943
rect 801 -948 811 -928
rect 821 -948 835 -928
rect 838 -941 847 -928
rect 863 -941 872 -928
rect 801 -959 835 -948
rect 838 -959 847 -943
rect 863 -959 872 -943
rect 879 -948 889 -928
rect 899 -948 913 -928
rect 914 -941 925 -928
rect 879 -959 913 -948
rect 914 -959 925 -943
rect 971 -952 987 -936
rect 994 -938 1024 -886
rect 1058 -890 1059 -883
rect 1043 -898 1059 -890
rect 1030 -930 1043 -911
rect 1058 -930 1088 -914
rect 1030 -946 1104 -930
rect 1030 -948 1043 -946
rect 1058 -948 1092 -946
rect 695 -970 708 -968
rect 723 -970 757 -968
rect 695 -986 757 -970
rect 801 -975 817 -968
rect 879 -975 909 -964
rect 957 -968 1003 -952
rect 1030 -964 1104 -948
rect 957 -970 991 -968
rect 956 -986 1003 -970
rect 1030 -986 1043 -964
rect 1058 -986 1088 -964
rect 1115 -986 1116 -970
rect 1131 -986 1144 -826
rect 1174 -930 1187 -826
rect 1232 -848 1233 -838
rect 1248 -848 1261 -838
rect 1232 -854 1261 -848
rect 1216 -862 1261 -854
rect 1216 -874 1241 -862
rect 1248 -874 1261 -862
rect 1216 -882 1261 -874
rect 1232 -890 1233 -882
rect 1248 -890 1261 -882
rect 1232 -898 1248 -890
rect 1229 -905 1248 -902
rect 1229 -914 1251 -905
rect 1202 -924 1251 -914
rect 1202 -930 1232 -924
rect 1251 -929 1256 -924
rect 3379 -930 3408 -914
rect 1174 -946 1248 -930
rect 3379 -946 3424 -930
rect 1174 -948 1187 -946
rect 1202 -948 1236 -946
rect 3379 -948 3412 -946
rect 1174 -964 1248 -948
rect 3379 -964 3424 -948
rect 1158 -986 1159 -970
rect 1174 -986 1187 -964
rect 1202 -986 1232 -964
rect 3379 -986 3408 -964
rect 3435 -986 3436 -970
rect 3451 -986 3464 -887
rect 3494 -930 3507 -887
rect 3552 -890 3553 -887
rect 3568 -890 3581 -887
rect 3552 -898 3568 -890
rect 3549 -905 3568 -902
rect 3549 -914 3571 -905
rect 3522 -924 3571 -914
rect 3522 -930 3552 -924
rect 3571 -929 3576 -924
rect 3494 -946 3568 -930
rect 3586 -938 3616 -887
rect 3651 -892 3859 -887
rect 3677 -922 3866 -892
rect 3692 -925 3866 -922
rect 3685 -928 3866 -925
rect 3494 -948 3507 -946
rect 3522 -948 3556 -946
rect 3494 -964 3568 -948
rect 3595 -952 3608 -938
rect 3623 -952 3639 -936
rect 3685 -941 3696 -928
rect 3478 -986 3479 -970
rect 3494 -986 3507 -964
rect 3522 -986 3552 -964
rect 3595 -968 3657 -952
rect 3685 -959 3696 -943
rect 3701 -948 3711 -928
rect 3721 -948 3735 -928
rect 3738 -941 3747 -928
rect 3763 -941 3772 -928
rect 3701 -959 3735 -948
rect 3738 -959 3747 -943
rect 3763 -959 3772 -943
rect 3779 -948 3789 -928
rect 3799 -948 3813 -928
rect 3814 -941 3825 -928
rect 3779 -959 3813 -948
rect 3814 -959 3825 -943
rect 3871 -952 3887 -936
rect 3894 -938 3924 -887
rect 3958 -890 3959 -887
rect 3943 -898 3959 -890
rect 3930 -930 3943 -911
rect 3958 -930 3988 -914
rect 3930 -946 4004 -930
rect 3930 -948 3943 -946
rect 3958 -948 3992 -946
rect 3595 -970 3608 -968
rect 3623 -970 3657 -968
rect 3595 -986 3657 -970
rect 3701 -975 3717 -968
rect 3779 -975 3809 -964
rect 3857 -968 3903 -952
rect 3930 -964 4004 -948
rect 3857 -970 3891 -968
rect 3856 -986 3903 -970
rect 3930 -986 3943 -964
rect 3958 -986 3988 -964
rect 4015 -986 4016 -970
rect 4031 -986 4044 -887
rect 4074 -930 4087 -887
rect 4132 -890 4133 -887
rect 4148 -890 4161 -887
rect 4132 -898 4148 -890
rect 4129 -905 4148 -902
rect 4129 -914 4151 -905
rect 4102 -924 4151 -914
rect 4102 -930 4132 -924
rect 4151 -929 4156 -924
rect 4074 -946 4148 -930
rect 4166 -938 4196 -887
rect 4231 -892 4439 -887
rect 4257 -922 4446 -892
rect 4272 -925 4446 -922
rect 4265 -928 4446 -925
rect 4074 -948 4087 -946
rect 4102 -948 4136 -946
rect 4074 -964 4148 -948
rect 4175 -952 4188 -938
rect 4203 -952 4219 -936
rect 4265 -941 4276 -928
rect 4058 -986 4059 -970
rect 4074 -986 4087 -964
rect 4102 -986 4132 -964
rect 4175 -968 4237 -952
rect 4265 -959 4276 -943
rect 4281 -948 4291 -928
rect 4301 -948 4315 -928
rect 4318 -941 4327 -928
rect 4343 -941 4352 -928
rect 4281 -959 4315 -948
rect 4318 -959 4327 -943
rect 4343 -959 4352 -943
rect 4359 -948 4369 -928
rect 4379 -948 4393 -928
rect 4394 -941 4405 -928
rect 4359 -959 4393 -948
rect 4394 -959 4405 -943
rect 4451 -952 4467 -936
rect 4474 -938 4504 -887
rect 4538 -890 4539 -887
rect 4523 -898 4539 -890
rect 4510 -930 4523 -911
rect 4538 -930 4568 -914
rect 4510 -946 4584 -930
rect 4510 -948 4523 -946
rect 4538 -948 4572 -946
rect 4175 -970 4188 -968
rect 4203 -970 4237 -968
rect 4175 -986 4237 -970
rect 4281 -975 4297 -968
rect 4359 -975 4389 -964
rect 4437 -968 4483 -952
rect 4510 -964 4584 -948
rect 4437 -970 4471 -968
rect 4436 -986 4483 -970
rect 4510 -986 4523 -964
rect 4538 -986 4568 -964
rect 4595 -986 4596 -970
rect 4611 -986 4624 -887
rect 4654 -931 4667 -887
rect 4712 -891 4713 -887
rect 4728 -891 4741 -887
rect 4712 -899 4728 -891
rect 4709 -906 4728 -903
rect 4709 -915 4731 -906
rect 4682 -925 4731 -915
rect 4682 -931 4712 -925
rect 4731 -930 4736 -925
rect 4654 -947 4728 -931
rect 4746 -939 4776 -887
rect 4811 -893 5019 -887
rect 4837 -923 5026 -893
rect 4852 -926 5026 -923
rect 4845 -929 5026 -926
rect 4654 -949 4667 -947
rect 4682 -949 4716 -947
rect 4654 -965 4728 -949
rect 4755 -953 4768 -939
rect 4783 -953 4799 -937
rect 4845 -942 4856 -929
rect -8 -994 33 -986
rect -8 -1020 7 -994
rect 14 -1020 33 -994
rect 97 -998 159 -986
rect 171 -998 246 -986
rect 304 -998 379 -986
rect 391 -998 422 -986
rect 428 -998 463 -986
rect 97 -1000 259 -998
rect -8 -1028 33 -1020
rect 115 -1024 128 -1000
rect 143 -1002 158 -1000
rect -2 -1038 -1 -1028
rect 14 -1038 27 -1028
rect 42 -1038 72 -1024
rect 115 -1038 158 -1024
rect 182 -1027 189 -1020
rect 192 -1024 259 -1000
rect 291 -1000 463 -998
rect 261 -1022 289 -1018
rect 291 -1022 371 -1000
rect 392 -1002 407 -1000
rect 261 -1024 371 -1022
rect 192 -1028 371 -1024
rect 165 -1038 195 -1028
rect 197 -1038 350 -1028
rect 358 -1038 388 -1028
rect 392 -1038 422 -1024
rect 450 -1038 463 -1000
rect 535 -994 570 -986
rect 535 -1020 536 -994
rect 543 -1020 570 -994
rect 478 -1038 508 -1024
rect 535 -1028 570 -1020
rect 572 -994 613 -986
rect 572 -1020 587 -994
rect 594 -1020 613 -994
rect 677 -998 739 -986
rect 751 -998 826 -986
rect 884 -998 959 -986
rect 971 -998 1002 -986
rect 1008 -998 1043 -986
rect 677 -1000 839 -998
rect 572 -1028 613 -1020
rect 695 -1024 708 -1000
rect 723 -1002 738 -1000
rect 535 -1038 536 -1028
rect 551 -1038 564 -1028
rect 578 -1038 579 -1028
rect 594 -1038 607 -1028
rect 622 -1038 652 -1024
rect 695 -1038 738 -1024
rect 762 -1027 769 -1020
rect 772 -1024 839 -1000
rect 871 -1000 1043 -998
rect 841 -1022 869 -1018
rect 871 -1022 951 -1000
rect 972 -1002 987 -1000
rect 841 -1024 951 -1022
rect 772 -1028 951 -1024
rect 745 -1038 775 -1028
rect 777 -1038 930 -1028
rect 938 -1038 968 -1028
rect 972 -1038 1002 -1024
rect 1030 -1038 1043 -1000
rect 1115 -994 1150 -986
rect 1115 -1020 1116 -994
rect 1123 -1020 1150 -994
rect 1058 -1038 1088 -1024
rect 1115 -1028 1150 -1020
rect 1152 -994 1193 -986
rect 1152 -1020 1167 -994
rect 1174 -1020 1193 -994
rect 1257 -1000 1261 -986
rect 3435 -994 3470 -986
rect 1152 -1028 1193 -1020
rect 3435 -1020 3436 -994
rect 3443 -1020 3470 -994
rect 1115 -1038 1116 -1028
rect 1131 -1038 1144 -1028
rect 1158 -1038 1159 -1028
rect 1174 -1038 1187 -1028
rect 1202 -1038 1232 -1024
rect 3379 -1038 3408 -1024
rect 3435 -1028 3470 -1020
rect 3472 -994 3513 -986
rect 3472 -1020 3487 -994
rect 3494 -1020 3513 -994
rect 3577 -998 3639 -986
rect 3651 -998 3726 -986
rect 3784 -998 3859 -986
rect 3871 -998 3902 -986
rect 3908 -998 3943 -986
rect 3577 -1000 3739 -998
rect 3472 -1028 3513 -1020
rect 3595 -1024 3608 -1000
rect 3623 -1002 3638 -1000
rect 3435 -1038 3436 -1028
rect 3451 -1038 3464 -1028
rect 3478 -1038 3479 -1028
rect 3494 -1038 3507 -1028
rect 3522 -1038 3552 -1024
rect 3595 -1038 3638 -1024
rect 3662 -1027 3669 -1020
rect 3672 -1024 3739 -1000
rect 3771 -1000 3943 -998
rect 3741 -1022 3769 -1018
rect 3771 -1022 3851 -1000
rect 3872 -1002 3887 -1000
rect 3741 -1024 3851 -1022
rect 3672 -1028 3851 -1024
rect 3645 -1038 3675 -1028
rect 3677 -1038 3830 -1028
rect 3838 -1038 3868 -1028
rect 3872 -1038 3902 -1024
rect 3930 -1038 3943 -1000
rect 4015 -994 4050 -986
rect 4015 -1020 4016 -994
rect 4023 -1020 4050 -994
rect 3958 -1038 3988 -1024
rect 4015 -1028 4050 -1020
rect 4052 -994 4093 -986
rect 4052 -1020 4067 -994
rect 4074 -1020 4093 -994
rect 4157 -998 4219 -986
rect 4231 -998 4306 -986
rect 4364 -998 4439 -986
rect 4451 -998 4482 -986
rect 4488 -998 4523 -986
rect 4157 -1000 4319 -998
rect 4052 -1028 4093 -1020
rect 4175 -1024 4188 -1000
rect 4203 -1002 4218 -1000
rect 4015 -1038 4016 -1028
rect 4031 -1038 4044 -1028
rect 4058 -1038 4059 -1028
rect 4074 -1038 4087 -1028
rect 4102 -1038 4132 -1024
rect 4175 -1038 4218 -1024
rect 4242 -1027 4249 -1020
rect 4252 -1024 4319 -1000
rect 4351 -1000 4523 -998
rect 4321 -1022 4349 -1018
rect 4351 -1022 4431 -1000
rect 4452 -1002 4467 -1000
rect 4321 -1024 4431 -1022
rect 4252 -1028 4431 -1024
rect 4225 -1038 4255 -1028
rect 4257 -1038 4410 -1028
rect 4418 -1038 4448 -1028
rect 4452 -1038 4482 -1024
rect 4510 -1038 4523 -1000
rect 4595 -994 4630 -986
rect 4638 -987 4639 -971
rect 4654 -987 4667 -965
rect 4682 -987 4712 -965
rect 4755 -969 4817 -953
rect 4845 -960 4856 -944
rect 4861 -949 4871 -929
rect 4881 -949 4895 -929
rect 4898 -942 4907 -929
rect 4923 -942 4932 -929
rect 4861 -960 4895 -949
rect 4898 -960 4907 -944
rect 4923 -960 4932 -944
rect 4939 -949 4949 -929
rect 4959 -949 4973 -929
rect 4974 -942 4985 -929
rect 4939 -960 4973 -949
rect 4974 -960 4985 -944
rect 5031 -953 5047 -937
rect 5054 -939 5084 -887
rect 5118 -891 5119 -887
rect 5103 -899 5119 -891
rect 5090 -931 5103 -912
rect 5118 -931 5148 -915
rect 5090 -947 5164 -931
rect 5090 -949 5103 -947
rect 5118 -949 5152 -947
rect 4755 -971 4768 -969
rect 4783 -971 4817 -969
rect 4755 -987 4817 -971
rect 4861 -976 4877 -969
rect 4939 -976 4969 -965
rect 5017 -969 5063 -953
rect 5090 -965 5164 -949
rect 5017 -971 5051 -969
rect 5016 -987 5063 -971
rect 5090 -987 5103 -965
rect 5118 -987 5148 -965
rect 5175 -987 5176 -971
rect 5191 -987 5204 -887
rect 5234 -931 5247 -887
rect 5292 -891 5293 -887
rect 5308 -891 5321 -887
rect 5292 -899 5308 -891
rect 5289 -906 5308 -903
rect 5289 -915 5311 -906
rect 5262 -925 5311 -915
rect 5262 -931 5292 -925
rect 5311 -930 5316 -925
rect 5234 -947 5308 -931
rect 5326 -939 5356 -887
rect 5391 -893 5599 -887
rect 5417 -923 5606 -893
rect 5432 -926 5606 -923
rect 5425 -929 5606 -926
rect 5234 -949 5247 -947
rect 5262 -949 5296 -947
rect 5234 -965 5308 -949
rect 5335 -953 5348 -939
rect 5363 -953 5379 -937
rect 5425 -942 5436 -929
rect 5218 -987 5219 -971
rect 5234 -987 5247 -965
rect 5262 -987 5292 -965
rect 5335 -969 5397 -953
rect 5425 -960 5436 -944
rect 5441 -949 5451 -929
rect 5461 -949 5475 -929
rect 5478 -942 5487 -929
rect 5503 -942 5512 -929
rect 5441 -960 5475 -949
rect 5478 -960 5487 -944
rect 5503 -960 5512 -944
rect 5519 -949 5529 -929
rect 5539 -949 5553 -929
rect 5554 -942 5565 -929
rect 5519 -960 5553 -949
rect 5554 -960 5565 -944
rect 5611 -953 5627 -937
rect 5634 -939 5664 -887
rect 5698 -891 5699 -887
rect 5683 -899 5699 -891
rect 5670 -931 5683 -912
rect 5698 -931 5728 -915
rect 5670 -947 5744 -931
rect 5670 -949 5683 -947
rect 5698 -949 5732 -947
rect 5335 -971 5348 -969
rect 5363 -971 5397 -969
rect 5335 -987 5397 -971
rect 5441 -976 5457 -969
rect 5519 -976 5549 -965
rect 5597 -969 5643 -953
rect 5670 -965 5744 -949
rect 5597 -971 5631 -969
rect 5596 -987 5643 -971
rect 5670 -987 5683 -965
rect 5698 -987 5728 -965
rect 5755 -987 5756 -971
rect 5771 -987 5784 -887
rect 5814 -931 5827 -887
rect 5872 -891 5873 -887
rect 5888 -891 5901 -887
rect 5872 -899 5888 -891
rect 5869 -906 5888 -903
rect 5869 -915 5891 -906
rect 5842 -925 5891 -915
rect 5842 -931 5872 -925
rect 5891 -930 5896 -925
rect 5814 -947 5888 -931
rect 5906 -939 5936 -887
rect 5971 -893 6179 -887
rect 5997 -923 6186 -893
rect 6012 -926 6186 -923
rect 6005 -929 6186 -926
rect 5814 -949 5827 -947
rect 5842 -949 5876 -947
rect 5814 -965 5888 -949
rect 5915 -953 5928 -939
rect 5943 -953 5959 -937
rect 6005 -942 6016 -929
rect 5798 -987 5799 -971
rect 5814 -987 5827 -965
rect 5842 -987 5872 -965
rect 5915 -969 5977 -953
rect 6005 -960 6016 -944
rect 6021 -949 6031 -929
rect 6041 -949 6055 -929
rect 6058 -942 6067 -929
rect 6083 -942 6092 -929
rect 6021 -960 6055 -949
rect 6058 -960 6067 -944
rect 6083 -960 6092 -944
rect 6099 -949 6109 -929
rect 6119 -949 6133 -929
rect 6134 -942 6145 -929
rect 6099 -960 6133 -949
rect 6134 -960 6145 -944
rect 6191 -953 6207 -937
rect 6214 -939 6244 -887
rect 6278 -891 6279 -887
rect 6263 -899 6279 -891
rect 6250 -931 6263 -912
rect 6278 -931 6308 -915
rect 6250 -947 6324 -931
rect 6250 -949 6263 -947
rect 6278 -949 6312 -947
rect 5915 -971 5928 -969
rect 5943 -971 5977 -969
rect 5915 -987 5977 -971
rect 6021 -976 6037 -969
rect 6099 -976 6129 -965
rect 6177 -969 6223 -953
rect 6250 -965 6324 -949
rect 6177 -971 6211 -969
rect 6176 -987 6223 -971
rect 6250 -987 6263 -965
rect 6278 -987 6308 -965
rect 6335 -987 6336 -971
rect 6351 -987 6364 -887
rect 6394 -931 6407 -887
rect 6452 -891 6453 -887
rect 6468 -891 6481 -887
rect 6452 -899 6468 -891
rect 6449 -906 6468 -903
rect 6449 -915 6471 -906
rect 6422 -925 6471 -915
rect 6422 -931 6452 -925
rect 6471 -930 6476 -925
rect 6394 -947 6468 -931
rect 6486 -939 6516 -887
rect 6551 -893 6759 -887
rect 6577 -923 6766 -893
rect 6592 -926 6766 -923
rect 6585 -929 6766 -926
rect 6394 -949 6407 -947
rect 6422 -949 6456 -947
rect 6394 -965 6468 -949
rect 6495 -953 6508 -939
rect 6523 -953 6539 -937
rect 6585 -942 6596 -929
rect 6378 -987 6379 -971
rect 6394 -987 6407 -965
rect 6422 -987 6452 -965
rect 6495 -969 6557 -953
rect 6585 -960 6596 -944
rect 6601 -949 6611 -929
rect 6621 -949 6635 -929
rect 6638 -942 6647 -929
rect 6663 -942 6672 -929
rect 6601 -960 6635 -949
rect 6638 -960 6647 -944
rect 6663 -960 6672 -944
rect 6679 -949 6689 -929
rect 6699 -949 6713 -929
rect 6714 -942 6725 -929
rect 6679 -960 6713 -949
rect 6714 -960 6725 -944
rect 6771 -953 6787 -937
rect 6794 -939 6824 -887
rect 6858 -891 6859 -887
rect 6843 -899 6859 -891
rect 6830 -931 6843 -912
rect 6858 -931 6888 -915
rect 6830 -947 6904 -931
rect 6830 -949 6843 -947
rect 6858 -949 6892 -947
rect 6495 -971 6508 -969
rect 6523 -971 6557 -969
rect 6495 -987 6557 -971
rect 6601 -976 6617 -969
rect 6679 -976 6709 -965
rect 6757 -969 6803 -953
rect 6830 -965 6904 -949
rect 6757 -971 6791 -969
rect 6756 -987 6803 -971
rect 6830 -987 6843 -965
rect 6858 -987 6888 -965
rect 6915 -987 6916 -971
rect 6931 -987 6944 -887
rect 4595 -1020 4596 -994
rect 4603 -1020 4630 -994
rect 4538 -1038 4568 -1024
rect 4595 -1028 4630 -1020
rect 4632 -995 4673 -987
rect 4632 -1021 4647 -995
rect 4654 -1021 4673 -995
rect 4737 -999 4799 -987
rect 4811 -999 4886 -987
rect 4944 -999 5019 -987
rect 5031 -999 5062 -987
rect 5068 -999 5103 -987
rect 4737 -1001 4899 -999
rect 4755 -1019 4768 -1001
rect 4783 -1003 4798 -1001
rect 4595 -1038 4596 -1028
rect 4611 -1038 4624 -1028
rect 4632 -1029 4673 -1021
rect 4756 -1025 4768 -1019
rect -2 -1044 1261 -1038
rect -1 -1052 1261 -1044
rect 3379 -1039 4624 -1038
rect 4638 -1039 4639 -1029
rect 4654 -1039 4667 -1029
rect 4682 -1039 4712 -1025
rect 4756 -1039 4798 -1025
rect 4822 -1028 4829 -1021
rect 4832 -1025 4899 -1001
rect 4931 -1001 5103 -999
rect 4901 -1023 4929 -1019
rect 4931 -1023 5011 -1001
rect 5032 -1003 5047 -1001
rect 4901 -1025 5011 -1023
rect 4832 -1029 5011 -1025
rect 4805 -1039 4835 -1029
rect 4837 -1039 4990 -1029
rect 4998 -1039 5028 -1029
rect 5032 -1039 5062 -1025
rect 5090 -1039 5103 -1001
rect 5175 -995 5210 -987
rect 5175 -1021 5176 -995
rect 5183 -1021 5210 -995
rect 5118 -1039 5148 -1025
rect 5175 -1029 5210 -1021
rect 5212 -995 5253 -987
rect 5212 -1021 5227 -995
rect 5234 -1021 5253 -995
rect 5317 -999 5379 -987
rect 5391 -999 5466 -987
rect 5524 -999 5599 -987
rect 5611 -999 5642 -987
rect 5648 -999 5683 -987
rect 5317 -1001 5479 -999
rect 5335 -1019 5348 -1001
rect 5363 -1003 5378 -1001
rect 5212 -1029 5253 -1021
rect 5336 -1025 5348 -1019
rect 5175 -1039 5176 -1029
rect 5191 -1039 5204 -1029
rect 5218 -1039 5219 -1029
rect 5234 -1039 5247 -1029
rect 5262 -1039 5292 -1025
rect 5336 -1039 5378 -1025
rect 5402 -1028 5409 -1021
rect 5412 -1025 5479 -1001
rect 5511 -1001 5683 -999
rect 5481 -1023 5509 -1019
rect 5511 -1023 5591 -1001
rect 5612 -1003 5627 -1001
rect 5481 -1025 5591 -1023
rect 5412 -1029 5591 -1025
rect 5385 -1039 5415 -1029
rect 5417 -1039 5570 -1029
rect 5578 -1039 5608 -1029
rect 5612 -1039 5642 -1025
rect 5670 -1039 5683 -1001
rect 5755 -995 5790 -987
rect 5755 -1021 5756 -995
rect 5763 -1021 5790 -995
rect 5698 -1039 5728 -1025
rect 5755 -1029 5790 -1021
rect 5792 -995 5833 -987
rect 5792 -1021 5807 -995
rect 5814 -1021 5833 -995
rect 5897 -999 5959 -987
rect 5971 -999 6046 -987
rect 6104 -999 6179 -987
rect 6191 -999 6222 -987
rect 6228 -999 6263 -987
rect 5897 -1001 6059 -999
rect 5915 -1019 5928 -1001
rect 5943 -1003 5958 -1001
rect 5792 -1029 5833 -1021
rect 5916 -1025 5928 -1019
rect 5755 -1039 5756 -1029
rect 5771 -1039 5784 -1029
rect 5798 -1039 5799 -1029
rect 5814 -1039 5827 -1029
rect 5842 -1039 5872 -1025
rect 5916 -1039 5958 -1025
rect 5982 -1028 5989 -1021
rect 5992 -1025 6059 -1001
rect 6091 -1001 6263 -999
rect 6061 -1023 6089 -1019
rect 6091 -1023 6171 -1001
rect 6192 -1003 6207 -1001
rect 6061 -1025 6171 -1023
rect 5992 -1029 6171 -1025
rect 5965 -1039 5995 -1029
rect 5997 -1039 6150 -1029
rect 6158 -1039 6188 -1029
rect 6192 -1039 6222 -1025
rect 6250 -1039 6263 -1001
rect 6335 -995 6370 -987
rect 6335 -1021 6336 -995
rect 6343 -1021 6370 -995
rect 6278 -1039 6308 -1025
rect 6335 -1029 6370 -1021
rect 6372 -995 6413 -987
rect 6372 -1021 6387 -995
rect 6394 -1021 6413 -995
rect 6477 -999 6539 -987
rect 6551 -999 6626 -987
rect 6684 -999 6759 -987
rect 6771 -999 6802 -987
rect 6808 -999 6843 -987
rect 6477 -1001 6639 -999
rect 6495 -1019 6508 -1001
rect 6523 -1003 6538 -1001
rect 6372 -1029 6413 -1021
rect 6496 -1025 6508 -1019
rect 6335 -1039 6336 -1029
rect 6351 -1039 6364 -1029
rect 6378 -1039 6379 -1029
rect 6394 -1039 6407 -1029
rect 6422 -1039 6452 -1025
rect 6496 -1039 6538 -1025
rect 6562 -1028 6569 -1021
rect 6572 -1025 6639 -1001
rect 6671 -1001 6843 -999
rect 6641 -1023 6669 -1019
rect 6671 -1023 6751 -1001
rect 6772 -1003 6787 -1001
rect 6641 -1025 6751 -1023
rect 6572 -1029 6751 -1025
rect 6545 -1039 6575 -1029
rect 6577 -1039 6730 -1029
rect 6738 -1039 6768 -1029
rect 6772 -1039 6802 -1025
rect 6830 -1039 6843 -1001
rect 6915 -995 6950 -987
rect 6915 -1021 6916 -995
rect 6923 -1021 6950 -995
rect 6858 -1039 6888 -1025
rect 6915 -1029 6950 -1021
rect 6915 -1039 6916 -1029
rect 6931 -1039 6944 -1029
rect 3379 -1052 6944 -1039
rect 14 -1082 27 -1052
rect 42 -1070 72 -1052
rect 115 -1066 129 -1052
rect 165 -1066 385 -1052
rect 116 -1068 129 -1066
rect 82 -1080 97 -1068
rect 79 -1082 101 -1080
rect 106 -1082 136 -1068
rect 197 -1070 350 -1066
rect 179 -1082 371 -1070
rect 414 -1082 444 -1068
rect 450 -1082 463 -1052
rect 478 -1070 508 -1052
rect 551 -1082 564 -1052
rect 594 -1082 607 -1052
rect 622 -1070 652 -1052
rect 695 -1066 709 -1052
rect 745 -1066 965 -1052
rect 696 -1068 709 -1066
rect 662 -1080 677 -1068
rect 659 -1082 681 -1080
rect 686 -1082 716 -1068
rect 777 -1070 930 -1066
rect 759 -1082 951 -1070
rect 994 -1082 1024 -1068
rect 1030 -1082 1043 -1052
rect 1058 -1070 1088 -1052
rect 1131 -1082 1144 -1052
rect 1174 -1082 1187 -1052
rect 1202 -1070 1232 -1052
rect 1242 -1080 1257 -1068
rect 3379 -1070 3408 -1052
rect 1239 -1082 1261 -1080
rect 3451 -1082 3464 -1052
rect 3494 -1082 3507 -1052
rect 3522 -1070 3552 -1052
rect 3595 -1066 3609 -1052
rect 3645 -1066 3865 -1052
rect 3596 -1068 3609 -1066
rect 3562 -1080 3577 -1068
rect 3559 -1082 3581 -1080
rect 3586 -1082 3616 -1068
rect 3677 -1070 3830 -1066
rect 3659 -1082 3851 -1070
rect 3894 -1082 3924 -1068
rect 3930 -1082 3943 -1052
rect 3958 -1070 3988 -1052
rect 4031 -1082 4044 -1052
rect 4074 -1082 4087 -1052
rect 4102 -1070 4132 -1052
rect 4175 -1066 4189 -1052
rect 4225 -1066 4445 -1052
rect 4176 -1068 4189 -1066
rect 4142 -1080 4157 -1068
rect 4139 -1082 4161 -1080
rect 4166 -1082 4196 -1068
rect 4257 -1070 4410 -1066
rect 4239 -1082 4431 -1070
rect 4474 -1082 4504 -1068
rect 4510 -1082 4523 -1052
rect 4538 -1070 4568 -1052
rect 4611 -1053 6944 -1052
rect 4611 -1082 4624 -1053
rect -1 -1096 1261 -1082
rect 3379 -1083 4624 -1082
rect 4654 -1083 4667 -1053
rect 4682 -1071 4712 -1053
rect 4756 -1069 4769 -1053
rect 4805 -1067 5025 -1053
rect 4722 -1081 4737 -1069
rect 4719 -1083 4741 -1081
rect 4746 -1083 4776 -1069
rect 4837 -1071 4990 -1067
rect 4819 -1083 5011 -1071
rect 5054 -1083 5084 -1069
rect 5090 -1083 5103 -1053
rect 5118 -1071 5148 -1053
rect 5191 -1083 5204 -1053
rect 5234 -1083 5247 -1053
rect 5262 -1071 5292 -1053
rect 5336 -1069 5349 -1053
rect 5385 -1067 5605 -1053
rect 5302 -1081 5317 -1069
rect 5299 -1083 5321 -1081
rect 5326 -1083 5356 -1069
rect 5417 -1071 5570 -1067
rect 5399 -1083 5591 -1071
rect 5634 -1083 5664 -1069
rect 5670 -1083 5683 -1053
rect 5698 -1071 5728 -1053
rect 5771 -1083 5784 -1053
rect 5814 -1083 5827 -1053
rect 5842 -1071 5872 -1053
rect 5916 -1069 5929 -1053
rect 5965 -1067 6185 -1053
rect 5882 -1081 5897 -1069
rect 5879 -1083 5901 -1081
rect 5906 -1083 5936 -1069
rect 5997 -1071 6150 -1067
rect 5979 -1083 6171 -1071
rect 6214 -1083 6244 -1069
rect 6250 -1083 6263 -1053
rect 6278 -1071 6308 -1053
rect 6351 -1083 6364 -1053
rect 6394 -1083 6407 -1053
rect 6422 -1071 6452 -1053
rect 6496 -1069 6509 -1053
rect 6545 -1067 6765 -1053
rect 6462 -1081 6477 -1069
rect 6459 -1083 6481 -1081
rect 6486 -1083 6516 -1069
rect 6577 -1071 6730 -1067
rect 6559 -1083 6751 -1071
rect 6794 -1083 6824 -1069
rect 6830 -1083 6843 -1053
rect 6858 -1071 6888 -1053
rect 6931 -1083 6944 -1053
rect 3379 -1096 6944 -1083
rect 14 -1200 27 -1096
rect 72 -1118 73 -1108
rect 88 -1118 101 -1108
rect 72 -1122 101 -1118
rect 106 -1122 136 -1096
rect 154 -1110 170 -1108
rect 242 -1110 295 -1096
rect 243 -1112 307 -1110
rect 350 -1112 365 -1096
rect 414 -1099 444 -1096
rect 414 -1102 450 -1099
rect 380 -1110 396 -1108
rect 154 -1122 169 -1118
rect 72 -1124 169 -1122
rect 197 -1124 365 -1112
rect 381 -1122 396 -1118
rect 414 -1121 453 -1102
rect 472 -1108 479 -1107
rect 478 -1115 479 -1108
rect 462 -1118 463 -1115
rect 478 -1118 491 -1115
rect 414 -1122 444 -1121
rect 453 -1122 459 -1121
rect 462 -1122 491 -1118
rect 381 -1123 491 -1122
rect 381 -1124 497 -1123
rect 56 -1132 107 -1124
rect 56 -1144 81 -1132
rect 88 -1144 107 -1132
rect 138 -1132 188 -1124
rect 138 -1140 154 -1132
rect 161 -1134 188 -1132
rect 197 -1134 418 -1124
rect 161 -1144 418 -1134
rect 447 -1132 497 -1124
rect 447 -1141 463 -1132
rect 56 -1152 107 -1144
rect 154 -1152 418 -1144
rect 444 -1144 463 -1141
rect 470 -1144 497 -1132
rect 444 -1152 497 -1144
rect 72 -1160 73 -1152
rect 88 -1160 101 -1152
rect 72 -1168 88 -1160
rect 69 -1175 88 -1172
rect 69 -1184 91 -1175
rect 42 -1194 91 -1184
rect 42 -1200 72 -1194
rect 91 -1199 96 -1194
rect 14 -1216 88 -1200
rect 106 -1208 136 -1152
rect 171 -1162 379 -1152
rect 414 -1156 459 -1152
rect 462 -1153 463 -1152
rect 478 -1153 491 -1152
rect 197 -1192 386 -1162
rect 212 -1195 386 -1192
rect 205 -1198 386 -1195
rect 14 -1218 27 -1216
rect 42 -1218 76 -1216
rect 14 -1234 88 -1218
rect 115 -1222 128 -1208
rect 143 -1222 159 -1206
rect 205 -1211 216 -1198
rect -2 -1256 -1 -1240
rect 14 -1256 27 -1234
rect 42 -1256 72 -1234
rect 115 -1238 177 -1222
rect 205 -1229 216 -1213
rect 221 -1218 231 -1198
rect 241 -1218 255 -1198
rect 258 -1211 267 -1198
rect 283 -1211 292 -1198
rect 221 -1229 255 -1218
rect 258 -1229 267 -1213
rect 283 -1229 292 -1213
rect 299 -1218 309 -1198
rect 319 -1218 333 -1198
rect 334 -1211 345 -1198
rect 299 -1229 333 -1218
rect 334 -1229 345 -1213
rect 391 -1222 407 -1206
rect 414 -1208 444 -1156
rect 478 -1160 479 -1153
rect 463 -1168 479 -1160
rect 450 -1200 463 -1181
rect 478 -1200 508 -1184
rect 450 -1216 524 -1200
rect 450 -1218 463 -1216
rect 478 -1218 512 -1216
rect 115 -1240 128 -1238
rect 143 -1240 177 -1238
rect 115 -1256 177 -1240
rect 221 -1245 237 -1238
rect 299 -1245 329 -1234
rect 377 -1238 423 -1222
rect 450 -1234 524 -1218
rect 377 -1240 411 -1238
rect 376 -1256 423 -1240
rect 450 -1256 463 -1234
rect 478 -1256 508 -1234
rect 535 -1256 536 -1240
rect 551 -1256 564 -1096
rect 594 -1200 607 -1096
rect 652 -1118 653 -1108
rect 668 -1118 681 -1108
rect 652 -1122 681 -1118
rect 686 -1122 716 -1096
rect 734 -1110 750 -1108
rect 822 -1110 875 -1096
rect 823 -1112 887 -1110
rect 930 -1112 945 -1096
rect 994 -1099 1024 -1096
rect 994 -1102 1030 -1099
rect 960 -1110 976 -1108
rect 734 -1122 749 -1118
rect 652 -1124 749 -1122
rect 777 -1124 945 -1112
rect 961 -1122 976 -1118
rect 994 -1121 1033 -1102
rect 1052 -1108 1059 -1107
rect 1058 -1115 1059 -1108
rect 1042 -1118 1043 -1115
rect 1058 -1118 1071 -1115
rect 994 -1122 1024 -1121
rect 1033 -1122 1039 -1121
rect 1042 -1122 1071 -1118
rect 961 -1123 1071 -1122
rect 961 -1124 1077 -1123
rect 636 -1132 687 -1124
rect 636 -1144 661 -1132
rect 668 -1144 687 -1132
rect 718 -1132 768 -1124
rect 718 -1140 734 -1132
rect 741 -1134 768 -1132
rect 777 -1134 998 -1124
rect 741 -1144 998 -1134
rect 1027 -1132 1077 -1124
rect 1027 -1141 1043 -1132
rect 636 -1152 687 -1144
rect 734 -1152 998 -1144
rect 1024 -1144 1043 -1141
rect 1050 -1144 1077 -1132
rect 1024 -1152 1077 -1144
rect 652 -1160 653 -1152
rect 668 -1160 681 -1152
rect 652 -1168 668 -1160
rect 649 -1175 668 -1172
rect 649 -1184 671 -1175
rect 622 -1194 671 -1184
rect 622 -1200 652 -1194
rect 671 -1199 676 -1194
rect 594 -1216 668 -1200
rect 686 -1208 716 -1152
rect 751 -1162 959 -1152
rect 994 -1156 1039 -1152
rect 1042 -1153 1043 -1152
rect 1058 -1153 1071 -1152
rect 777 -1192 966 -1162
rect 792 -1195 966 -1192
rect 785 -1198 966 -1195
rect 594 -1218 607 -1216
rect 622 -1218 656 -1216
rect 594 -1234 668 -1218
rect 695 -1222 708 -1208
rect 723 -1222 739 -1206
rect 785 -1211 796 -1198
rect 578 -1256 579 -1240
rect 594 -1256 607 -1234
rect 622 -1256 652 -1234
rect 695 -1238 757 -1222
rect 785 -1229 796 -1213
rect 801 -1218 811 -1198
rect 821 -1218 835 -1198
rect 838 -1211 847 -1198
rect 863 -1211 872 -1198
rect 801 -1229 835 -1218
rect 838 -1229 847 -1213
rect 863 -1229 872 -1213
rect 879 -1218 889 -1198
rect 899 -1218 913 -1198
rect 914 -1211 925 -1198
rect 879 -1229 913 -1218
rect 914 -1229 925 -1213
rect 971 -1222 987 -1206
rect 994 -1208 1024 -1156
rect 1058 -1160 1059 -1153
rect 1043 -1168 1059 -1160
rect 1030 -1200 1043 -1181
rect 1058 -1200 1088 -1184
rect 1030 -1216 1104 -1200
rect 1030 -1218 1043 -1216
rect 1058 -1218 1092 -1216
rect 695 -1240 708 -1238
rect 723 -1240 757 -1238
rect 695 -1256 757 -1240
rect 801 -1245 817 -1238
rect 879 -1245 909 -1234
rect 957 -1238 1003 -1222
rect 1030 -1234 1104 -1218
rect 957 -1240 991 -1238
rect 956 -1256 1003 -1240
rect 1030 -1256 1043 -1234
rect 1058 -1256 1088 -1234
rect 1115 -1256 1116 -1240
rect 1131 -1256 1144 -1096
rect 1174 -1200 1187 -1096
rect 1232 -1118 1233 -1108
rect 1248 -1118 1261 -1108
rect 1232 -1124 1261 -1118
rect 1216 -1132 1261 -1124
rect 1216 -1144 1241 -1132
rect 1248 -1144 1261 -1132
rect 1216 -1152 1261 -1144
rect 1232 -1160 1233 -1152
rect 1248 -1160 1261 -1152
rect 3379 -1123 3391 -1115
rect 3379 -1152 3397 -1123
rect 3379 -1153 3391 -1152
rect 1232 -1168 1248 -1160
rect 1229 -1175 1248 -1172
rect 1229 -1184 1251 -1175
rect 1202 -1194 1251 -1184
rect 1202 -1200 1232 -1194
rect 1251 -1199 1256 -1194
rect 3379 -1200 3408 -1184
rect 1174 -1216 1248 -1200
rect 3379 -1216 3424 -1200
rect 1174 -1218 1187 -1216
rect 1202 -1218 1236 -1216
rect 3379 -1218 3412 -1216
rect 1174 -1234 1248 -1218
rect 3379 -1234 3424 -1218
rect 1158 -1256 1159 -1240
rect 1174 -1256 1187 -1234
rect 1202 -1256 1232 -1234
rect 3379 -1256 3408 -1234
rect 3435 -1256 3436 -1240
rect 3451 -1256 3464 -1096
rect 3494 -1200 3507 -1096
rect 3552 -1118 3553 -1108
rect 3568 -1118 3581 -1108
rect 3552 -1122 3581 -1118
rect 3586 -1122 3616 -1096
rect 3634 -1110 3650 -1108
rect 3722 -1110 3775 -1096
rect 3723 -1112 3787 -1110
rect 3830 -1112 3845 -1096
rect 3894 -1099 3924 -1096
rect 3894 -1102 3930 -1099
rect 3860 -1110 3876 -1108
rect 3634 -1122 3649 -1118
rect 3552 -1124 3649 -1122
rect 3677 -1124 3845 -1112
rect 3861 -1122 3876 -1118
rect 3894 -1121 3933 -1102
rect 3952 -1108 3959 -1107
rect 3958 -1115 3959 -1108
rect 3942 -1118 3943 -1115
rect 3958 -1118 3971 -1115
rect 3894 -1122 3924 -1121
rect 3933 -1122 3939 -1121
rect 3942 -1122 3971 -1118
rect 3861 -1123 3971 -1122
rect 3861 -1124 3977 -1123
rect 3536 -1132 3587 -1124
rect 3536 -1144 3561 -1132
rect 3568 -1144 3587 -1132
rect 3618 -1132 3668 -1124
rect 3618 -1140 3634 -1132
rect 3641 -1134 3668 -1132
rect 3677 -1134 3898 -1124
rect 3641 -1144 3898 -1134
rect 3927 -1132 3977 -1124
rect 3927 -1141 3943 -1132
rect 3536 -1152 3587 -1144
rect 3634 -1152 3898 -1144
rect 3924 -1144 3943 -1141
rect 3950 -1144 3977 -1132
rect 3924 -1152 3977 -1144
rect 3552 -1160 3553 -1152
rect 3568 -1160 3581 -1152
rect 3552 -1168 3568 -1160
rect 3549 -1175 3568 -1172
rect 3549 -1184 3571 -1175
rect 3522 -1194 3571 -1184
rect 3522 -1200 3552 -1194
rect 3571 -1199 3576 -1194
rect 3494 -1216 3568 -1200
rect 3586 -1208 3616 -1152
rect 3651 -1162 3859 -1152
rect 3894 -1156 3939 -1152
rect 3942 -1153 3943 -1152
rect 3958 -1153 3971 -1152
rect 3677 -1192 3866 -1162
rect 3692 -1195 3866 -1192
rect 3685 -1198 3866 -1195
rect 3494 -1218 3507 -1216
rect 3522 -1218 3556 -1216
rect 3494 -1234 3568 -1218
rect 3595 -1222 3608 -1208
rect 3623 -1222 3639 -1206
rect 3685 -1211 3696 -1198
rect 3478 -1256 3479 -1240
rect 3494 -1256 3507 -1234
rect 3522 -1256 3552 -1234
rect 3595 -1238 3657 -1222
rect 3685 -1229 3696 -1213
rect 3701 -1218 3711 -1198
rect 3721 -1218 3735 -1198
rect 3738 -1211 3747 -1198
rect 3763 -1211 3772 -1198
rect 3701 -1229 3735 -1218
rect 3738 -1229 3747 -1213
rect 3763 -1229 3772 -1213
rect 3779 -1218 3789 -1198
rect 3799 -1218 3813 -1198
rect 3814 -1211 3825 -1198
rect 3779 -1229 3813 -1218
rect 3814 -1229 3825 -1213
rect 3871 -1222 3887 -1206
rect 3894 -1208 3924 -1156
rect 3958 -1160 3959 -1153
rect 3943 -1168 3959 -1160
rect 3930 -1200 3943 -1181
rect 3958 -1200 3988 -1184
rect 3930 -1216 4004 -1200
rect 3930 -1218 3943 -1216
rect 3958 -1218 3992 -1216
rect 3595 -1240 3608 -1238
rect 3623 -1240 3657 -1238
rect 3595 -1256 3657 -1240
rect 3701 -1245 3717 -1238
rect 3779 -1245 3809 -1234
rect 3857 -1238 3903 -1222
rect 3930 -1234 4004 -1218
rect 3857 -1240 3891 -1238
rect 3856 -1256 3903 -1240
rect 3930 -1256 3943 -1234
rect 3958 -1256 3988 -1234
rect 4015 -1256 4016 -1240
rect 4031 -1256 4044 -1096
rect 4074 -1200 4087 -1096
rect 4132 -1118 4133 -1108
rect 4148 -1118 4161 -1108
rect 4132 -1122 4161 -1118
rect 4166 -1122 4196 -1096
rect 4214 -1110 4230 -1108
rect 4302 -1110 4355 -1096
rect 4303 -1112 4367 -1110
rect 4410 -1112 4425 -1096
rect 4474 -1099 4504 -1096
rect 4611 -1097 6944 -1096
rect 4474 -1102 4510 -1099
rect 4440 -1110 4456 -1108
rect 4214 -1122 4229 -1118
rect 4132 -1124 4229 -1122
rect 4257 -1124 4425 -1112
rect 4441 -1122 4456 -1118
rect 4474 -1121 4513 -1102
rect 4532 -1108 4539 -1107
rect 4538 -1115 4539 -1108
rect 4522 -1118 4523 -1115
rect 4538 -1118 4551 -1115
rect 4474 -1122 4504 -1121
rect 4513 -1122 4519 -1121
rect 4522 -1122 4551 -1118
rect 4441 -1123 4551 -1122
rect 4441 -1124 4557 -1123
rect 4116 -1132 4167 -1124
rect 4116 -1144 4141 -1132
rect 4148 -1144 4167 -1132
rect 4198 -1132 4248 -1124
rect 4198 -1140 4214 -1132
rect 4221 -1134 4248 -1132
rect 4257 -1134 4478 -1124
rect 4221 -1144 4478 -1134
rect 4507 -1132 4557 -1124
rect 4507 -1141 4523 -1132
rect 4116 -1152 4167 -1144
rect 4214 -1152 4478 -1144
rect 4504 -1144 4523 -1141
rect 4530 -1144 4557 -1132
rect 4504 -1152 4557 -1144
rect 4132 -1160 4133 -1152
rect 4148 -1160 4161 -1152
rect 4132 -1168 4148 -1160
rect 4129 -1175 4148 -1172
rect 4129 -1184 4151 -1175
rect 4102 -1194 4151 -1184
rect 4102 -1200 4132 -1194
rect 4151 -1199 4156 -1194
rect 4074 -1216 4148 -1200
rect 4166 -1208 4196 -1152
rect 4231 -1162 4439 -1152
rect 4474 -1156 4519 -1152
rect 4522 -1153 4523 -1152
rect 4538 -1153 4551 -1152
rect 4257 -1192 4446 -1162
rect 4272 -1195 4446 -1192
rect 4265 -1198 4446 -1195
rect 4074 -1218 4087 -1216
rect 4102 -1218 4136 -1216
rect 4074 -1234 4148 -1218
rect 4175 -1222 4188 -1208
rect 4203 -1222 4219 -1206
rect 4265 -1211 4276 -1198
rect 4058 -1256 4059 -1240
rect 4074 -1256 4087 -1234
rect 4102 -1256 4132 -1234
rect 4175 -1238 4237 -1222
rect 4265 -1229 4276 -1213
rect 4281 -1218 4291 -1198
rect 4301 -1218 4315 -1198
rect 4318 -1211 4327 -1198
rect 4343 -1211 4352 -1198
rect 4281 -1229 4315 -1218
rect 4318 -1229 4327 -1213
rect 4343 -1229 4352 -1213
rect 4359 -1218 4369 -1198
rect 4379 -1218 4393 -1198
rect 4394 -1211 4405 -1198
rect 4359 -1229 4393 -1218
rect 4394 -1229 4405 -1213
rect 4451 -1222 4467 -1206
rect 4474 -1208 4504 -1156
rect 4538 -1160 4539 -1153
rect 4523 -1168 4539 -1160
rect 4510 -1200 4523 -1181
rect 4538 -1200 4568 -1184
rect 4510 -1216 4584 -1200
rect 4510 -1218 4523 -1216
rect 4538 -1218 4572 -1216
rect 4175 -1240 4188 -1238
rect 4203 -1240 4237 -1238
rect 4175 -1256 4237 -1240
rect 4281 -1245 4297 -1238
rect 4359 -1245 4389 -1234
rect 4437 -1238 4483 -1222
rect 4510 -1234 4584 -1218
rect 4437 -1240 4471 -1238
rect 4436 -1256 4483 -1240
rect 4510 -1256 4523 -1234
rect 4538 -1256 4568 -1234
rect 4595 -1256 4596 -1240
rect 4611 -1256 4624 -1097
rect 4654 -1201 4667 -1097
rect 4712 -1119 4713 -1109
rect 4728 -1119 4741 -1109
rect 4712 -1123 4741 -1119
rect 4746 -1123 4776 -1097
rect 4794 -1111 4810 -1109
rect 4882 -1111 4935 -1097
rect 4883 -1113 4947 -1111
rect 4990 -1113 5005 -1097
rect 5054 -1100 5084 -1097
rect 5054 -1103 5090 -1100
rect 5020 -1111 5036 -1109
rect 4794 -1123 4809 -1119
rect 4712 -1125 4809 -1123
rect 4837 -1125 5005 -1113
rect 5021 -1123 5036 -1119
rect 5054 -1122 5093 -1103
rect 5112 -1109 5119 -1108
rect 5118 -1116 5119 -1109
rect 5102 -1119 5103 -1116
rect 5118 -1119 5131 -1116
rect 5054 -1123 5084 -1122
rect 5093 -1123 5099 -1122
rect 5102 -1123 5131 -1119
rect 5021 -1124 5131 -1123
rect 5021 -1125 5137 -1124
rect 4696 -1133 4747 -1125
rect 4696 -1145 4721 -1133
rect 4728 -1145 4747 -1133
rect 4778 -1133 4828 -1125
rect 4778 -1141 4794 -1133
rect 4801 -1135 4828 -1133
rect 4837 -1135 5058 -1125
rect 4801 -1145 5058 -1135
rect 5087 -1133 5137 -1125
rect 5087 -1142 5103 -1133
rect 4696 -1153 4747 -1145
rect 4794 -1153 5058 -1145
rect 5084 -1145 5103 -1142
rect 5110 -1145 5137 -1133
rect 5084 -1153 5137 -1145
rect 4712 -1161 4713 -1153
rect 4728 -1161 4741 -1153
rect 4712 -1169 4728 -1161
rect 4709 -1176 4728 -1173
rect 4709 -1185 4731 -1176
rect 4682 -1195 4731 -1185
rect 4682 -1201 4712 -1195
rect 4731 -1200 4736 -1195
rect 4654 -1217 4728 -1201
rect 4746 -1209 4776 -1153
rect 4811 -1163 5019 -1153
rect 5054 -1157 5099 -1153
rect 5102 -1154 5103 -1153
rect 5118 -1154 5131 -1153
rect 4837 -1193 5026 -1163
rect 4852 -1196 5026 -1193
rect 4845 -1199 5026 -1196
rect 4654 -1219 4667 -1217
rect 4682 -1219 4716 -1217
rect 4654 -1235 4728 -1219
rect 4755 -1223 4768 -1209
rect 4783 -1223 4799 -1207
rect 4845 -1212 4856 -1199
rect -8 -1260 33 -1256
rect 97 -1260 159 -1256
rect 171 -1260 246 -1256
rect 304 -1260 379 -1256
rect 391 -1260 422 -1256
rect 428 -1260 463 -1256
rect 535 -1260 570 -1256
rect 572 -1260 613 -1256
rect 677 -1260 739 -1256
rect 751 -1260 826 -1256
rect 884 -1260 959 -1256
rect 971 -1260 1002 -1256
rect 1008 -1260 1043 -1256
rect 1115 -1260 1150 -1256
rect 1152 -1260 1193 -1256
rect 1257 -1260 1261 -1256
rect 3435 -1264 3470 -1256
rect 3435 -1290 3436 -1264
rect 3443 -1290 3470 -1264
rect 3379 -1308 3408 -1294
rect 3435 -1298 3470 -1290
rect 3472 -1264 3513 -1256
rect 3472 -1290 3487 -1264
rect 3494 -1290 3513 -1264
rect 3577 -1268 3639 -1256
rect 3651 -1268 3726 -1256
rect 3784 -1268 3859 -1256
rect 3871 -1268 3902 -1256
rect 3908 -1268 3943 -1256
rect 3577 -1270 3739 -1268
rect 3472 -1298 3513 -1290
rect 3595 -1294 3608 -1270
rect 3623 -1272 3638 -1270
rect 3435 -1308 3436 -1298
rect 3451 -1308 3464 -1298
rect 3478 -1308 3479 -1298
rect 3494 -1308 3507 -1298
rect 3522 -1308 3552 -1294
rect 3595 -1308 3638 -1294
rect 3662 -1297 3669 -1290
rect 3672 -1294 3739 -1270
rect 3771 -1270 3943 -1268
rect 3741 -1292 3769 -1288
rect 3771 -1292 3851 -1270
rect 3872 -1272 3887 -1270
rect 3741 -1294 3851 -1292
rect 3672 -1298 3851 -1294
rect 3645 -1308 3675 -1298
rect 3677 -1308 3830 -1298
rect 3838 -1308 3868 -1298
rect 3872 -1308 3902 -1294
rect 3930 -1308 3943 -1270
rect 4015 -1264 4050 -1256
rect 4015 -1290 4016 -1264
rect 4023 -1290 4050 -1264
rect 3958 -1308 3988 -1294
rect 4015 -1298 4050 -1290
rect 4052 -1264 4093 -1256
rect 4052 -1290 4067 -1264
rect 4074 -1290 4093 -1264
rect 4157 -1268 4219 -1256
rect 4231 -1268 4306 -1256
rect 4364 -1268 4439 -1256
rect 4451 -1268 4482 -1256
rect 4488 -1268 4523 -1256
rect 4157 -1270 4319 -1268
rect 4052 -1298 4093 -1290
rect 4175 -1294 4188 -1270
rect 4203 -1272 4218 -1270
rect 4015 -1308 4016 -1298
rect 4031 -1308 4044 -1298
rect 4058 -1308 4059 -1298
rect 4074 -1308 4087 -1298
rect 4102 -1308 4132 -1294
rect 4175 -1308 4218 -1294
rect 4242 -1297 4249 -1290
rect 4252 -1294 4319 -1270
rect 4351 -1270 4523 -1268
rect 4321 -1292 4349 -1288
rect 4351 -1292 4431 -1270
rect 4452 -1272 4467 -1270
rect 4321 -1294 4431 -1292
rect 4252 -1298 4431 -1294
rect 4225 -1308 4255 -1298
rect 4257 -1308 4410 -1298
rect 4418 -1308 4448 -1298
rect 4452 -1308 4482 -1294
rect 4510 -1308 4523 -1270
rect 4595 -1264 4630 -1256
rect 4638 -1257 4639 -1241
rect 4654 -1257 4667 -1235
rect 4682 -1257 4712 -1235
rect 4755 -1239 4817 -1223
rect 4845 -1230 4856 -1214
rect 4861 -1219 4871 -1199
rect 4881 -1219 4895 -1199
rect 4898 -1212 4907 -1199
rect 4923 -1212 4932 -1199
rect 4861 -1230 4895 -1219
rect 4898 -1230 4907 -1214
rect 4923 -1230 4932 -1214
rect 4939 -1219 4949 -1199
rect 4959 -1219 4973 -1199
rect 4974 -1212 4985 -1199
rect 4939 -1230 4973 -1219
rect 4974 -1230 4985 -1214
rect 5031 -1223 5047 -1207
rect 5054 -1209 5084 -1157
rect 5118 -1161 5119 -1154
rect 5103 -1169 5119 -1161
rect 5090 -1201 5103 -1182
rect 5118 -1201 5148 -1185
rect 5090 -1217 5164 -1201
rect 5090 -1219 5103 -1217
rect 5118 -1219 5152 -1217
rect 4755 -1241 4768 -1239
rect 4783 -1241 4817 -1239
rect 4755 -1257 4817 -1241
rect 4861 -1246 4877 -1239
rect 4939 -1246 4969 -1235
rect 5017 -1239 5063 -1223
rect 5090 -1235 5164 -1219
rect 5017 -1241 5051 -1239
rect 5016 -1257 5063 -1241
rect 5090 -1257 5103 -1235
rect 5118 -1257 5148 -1235
rect 5175 -1257 5176 -1241
rect 5191 -1257 5204 -1097
rect 5234 -1201 5247 -1097
rect 5292 -1119 5293 -1109
rect 5308 -1119 5321 -1109
rect 5292 -1123 5321 -1119
rect 5326 -1123 5356 -1097
rect 5374 -1111 5390 -1109
rect 5462 -1111 5515 -1097
rect 5463 -1113 5527 -1111
rect 5570 -1113 5585 -1097
rect 5634 -1100 5664 -1097
rect 5634 -1103 5670 -1100
rect 5600 -1111 5616 -1109
rect 5374 -1123 5389 -1119
rect 5292 -1125 5389 -1123
rect 5417 -1125 5585 -1113
rect 5601 -1123 5616 -1119
rect 5634 -1122 5673 -1103
rect 5692 -1109 5699 -1108
rect 5698 -1116 5699 -1109
rect 5682 -1119 5683 -1116
rect 5698 -1119 5711 -1116
rect 5634 -1123 5664 -1122
rect 5673 -1123 5679 -1122
rect 5682 -1123 5711 -1119
rect 5601 -1124 5711 -1123
rect 5601 -1125 5717 -1124
rect 5276 -1133 5327 -1125
rect 5276 -1145 5301 -1133
rect 5308 -1145 5327 -1133
rect 5358 -1133 5408 -1125
rect 5358 -1141 5374 -1133
rect 5381 -1135 5408 -1133
rect 5417 -1135 5638 -1125
rect 5381 -1145 5638 -1135
rect 5667 -1133 5717 -1125
rect 5667 -1142 5683 -1133
rect 5276 -1153 5327 -1145
rect 5374 -1153 5638 -1145
rect 5664 -1145 5683 -1142
rect 5690 -1145 5717 -1133
rect 5664 -1153 5717 -1145
rect 5292 -1161 5293 -1153
rect 5308 -1161 5321 -1153
rect 5292 -1169 5308 -1161
rect 5289 -1176 5308 -1173
rect 5289 -1185 5311 -1176
rect 5262 -1195 5311 -1185
rect 5262 -1201 5292 -1195
rect 5311 -1200 5316 -1195
rect 5234 -1217 5308 -1201
rect 5326 -1209 5356 -1153
rect 5391 -1163 5599 -1153
rect 5634 -1157 5679 -1153
rect 5682 -1154 5683 -1153
rect 5698 -1154 5711 -1153
rect 5417 -1193 5606 -1163
rect 5432 -1196 5606 -1193
rect 5425 -1199 5606 -1196
rect 5234 -1219 5247 -1217
rect 5262 -1219 5296 -1217
rect 5234 -1235 5308 -1219
rect 5335 -1223 5348 -1209
rect 5363 -1223 5379 -1207
rect 5425 -1212 5436 -1199
rect 5218 -1257 5219 -1241
rect 5234 -1257 5247 -1235
rect 5262 -1257 5292 -1235
rect 5335 -1239 5397 -1223
rect 5425 -1230 5436 -1214
rect 5441 -1219 5451 -1199
rect 5461 -1219 5475 -1199
rect 5478 -1212 5487 -1199
rect 5503 -1212 5512 -1199
rect 5441 -1230 5475 -1219
rect 5478 -1230 5487 -1214
rect 5503 -1230 5512 -1214
rect 5519 -1219 5529 -1199
rect 5539 -1219 5553 -1199
rect 5554 -1212 5565 -1199
rect 5519 -1230 5553 -1219
rect 5554 -1230 5565 -1214
rect 5611 -1223 5627 -1207
rect 5634 -1209 5664 -1157
rect 5698 -1161 5699 -1154
rect 5683 -1169 5699 -1161
rect 5670 -1201 5683 -1182
rect 5698 -1201 5728 -1185
rect 5670 -1217 5744 -1201
rect 5670 -1219 5683 -1217
rect 5698 -1219 5732 -1217
rect 5335 -1241 5348 -1239
rect 5363 -1241 5397 -1239
rect 5335 -1257 5397 -1241
rect 5441 -1246 5457 -1239
rect 5519 -1246 5549 -1235
rect 5597 -1239 5643 -1223
rect 5670 -1235 5744 -1219
rect 5597 -1241 5631 -1239
rect 5596 -1257 5643 -1241
rect 5670 -1257 5683 -1235
rect 5698 -1257 5728 -1235
rect 5755 -1257 5756 -1241
rect 5771 -1257 5784 -1097
rect 5814 -1201 5827 -1097
rect 5872 -1119 5873 -1109
rect 5888 -1119 5901 -1109
rect 5872 -1123 5901 -1119
rect 5906 -1123 5936 -1097
rect 5954 -1111 5970 -1109
rect 6042 -1111 6095 -1097
rect 6043 -1113 6107 -1111
rect 6150 -1113 6165 -1097
rect 6214 -1100 6244 -1097
rect 6214 -1103 6250 -1100
rect 6180 -1111 6196 -1109
rect 5954 -1123 5969 -1119
rect 5872 -1125 5969 -1123
rect 5997 -1125 6165 -1113
rect 6181 -1123 6196 -1119
rect 6214 -1122 6253 -1103
rect 6272 -1109 6279 -1108
rect 6278 -1116 6279 -1109
rect 6262 -1119 6263 -1116
rect 6278 -1119 6291 -1116
rect 6214 -1123 6244 -1122
rect 6253 -1123 6259 -1122
rect 6262 -1123 6291 -1119
rect 6181 -1124 6291 -1123
rect 6181 -1125 6297 -1124
rect 5856 -1133 5907 -1125
rect 5856 -1145 5881 -1133
rect 5888 -1145 5907 -1133
rect 5938 -1133 5988 -1125
rect 5938 -1141 5954 -1133
rect 5961 -1135 5988 -1133
rect 5997 -1135 6218 -1125
rect 5961 -1145 6218 -1135
rect 6247 -1133 6297 -1125
rect 6247 -1142 6263 -1133
rect 5856 -1153 5907 -1145
rect 5954 -1153 6218 -1145
rect 6244 -1145 6263 -1142
rect 6270 -1145 6297 -1133
rect 6244 -1153 6297 -1145
rect 5872 -1161 5873 -1153
rect 5888 -1161 5901 -1153
rect 5872 -1169 5888 -1161
rect 5869 -1176 5888 -1173
rect 5869 -1185 5891 -1176
rect 5842 -1195 5891 -1185
rect 5842 -1201 5872 -1195
rect 5891 -1200 5896 -1195
rect 5814 -1217 5888 -1201
rect 5906 -1209 5936 -1153
rect 5971 -1163 6179 -1153
rect 6214 -1157 6259 -1153
rect 6262 -1154 6263 -1153
rect 6278 -1154 6291 -1153
rect 5997 -1193 6186 -1163
rect 6012 -1196 6186 -1193
rect 6005 -1199 6186 -1196
rect 5814 -1219 5827 -1217
rect 5842 -1219 5876 -1217
rect 5814 -1235 5888 -1219
rect 5915 -1223 5928 -1209
rect 5943 -1223 5959 -1207
rect 6005 -1212 6016 -1199
rect 5798 -1257 5799 -1241
rect 5814 -1257 5827 -1235
rect 5842 -1257 5872 -1235
rect 5915 -1239 5977 -1223
rect 6005 -1230 6016 -1214
rect 6021 -1219 6031 -1199
rect 6041 -1219 6055 -1199
rect 6058 -1212 6067 -1199
rect 6083 -1212 6092 -1199
rect 6021 -1230 6055 -1219
rect 6058 -1230 6067 -1214
rect 6083 -1230 6092 -1214
rect 6099 -1219 6109 -1199
rect 6119 -1219 6133 -1199
rect 6134 -1212 6145 -1199
rect 6099 -1230 6133 -1219
rect 6134 -1230 6145 -1214
rect 6191 -1223 6207 -1207
rect 6214 -1209 6244 -1157
rect 6278 -1161 6279 -1154
rect 6263 -1169 6279 -1161
rect 6250 -1201 6263 -1182
rect 6278 -1201 6308 -1185
rect 6250 -1217 6324 -1201
rect 6250 -1219 6263 -1217
rect 6278 -1219 6312 -1217
rect 5915 -1241 5928 -1239
rect 5943 -1241 5977 -1239
rect 5915 -1257 5977 -1241
rect 6021 -1246 6037 -1239
rect 6099 -1246 6129 -1235
rect 6177 -1239 6223 -1223
rect 6250 -1235 6324 -1219
rect 6177 -1241 6211 -1239
rect 6176 -1257 6223 -1241
rect 6250 -1257 6263 -1235
rect 6278 -1257 6308 -1235
rect 6335 -1257 6336 -1241
rect 6351 -1257 6364 -1097
rect 6394 -1201 6407 -1097
rect 6452 -1119 6453 -1109
rect 6468 -1119 6481 -1109
rect 6452 -1123 6481 -1119
rect 6486 -1123 6516 -1097
rect 6534 -1111 6550 -1109
rect 6622 -1111 6675 -1097
rect 6623 -1113 6687 -1111
rect 6730 -1113 6745 -1097
rect 6794 -1100 6824 -1097
rect 6794 -1103 6830 -1100
rect 6760 -1111 6776 -1109
rect 6534 -1123 6549 -1119
rect 6452 -1125 6549 -1123
rect 6577 -1125 6745 -1113
rect 6761 -1123 6776 -1119
rect 6794 -1122 6833 -1103
rect 6852 -1109 6859 -1108
rect 6858 -1116 6859 -1109
rect 6842 -1119 6843 -1116
rect 6858 -1119 6871 -1116
rect 6794 -1123 6824 -1122
rect 6833 -1123 6839 -1122
rect 6842 -1123 6871 -1119
rect 6761 -1124 6871 -1123
rect 6761 -1125 6877 -1124
rect 6436 -1133 6487 -1125
rect 6436 -1145 6461 -1133
rect 6468 -1145 6487 -1133
rect 6518 -1133 6568 -1125
rect 6518 -1141 6534 -1133
rect 6541 -1135 6568 -1133
rect 6577 -1135 6798 -1125
rect 6541 -1145 6798 -1135
rect 6827 -1133 6877 -1125
rect 6827 -1142 6843 -1133
rect 6436 -1153 6487 -1145
rect 6534 -1153 6798 -1145
rect 6824 -1145 6843 -1142
rect 6850 -1145 6877 -1133
rect 6824 -1153 6877 -1145
rect 6452 -1161 6453 -1153
rect 6468 -1161 6481 -1153
rect 6452 -1169 6468 -1161
rect 6449 -1176 6468 -1173
rect 6449 -1185 6471 -1176
rect 6422 -1195 6471 -1185
rect 6422 -1201 6452 -1195
rect 6471 -1200 6476 -1195
rect 6394 -1217 6468 -1201
rect 6486 -1209 6516 -1153
rect 6551 -1163 6759 -1153
rect 6794 -1157 6839 -1153
rect 6842 -1154 6843 -1153
rect 6858 -1154 6871 -1153
rect 6577 -1193 6766 -1163
rect 6592 -1196 6766 -1193
rect 6585 -1199 6766 -1196
rect 6394 -1219 6407 -1217
rect 6422 -1219 6456 -1217
rect 6394 -1235 6468 -1219
rect 6495 -1223 6508 -1209
rect 6523 -1223 6539 -1207
rect 6585 -1212 6596 -1199
rect 6378 -1257 6379 -1241
rect 6394 -1257 6407 -1235
rect 6422 -1257 6452 -1235
rect 6495 -1239 6557 -1223
rect 6585 -1230 6596 -1214
rect 6601 -1219 6611 -1199
rect 6621 -1219 6635 -1199
rect 6638 -1212 6647 -1199
rect 6663 -1212 6672 -1199
rect 6601 -1230 6635 -1219
rect 6638 -1230 6647 -1214
rect 6663 -1230 6672 -1214
rect 6679 -1219 6689 -1199
rect 6699 -1219 6713 -1199
rect 6714 -1212 6725 -1199
rect 6679 -1230 6713 -1219
rect 6714 -1230 6725 -1214
rect 6771 -1223 6787 -1207
rect 6794 -1209 6824 -1157
rect 6858 -1161 6859 -1154
rect 6843 -1169 6859 -1161
rect 6830 -1201 6843 -1182
rect 6858 -1201 6888 -1185
rect 6830 -1217 6904 -1201
rect 6830 -1219 6843 -1217
rect 6858 -1219 6892 -1217
rect 6495 -1241 6508 -1239
rect 6523 -1241 6557 -1239
rect 6495 -1257 6557 -1241
rect 6601 -1246 6617 -1239
rect 6679 -1246 6709 -1235
rect 6757 -1239 6803 -1223
rect 6830 -1235 6904 -1219
rect 6757 -1241 6791 -1239
rect 6756 -1257 6803 -1241
rect 6830 -1257 6843 -1235
rect 6858 -1257 6888 -1235
rect 6915 -1257 6916 -1241
rect 6931 -1257 6944 -1097
rect 4595 -1290 4596 -1264
rect 4603 -1290 4630 -1264
rect 4538 -1308 4568 -1294
rect 4595 -1298 4630 -1290
rect 4632 -1265 4673 -1257
rect 4632 -1291 4647 -1265
rect 4654 -1291 4673 -1265
rect 4737 -1269 4799 -1257
rect 4811 -1269 4886 -1257
rect 4944 -1269 5019 -1257
rect 5031 -1269 5062 -1257
rect 5068 -1269 5103 -1257
rect 4737 -1271 4899 -1269
rect 4595 -1308 4596 -1298
rect 4611 -1308 4624 -1298
rect 4632 -1299 4673 -1291
rect 4755 -1295 4768 -1271
rect 4783 -1273 4798 -1271
rect 3379 -1309 4624 -1308
rect 4638 -1309 4639 -1299
rect 4654 -1309 4667 -1299
rect 4682 -1309 4712 -1295
rect 4755 -1309 4798 -1295
rect 4822 -1298 4829 -1291
rect 4832 -1295 4899 -1271
rect 4931 -1271 5103 -1269
rect 4901 -1293 4929 -1289
rect 4931 -1293 5011 -1271
rect 5032 -1273 5047 -1271
rect 4901 -1295 5011 -1293
rect 4832 -1299 5011 -1295
rect 4805 -1309 4835 -1299
rect 4837 -1309 4990 -1299
rect 4998 -1309 5028 -1299
rect 5032 -1309 5062 -1295
rect 5090 -1309 5103 -1271
rect 5175 -1265 5210 -1257
rect 5175 -1291 5176 -1265
rect 5183 -1291 5210 -1265
rect 5118 -1309 5148 -1295
rect 5175 -1299 5210 -1291
rect 5212 -1265 5253 -1257
rect 5212 -1291 5227 -1265
rect 5234 -1291 5253 -1265
rect 5317 -1269 5379 -1257
rect 5391 -1269 5466 -1257
rect 5524 -1269 5599 -1257
rect 5611 -1269 5642 -1257
rect 5648 -1269 5683 -1257
rect 5317 -1271 5479 -1269
rect 5212 -1299 5253 -1291
rect 5335 -1295 5348 -1271
rect 5363 -1273 5378 -1271
rect 5175 -1309 5176 -1299
rect 5191 -1309 5204 -1299
rect 5218 -1309 5219 -1299
rect 5234 -1309 5247 -1299
rect 5262 -1309 5292 -1295
rect 5335 -1309 5378 -1295
rect 5402 -1298 5409 -1291
rect 5412 -1295 5479 -1271
rect 5511 -1271 5683 -1269
rect 5481 -1293 5509 -1289
rect 5511 -1293 5591 -1271
rect 5612 -1273 5627 -1271
rect 5481 -1295 5591 -1293
rect 5412 -1299 5591 -1295
rect 5385 -1309 5415 -1299
rect 5417 -1309 5570 -1299
rect 5578 -1309 5608 -1299
rect 5612 -1309 5642 -1295
rect 5670 -1309 5683 -1271
rect 5755 -1265 5790 -1257
rect 5755 -1291 5756 -1265
rect 5763 -1291 5790 -1265
rect 5698 -1309 5728 -1295
rect 5755 -1299 5790 -1291
rect 5792 -1265 5833 -1257
rect 5792 -1291 5807 -1265
rect 5814 -1291 5833 -1265
rect 5897 -1269 5959 -1257
rect 5971 -1269 6046 -1257
rect 6104 -1269 6179 -1257
rect 6191 -1269 6222 -1257
rect 6228 -1269 6263 -1257
rect 5897 -1271 6059 -1269
rect 5792 -1299 5833 -1291
rect 5915 -1295 5928 -1271
rect 5943 -1273 5958 -1271
rect 5755 -1309 5756 -1299
rect 5771 -1309 5784 -1299
rect 5798 -1309 5799 -1299
rect 5814 -1309 5827 -1299
rect 5842 -1309 5872 -1295
rect 5915 -1309 5958 -1295
rect 5982 -1298 5989 -1291
rect 5992 -1295 6059 -1271
rect 6091 -1271 6263 -1269
rect 6061 -1293 6089 -1289
rect 6091 -1293 6171 -1271
rect 6192 -1273 6207 -1271
rect 6061 -1295 6171 -1293
rect 5992 -1299 6171 -1295
rect 5965 -1309 5995 -1299
rect 5997 -1309 6150 -1299
rect 6158 -1309 6188 -1299
rect 6192 -1309 6222 -1295
rect 6250 -1309 6263 -1271
rect 6335 -1265 6370 -1257
rect 6335 -1291 6336 -1265
rect 6343 -1291 6370 -1265
rect 6278 -1309 6308 -1295
rect 6335 -1299 6370 -1291
rect 6372 -1265 6413 -1257
rect 6372 -1291 6387 -1265
rect 6394 -1291 6413 -1265
rect 6477 -1269 6539 -1257
rect 6551 -1269 6626 -1257
rect 6684 -1269 6759 -1257
rect 6771 -1269 6802 -1257
rect 6808 -1269 6843 -1257
rect 6477 -1271 6639 -1269
rect 6372 -1299 6413 -1291
rect 6495 -1295 6508 -1271
rect 6523 -1273 6538 -1271
rect 6335 -1309 6336 -1299
rect 6351 -1309 6364 -1299
rect 6378 -1309 6379 -1299
rect 6394 -1309 6407 -1299
rect 6422 -1309 6452 -1295
rect 6495 -1309 6538 -1295
rect 6562 -1298 6569 -1291
rect 6572 -1295 6639 -1271
rect 6671 -1271 6843 -1269
rect 6641 -1293 6669 -1289
rect 6671 -1293 6751 -1271
rect 6772 -1273 6787 -1271
rect 6641 -1295 6751 -1293
rect 6572 -1299 6751 -1295
rect 6545 -1309 6575 -1299
rect 6577 -1309 6730 -1299
rect 6738 -1309 6768 -1299
rect 6772 -1309 6802 -1295
rect 6830 -1309 6843 -1271
rect 6915 -1265 6950 -1257
rect 6915 -1291 6916 -1265
rect 6923 -1291 6950 -1265
rect 6858 -1309 6888 -1295
rect 6915 -1299 6950 -1291
rect 6915 -1309 6916 -1299
rect 6931 -1309 6944 -1299
rect 3379 -1322 6944 -1309
rect 3379 -1340 3408 -1322
rect 3451 -1352 3464 -1322
rect 3494 -1352 3507 -1322
rect 3522 -1340 3552 -1322
rect 3595 -1336 3609 -1322
rect 3645 -1336 3865 -1322
rect 3596 -1338 3609 -1336
rect 3562 -1350 3577 -1338
rect 3559 -1352 3581 -1350
rect 3586 -1352 3616 -1338
rect 3677 -1340 3830 -1336
rect 3659 -1352 3851 -1340
rect 3894 -1352 3924 -1338
rect 3930 -1352 3943 -1322
rect 3958 -1340 3988 -1322
rect 4031 -1352 4044 -1322
rect 4074 -1352 4087 -1322
rect 4102 -1340 4132 -1322
rect 4175 -1336 4189 -1322
rect 4225 -1336 4445 -1322
rect 4176 -1338 4189 -1336
rect 4142 -1350 4157 -1338
rect 4139 -1352 4161 -1350
rect 4166 -1352 4196 -1338
rect 4257 -1340 4410 -1336
rect 4239 -1352 4431 -1340
rect 4474 -1352 4504 -1338
rect 4510 -1352 4523 -1322
rect 4538 -1340 4568 -1322
rect 4611 -1323 6944 -1322
rect 4611 -1352 4624 -1323
rect 3379 -1353 4624 -1352
rect 4654 -1353 4667 -1323
rect 4682 -1341 4712 -1323
rect 4755 -1337 4769 -1323
rect 4805 -1337 5025 -1323
rect 4756 -1339 4769 -1337
rect 4722 -1351 4737 -1339
rect 4719 -1353 4741 -1351
rect 4746 -1353 4776 -1339
rect 4837 -1341 4990 -1337
rect 4819 -1353 5011 -1341
rect 5054 -1353 5084 -1339
rect 5090 -1353 5103 -1323
rect 5118 -1341 5148 -1323
rect 5191 -1353 5204 -1323
rect 5234 -1353 5247 -1323
rect 5262 -1341 5292 -1323
rect 5335 -1337 5349 -1323
rect 5385 -1337 5605 -1323
rect 5336 -1339 5349 -1337
rect 5302 -1351 5317 -1339
rect 5299 -1353 5321 -1351
rect 5326 -1353 5356 -1339
rect 5417 -1341 5570 -1337
rect 5399 -1353 5591 -1341
rect 5634 -1353 5664 -1339
rect 5670 -1353 5683 -1323
rect 5698 -1341 5728 -1323
rect 5771 -1353 5784 -1323
rect 5814 -1353 5827 -1323
rect 5842 -1341 5872 -1323
rect 5915 -1337 5929 -1323
rect 5965 -1337 6185 -1323
rect 5916 -1339 5929 -1337
rect 5882 -1351 5897 -1339
rect 5879 -1353 5901 -1351
rect 5906 -1353 5936 -1339
rect 5997 -1341 6150 -1337
rect 5979 -1353 6171 -1341
rect 6214 -1353 6244 -1339
rect 6250 -1353 6263 -1323
rect 6278 -1341 6308 -1323
rect 6351 -1353 6364 -1323
rect 6394 -1353 6407 -1323
rect 6422 -1341 6452 -1323
rect 6495 -1337 6509 -1323
rect 6545 -1337 6765 -1323
rect 6496 -1339 6509 -1337
rect 6462 -1351 6477 -1339
rect 6459 -1353 6481 -1351
rect 6486 -1353 6516 -1339
rect 6577 -1341 6730 -1337
rect 6559 -1353 6751 -1341
rect 6794 -1353 6824 -1339
rect 6830 -1353 6843 -1323
rect 6858 -1341 6888 -1323
rect 6931 -1353 6944 -1323
rect 3379 -1366 6944 -1353
rect 3379 -1393 3391 -1385
rect 3379 -1422 3397 -1393
rect 3379 -1423 3391 -1422
rect 3379 -1470 3408 -1454
rect 3379 -1486 3424 -1470
rect 3379 -1488 3412 -1486
rect 3379 -1504 3424 -1488
rect 3379 -1526 3408 -1504
rect 3435 -1526 3436 -1510
rect 3451 -1526 3464 -1366
rect 3494 -1470 3507 -1366
rect 3552 -1388 3553 -1378
rect 3568 -1388 3581 -1378
rect 3552 -1392 3581 -1388
rect 3586 -1392 3616 -1366
rect 3634 -1380 3650 -1378
rect 3722 -1380 3775 -1366
rect 3723 -1382 3787 -1380
rect 3830 -1382 3845 -1366
rect 3894 -1369 3924 -1366
rect 3894 -1372 3930 -1369
rect 3860 -1380 3876 -1378
rect 3634 -1392 3649 -1388
rect 3552 -1394 3649 -1392
rect 3677 -1394 3845 -1382
rect 3861 -1392 3876 -1388
rect 3894 -1391 3933 -1372
rect 3952 -1378 3959 -1377
rect 3958 -1385 3959 -1378
rect 3942 -1388 3943 -1385
rect 3958 -1388 3971 -1385
rect 3894 -1392 3924 -1391
rect 3933 -1392 3939 -1391
rect 3942 -1392 3971 -1388
rect 3861 -1393 3971 -1392
rect 3861 -1394 3977 -1393
rect 3536 -1402 3587 -1394
rect 3536 -1414 3561 -1402
rect 3568 -1414 3587 -1402
rect 3618 -1402 3668 -1394
rect 3618 -1410 3634 -1402
rect 3641 -1404 3668 -1402
rect 3677 -1404 3898 -1394
rect 3641 -1414 3898 -1404
rect 3927 -1402 3977 -1394
rect 3927 -1411 3943 -1402
rect 3536 -1422 3587 -1414
rect 3634 -1422 3898 -1414
rect 3924 -1414 3943 -1411
rect 3950 -1414 3977 -1402
rect 3924 -1422 3977 -1414
rect 3552 -1430 3553 -1422
rect 3568 -1430 3581 -1422
rect 3552 -1438 3568 -1430
rect 3549 -1445 3568 -1442
rect 3549 -1454 3571 -1445
rect 3522 -1464 3571 -1454
rect 3522 -1470 3552 -1464
rect 3571 -1469 3576 -1464
rect 3494 -1486 3568 -1470
rect 3586 -1478 3616 -1422
rect 3651 -1432 3859 -1422
rect 3894 -1426 3939 -1422
rect 3942 -1423 3943 -1422
rect 3958 -1423 3971 -1422
rect 3677 -1462 3866 -1432
rect 3692 -1465 3866 -1462
rect 3685 -1468 3866 -1465
rect 3494 -1488 3507 -1486
rect 3522 -1488 3556 -1486
rect 3494 -1504 3568 -1488
rect 3595 -1492 3608 -1478
rect 3623 -1492 3639 -1476
rect 3685 -1481 3696 -1468
rect 3478 -1526 3479 -1510
rect 3494 -1526 3507 -1504
rect 3522 -1526 3552 -1504
rect 3595 -1508 3657 -1492
rect 3685 -1499 3696 -1483
rect 3701 -1488 3711 -1468
rect 3721 -1488 3735 -1468
rect 3738 -1481 3747 -1468
rect 3763 -1481 3772 -1468
rect 3701 -1499 3735 -1488
rect 3738 -1499 3747 -1483
rect 3763 -1499 3772 -1483
rect 3779 -1488 3789 -1468
rect 3799 -1488 3813 -1468
rect 3814 -1481 3825 -1468
rect 3779 -1499 3813 -1488
rect 3814 -1499 3825 -1483
rect 3871 -1492 3887 -1476
rect 3894 -1478 3924 -1426
rect 3958 -1430 3959 -1423
rect 3943 -1438 3959 -1430
rect 3930 -1470 3943 -1451
rect 3958 -1470 3988 -1454
rect 3930 -1486 4004 -1470
rect 3930 -1488 3943 -1486
rect 3958 -1488 3992 -1486
rect 3595 -1510 3608 -1508
rect 3623 -1510 3657 -1508
rect 3595 -1526 3657 -1510
rect 3701 -1515 3717 -1508
rect 3779 -1515 3809 -1504
rect 3857 -1508 3903 -1492
rect 3930 -1504 4004 -1488
rect 3857 -1510 3891 -1508
rect 3856 -1526 3903 -1510
rect 3930 -1526 3943 -1504
rect 3958 -1526 3988 -1504
rect 4015 -1526 4016 -1510
rect 4031 -1526 4044 -1366
rect 4074 -1470 4087 -1366
rect 4132 -1388 4133 -1378
rect 4148 -1388 4161 -1378
rect 4132 -1392 4161 -1388
rect 4166 -1392 4196 -1366
rect 4214 -1380 4230 -1378
rect 4302 -1380 4355 -1366
rect 4303 -1382 4367 -1380
rect 4410 -1382 4425 -1366
rect 4474 -1369 4504 -1366
rect 4611 -1367 6944 -1366
rect 4474 -1372 4510 -1369
rect 4440 -1380 4456 -1378
rect 4214 -1392 4229 -1388
rect 4132 -1394 4229 -1392
rect 4257 -1394 4425 -1382
rect 4441 -1392 4456 -1388
rect 4474 -1391 4513 -1372
rect 4532 -1378 4539 -1377
rect 4538 -1385 4539 -1378
rect 4522 -1388 4523 -1385
rect 4538 -1388 4551 -1385
rect 4474 -1392 4504 -1391
rect 4513 -1392 4519 -1391
rect 4522 -1392 4551 -1388
rect 4441 -1393 4551 -1392
rect 4441 -1394 4557 -1393
rect 4116 -1402 4167 -1394
rect 4116 -1414 4141 -1402
rect 4148 -1414 4167 -1402
rect 4198 -1402 4248 -1394
rect 4198 -1410 4214 -1402
rect 4221 -1404 4248 -1402
rect 4257 -1404 4478 -1394
rect 4221 -1414 4478 -1404
rect 4507 -1402 4557 -1394
rect 4507 -1411 4523 -1402
rect 4116 -1422 4167 -1414
rect 4214 -1422 4478 -1414
rect 4504 -1414 4523 -1411
rect 4530 -1414 4557 -1402
rect 4504 -1422 4557 -1414
rect 4132 -1430 4133 -1422
rect 4148 -1430 4161 -1422
rect 4132 -1438 4148 -1430
rect 4129 -1445 4148 -1442
rect 4129 -1454 4151 -1445
rect 4102 -1464 4151 -1454
rect 4102 -1470 4132 -1464
rect 4151 -1469 4156 -1464
rect 4074 -1486 4148 -1470
rect 4166 -1478 4196 -1422
rect 4231 -1432 4439 -1422
rect 4474 -1426 4519 -1422
rect 4522 -1423 4523 -1422
rect 4538 -1423 4551 -1422
rect 4257 -1462 4446 -1432
rect 4272 -1465 4446 -1462
rect 4265 -1468 4446 -1465
rect 4074 -1488 4087 -1486
rect 4102 -1488 4136 -1486
rect 4074 -1504 4148 -1488
rect 4175 -1492 4188 -1478
rect 4203 -1492 4219 -1476
rect 4265 -1481 4276 -1468
rect 4058 -1526 4059 -1510
rect 4074 -1526 4087 -1504
rect 4102 -1526 4132 -1504
rect 4175 -1508 4237 -1492
rect 4265 -1499 4276 -1483
rect 4281 -1488 4291 -1468
rect 4301 -1488 4315 -1468
rect 4318 -1481 4327 -1468
rect 4343 -1481 4352 -1468
rect 4281 -1499 4315 -1488
rect 4318 -1499 4327 -1483
rect 4343 -1499 4352 -1483
rect 4359 -1488 4369 -1468
rect 4379 -1488 4393 -1468
rect 4394 -1481 4405 -1468
rect 4359 -1499 4393 -1488
rect 4394 -1499 4405 -1483
rect 4451 -1492 4467 -1476
rect 4474 -1478 4504 -1426
rect 4538 -1430 4539 -1423
rect 4523 -1438 4539 -1430
rect 4510 -1470 4523 -1451
rect 4538 -1470 4568 -1454
rect 4510 -1486 4584 -1470
rect 4510 -1488 4523 -1486
rect 4538 -1488 4572 -1486
rect 4175 -1510 4188 -1508
rect 4203 -1510 4237 -1508
rect 4175 -1526 4237 -1510
rect 4281 -1515 4297 -1508
rect 4359 -1515 4389 -1504
rect 4437 -1508 4483 -1492
rect 4510 -1504 4584 -1488
rect 4437 -1510 4471 -1508
rect 4436 -1526 4483 -1510
rect 4510 -1526 4523 -1504
rect 4538 -1526 4568 -1504
rect 4595 -1526 4596 -1510
rect 4611 -1526 4624 -1367
rect 4654 -1471 4667 -1367
rect 4712 -1389 4713 -1379
rect 4728 -1389 4741 -1379
rect 4712 -1393 4741 -1389
rect 4746 -1393 4776 -1367
rect 4794 -1381 4810 -1379
rect 4882 -1381 4935 -1367
rect 4883 -1383 4947 -1381
rect 4990 -1383 5005 -1367
rect 5054 -1370 5084 -1367
rect 5054 -1373 5090 -1370
rect 5020 -1381 5036 -1379
rect 4794 -1393 4809 -1389
rect 4712 -1395 4809 -1393
rect 4837 -1395 5005 -1383
rect 5021 -1393 5036 -1389
rect 5054 -1392 5093 -1373
rect 5112 -1379 5119 -1378
rect 5118 -1386 5119 -1379
rect 5102 -1389 5103 -1386
rect 5118 -1389 5131 -1386
rect 5054 -1393 5084 -1392
rect 5093 -1393 5099 -1392
rect 5102 -1393 5131 -1389
rect 5021 -1394 5131 -1393
rect 5021 -1395 5137 -1394
rect 4696 -1403 4747 -1395
rect 4696 -1415 4721 -1403
rect 4728 -1415 4747 -1403
rect 4778 -1403 4828 -1395
rect 4778 -1411 4794 -1403
rect 4801 -1405 4828 -1403
rect 4837 -1405 5058 -1395
rect 4801 -1415 5058 -1405
rect 5087 -1403 5137 -1395
rect 5087 -1412 5103 -1403
rect 4696 -1423 4747 -1415
rect 4794 -1423 5058 -1415
rect 5084 -1415 5103 -1412
rect 5110 -1415 5137 -1403
rect 5084 -1423 5137 -1415
rect 4712 -1431 4713 -1423
rect 4728 -1431 4741 -1423
rect 4712 -1439 4728 -1431
rect 4709 -1446 4728 -1443
rect 4709 -1455 4731 -1446
rect 4682 -1465 4731 -1455
rect 4682 -1471 4712 -1465
rect 4731 -1470 4736 -1465
rect 4654 -1487 4728 -1471
rect 4746 -1479 4776 -1423
rect 4811 -1433 5019 -1423
rect 5054 -1427 5099 -1423
rect 5102 -1424 5103 -1423
rect 5118 -1424 5131 -1423
rect 4837 -1463 5026 -1433
rect 4852 -1466 5026 -1463
rect 4845 -1469 5026 -1466
rect 4654 -1489 4667 -1487
rect 4682 -1489 4716 -1487
rect 4654 -1505 4728 -1489
rect 4755 -1493 4768 -1479
rect 4783 -1493 4799 -1477
rect 4845 -1482 4856 -1469
rect 3435 -1534 3470 -1526
rect 3435 -1560 3436 -1534
rect 3443 -1560 3470 -1534
rect 3379 -1578 3408 -1564
rect 3435 -1568 3470 -1560
rect 3472 -1534 3513 -1526
rect 3472 -1560 3487 -1534
rect 3494 -1560 3513 -1534
rect 3577 -1538 3639 -1526
rect 3651 -1538 3726 -1526
rect 3784 -1538 3859 -1526
rect 3871 -1538 3902 -1526
rect 3908 -1538 3943 -1526
rect 3577 -1540 3739 -1538
rect 3472 -1568 3513 -1560
rect 3595 -1564 3608 -1540
rect 3623 -1542 3638 -1540
rect 3435 -1578 3436 -1568
rect 3451 -1578 3464 -1568
rect 3478 -1578 3479 -1568
rect 3494 -1578 3507 -1568
rect 3522 -1578 3552 -1564
rect 3595 -1578 3638 -1564
rect 3662 -1567 3669 -1560
rect 3672 -1564 3739 -1540
rect 3771 -1540 3943 -1538
rect 3741 -1562 3769 -1558
rect 3771 -1562 3851 -1540
rect 3872 -1542 3887 -1540
rect 3741 -1564 3851 -1562
rect 3672 -1568 3851 -1564
rect 3645 -1578 3675 -1568
rect 3677 -1578 3830 -1568
rect 3838 -1578 3868 -1568
rect 3872 -1578 3902 -1564
rect 3930 -1578 3943 -1540
rect 4015 -1534 4050 -1526
rect 4015 -1560 4016 -1534
rect 4023 -1560 4050 -1534
rect 3958 -1578 3988 -1564
rect 4015 -1568 4050 -1560
rect 4052 -1534 4093 -1526
rect 4052 -1560 4067 -1534
rect 4074 -1560 4093 -1534
rect 4157 -1538 4219 -1526
rect 4231 -1538 4306 -1526
rect 4364 -1538 4439 -1526
rect 4451 -1538 4482 -1526
rect 4488 -1538 4523 -1526
rect 4157 -1540 4319 -1538
rect 4052 -1568 4093 -1560
rect 4175 -1564 4188 -1540
rect 4203 -1542 4218 -1540
rect 4015 -1578 4016 -1568
rect 4031 -1578 4044 -1568
rect 4058 -1578 4059 -1568
rect 4074 -1578 4087 -1568
rect 4102 -1578 4132 -1564
rect 4175 -1578 4218 -1564
rect 4242 -1567 4249 -1560
rect 4252 -1564 4319 -1540
rect 4351 -1540 4523 -1538
rect 4321 -1562 4349 -1558
rect 4351 -1562 4431 -1540
rect 4452 -1542 4467 -1540
rect 4321 -1564 4431 -1562
rect 4252 -1568 4431 -1564
rect 4225 -1578 4255 -1568
rect 4257 -1578 4410 -1568
rect 4418 -1578 4448 -1568
rect 4452 -1578 4482 -1564
rect 4510 -1578 4523 -1540
rect 4595 -1534 4630 -1526
rect 4638 -1527 4639 -1511
rect 4654 -1527 4667 -1505
rect 4682 -1527 4712 -1505
rect 4755 -1509 4817 -1493
rect 4845 -1500 4856 -1484
rect 4861 -1489 4871 -1469
rect 4881 -1489 4895 -1469
rect 4898 -1482 4907 -1469
rect 4923 -1482 4932 -1469
rect 4861 -1500 4895 -1489
rect 4898 -1500 4907 -1484
rect 4923 -1500 4932 -1484
rect 4939 -1489 4949 -1469
rect 4959 -1489 4973 -1469
rect 4974 -1482 4985 -1469
rect 4939 -1500 4973 -1489
rect 4974 -1500 4985 -1484
rect 5031 -1493 5047 -1477
rect 5054 -1479 5084 -1427
rect 5118 -1431 5119 -1424
rect 5103 -1439 5119 -1431
rect 5090 -1471 5103 -1452
rect 5118 -1471 5148 -1455
rect 5090 -1487 5164 -1471
rect 5090 -1489 5103 -1487
rect 5118 -1489 5152 -1487
rect 4755 -1511 4768 -1509
rect 4783 -1511 4817 -1509
rect 4755 -1527 4817 -1511
rect 4861 -1516 4877 -1509
rect 4939 -1516 4969 -1505
rect 5017 -1509 5063 -1493
rect 5090 -1505 5164 -1489
rect 5017 -1511 5051 -1509
rect 5016 -1527 5063 -1511
rect 5090 -1527 5103 -1505
rect 5118 -1527 5148 -1505
rect 5175 -1527 5176 -1511
rect 5191 -1527 5204 -1367
rect 5234 -1471 5247 -1367
rect 5292 -1389 5293 -1379
rect 5308 -1389 5321 -1379
rect 5292 -1393 5321 -1389
rect 5326 -1393 5356 -1367
rect 5374 -1381 5390 -1379
rect 5462 -1381 5515 -1367
rect 5463 -1383 5527 -1381
rect 5570 -1383 5585 -1367
rect 5634 -1370 5664 -1367
rect 5634 -1373 5670 -1370
rect 5600 -1381 5616 -1379
rect 5374 -1393 5389 -1389
rect 5292 -1395 5389 -1393
rect 5417 -1395 5585 -1383
rect 5601 -1393 5616 -1389
rect 5634 -1392 5673 -1373
rect 5692 -1379 5699 -1378
rect 5698 -1386 5699 -1379
rect 5682 -1389 5683 -1386
rect 5698 -1389 5711 -1386
rect 5634 -1393 5664 -1392
rect 5673 -1393 5679 -1392
rect 5682 -1393 5711 -1389
rect 5601 -1394 5711 -1393
rect 5601 -1395 5717 -1394
rect 5276 -1403 5327 -1395
rect 5276 -1415 5301 -1403
rect 5308 -1415 5327 -1403
rect 5358 -1403 5408 -1395
rect 5358 -1411 5374 -1403
rect 5381 -1405 5408 -1403
rect 5417 -1405 5638 -1395
rect 5381 -1415 5638 -1405
rect 5667 -1403 5717 -1395
rect 5667 -1412 5683 -1403
rect 5276 -1423 5327 -1415
rect 5374 -1423 5638 -1415
rect 5664 -1415 5683 -1412
rect 5690 -1415 5717 -1403
rect 5664 -1423 5717 -1415
rect 5292 -1431 5293 -1423
rect 5308 -1431 5321 -1423
rect 5292 -1439 5308 -1431
rect 5289 -1446 5308 -1443
rect 5289 -1455 5311 -1446
rect 5262 -1465 5311 -1455
rect 5262 -1471 5292 -1465
rect 5311 -1470 5316 -1465
rect 5234 -1487 5308 -1471
rect 5326 -1479 5356 -1423
rect 5391 -1433 5599 -1423
rect 5634 -1427 5679 -1423
rect 5682 -1424 5683 -1423
rect 5698 -1424 5711 -1423
rect 5417 -1463 5606 -1433
rect 5432 -1466 5606 -1463
rect 5425 -1469 5606 -1466
rect 5234 -1489 5247 -1487
rect 5262 -1489 5296 -1487
rect 5234 -1505 5308 -1489
rect 5335 -1493 5348 -1479
rect 5363 -1493 5379 -1477
rect 5425 -1482 5436 -1469
rect 5218 -1527 5219 -1511
rect 5234 -1527 5247 -1505
rect 5262 -1527 5292 -1505
rect 5335 -1509 5397 -1493
rect 5425 -1500 5436 -1484
rect 5441 -1489 5451 -1469
rect 5461 -1489 5475 -1469
rect 5478 -1482 5487 -1469
rect 5503 -1482 5512 -1469
rect 5441 -1500 5475 -1489
rect 5478 -1500 5487 -1484
rect 5503 -1500 5512 -1484
rect 5519 -1489 5529 -1469
rect 5539 -1489 5553 -1469
rect 5554 -1482 5565 -1469
rect 5519 -1500 5553 -1489
rect 5554 -1500 5565 -1484
rect 5611 -1493 5627 -1477
rect 5634 -1479 5664 -1427
rect 5698 -1431 5699 -1424
rect 5683 -1439 5699 -1431
rect 5670 -1471 5683 -1452
rect 5698 -1471 5728 -1455
rect 5670 -1487 5744 -1471
rect 5670 -1489 5683 -1487
rect 5698 -1489 5732 -1487
rect 5335 -1511 5348 -1509
rect 5363 -1511 5397 -1509
rect 5335 -1527 5397 -1511
rect 5441 -1516 5457 -1509
rect 5519 -1516 5549 -1505
rect 5597 -1509 5643 -1493
rect 5670 -1505 5744 -1489
rect 5597 -1511 5631 -1509
rect 5596 -1527 5643 -1511
rect 5670 -1527 5683 -1505
rect 5698 -1527 5728 -1505
rect 5755 -1527 5756 -1511
rect 5771 -1527 5784 -1367
rect 5814 -1471 5827 -1367
rect 5872 -1389 5873 -1379
rect 5888 -1389 5901 -1379
rect 5872 -1393 5901 -1389
rect 5906 -1393 5936 -1367
rect 5954 -1381 5970 -1379
rect 6042 -1381 6095 -1367
rect 6043 -1383 6107 -1381
rect 6150 -1383 6165 -1367
rect 6214 -1370 6244 -1367
rect 6214 -1373 6250 -1370
rect 6180 -1381 6196 -1379
rect 5954 -1393 5969 -1389
rect 5872 -1395 5969 -1393
rect 5997 -1395 6165 -1383
rect 6181 -1393 6196 -1389
rect 6214 -1392 6253 -1373
rect 6272 -1379 6279 -1378
rect 6278 -1386 6279 -1379
rect 6262 -1389 6263 -1386
rect 6278 -1389 6291 -1386
rect 6214 -1393 6244 -1392
rect 6253 -1393 6259 -1392
rect 6262 -1393 6291 -1389
rect 6181 -1394 6291 -1393
rect 6181 -1395 6297 -1394
rect 5856 -1403 5907 -1395
rect 5856 -1415 5881 -1403
rect 5888 -1415 5907 -1403
rect 5938 -1403 5988 -1395
rect 5938 -1411 5954 -1403
rect 5961 -1405 5988 -1403
rect 5997 -1405 6218 -1395
rect 5961 -1415 6218 -1405
rect 6247 -1403 6297 -1395
rect 6247 -1412 6263 -1403
rect 5856 -1423 5907 -1415
rect 5954 -1423 6218 -1415
rect 6244 -1415 6263 -1412
rect 6270 -1415 6297 -1403
rect 6244 -1423 6297 -1415
rect 5872 -1431 5873 -1423
rect 5888 -1431 5901 -1423
rect 5872 -1439 5888 -1431
rect 5869 -1446 5888 -1443
rect 5869 -1455 5891 -1446
rect 5842 -1465 5891 -1455
rect 5842 -1471 5872 -1465
rect 5891 -1470 5896 -1465
rect 5814 -1487 5888 -1471
rect 5906 -1479 5936 -1423
rect 5971 -1433 6179 -1423
rect 6214 -1427 6259 -1423
rect 6262 -1424 6263 -1423
rect 6278 -1424 6291 -1423
rect 5997 -1463 6186 -1433
rect 6012 -1466 6186 -1463
rect 6005 -1469 6186 -1466
rect 5814 -1489 5827 -1487
rect 5842 -1489 5876 -1487
rect 5814 -1505 5888 -1489
rect 5915 -1493 5928 -1479
rect 5943 -1493 5959 -1477
rect 6005 -1482 6016 -1469
rect 5798 -1527 5799 -1511
rect 5814 -1527 5827 -1505
rect 5842 -1527 5872 -1505
rect 5915 -1509 5977 -1493
rect 6005 -1500 6016 -1484
rect 6021 -1489 6031 -1469
rect 6041 -1489 6055 -1469
rect 6058 -1482 6067 -1469
rect 6083 -1482 6092 -1469
rect 6021 -1500 6055 -1489
rect 6058 -1500 6067 -1484
rect 6083 -1500 6092 -1484
rect 6099 -1489 6109 -1469
rect 6119 -1489 6133 -1469
rect 6134 -1482 6145 -1469
rect 6099 -1500 6133 -1489
rect 6134 -1500 6145 -1484
rect 6191 -1493 6207 -1477
rect 6214 -1479 6244 -1427
rect 6278 -1431 6279 -1424
rect 6263 -1439 6279 -1431
rect 6250 -1471 6263 -1452
rect 6278 -1471 6308 -1455
rect 6250 -1487 6324 -1471
rect 6250 -1489 6263 -1487
rect 6278 -1489 6312 -1487
rect 5915 -1511 5928 -1509
rect 5943 -1511 5977 -1509
rect 5915 -1527 5977 -1511
rect 6021 -1516 6037 -1509
rect 6099 -1516 6129 -1505
rect 6177 -1509 6223 -1493
rect 6250 -1505 6324 -1489
rect 6177 -1511 6211 -1509
rect 6176 -1527 6223 -1511
rect 6250 -1527 6263 -1505
rect 6278 -1527 6308 -1505
rect 6335 -1527 6336 -1511
rect 6351 -1527 6364 -1367
rect 6394 -1471 6407 -1367
rect 6452 -1389 6453 -1379
rect 6468 -1389 6481 -1379
rect 6452 -1393 6481 -1389
rect 6486 -1393 6516 -1367
rect 6534 -1381 6550 -1379
rect 6622 -1381 6675 -1367
rect 6623 -1383 6687 -1381
rect 6730 -1383 6745 -1367
rect 6794 -1370 6824 -1367
rect 6794 -1373 6830 -1370
rect 6760 -1381 6776 -1379
rect 6534 -1393 6549 -1389
rect 6452 -1395 6549 -1393
rect 6577 -1395 6745 -1383
rect 6761 -1393 6776 -1389
rect 6794 -1392 6833 -1373
rect 6852 -1379 6859 -1378
rect 6858 -1386 6859 -1379
rect 6842 -1389 6843 -1386
rect 6858 -1389 6871 -1386
rect 6794 -1393 6824 -1392
rect 6833 -1393 6839 -1392
rect 6842 -1393 6871 -1389
rect 6761 -1394 6871 -1393
rect 6761 -1395 6877 -1394
rect 6436 -1403 6487 -1395
rect 6436 -1415 6461 -1403
rect 6468 -1415 6487 -1403
rect 6518 -1403 6568 -1395
rect 6518 -1411 6534 -1403
rect 6541 -1405 6568 -1403
rect 6577 -1405 6798 -1395
rect 6541 -1415 6798 -1405
rect 6827 -1403 6877 -1395
rect 6827 -1412 6843 -1403
rect 6436 -1423 6487 -1415
rect 6534 -1423 6798 -1415
rect 6824 -1415 6843 -1412
rect 6850 -1415 6877 -1403
rect 6824 -1423 6877 -1415
rect 6452 -1431 6453 -1423
rect 6468 -1431 6481 -1423
rect 6452 -1439 6468 -1431
rect 6449 -1446 6468 -1443
rect 6449 -1455 6471 -1446
rect 6422 -1465 6471 -1455
rect 6422 -1471 6452 -1465
rect 6471 -1470 6476 -1465
rect 6394 -1487 6468 -1471
rect 6486 -1479 6516 -1423
rect 6551 -1433 6759 -1423
rect 6794 -1427 6839 -1423
rect 6842 -1424 6843 -1423
rect 6858 -1424 6871 -1423
rect 6577 -1463 6766 -1433
rect 6592 -1466 6766 -1463
rect 6585 -1469 6766 -1466
rect 6394 -1489 6407 -1487
rect 6422 -1489 6456 -1487
rect 6394 -1505 6468 -1489
rect 6495 -1493 6508 -1479
rect 6523 -1493 6539 -1477
rect 6585 -1482 6596 -1469
rect 6378 -1527 6379 -1511
rect 6394 -1527 6407 -1505
rect 6422 -1527 6452 -1505
rect 6495 -1509 6557 -1493
rect 6585 -1500 6596 -1484
rect 6601 -1489 6611 -1469
rect 6621 -1489 6635 -1469
rect 6638 -1482 6647 -1469
rect 6663 -1482 6672 -1469
rect 6601 -1500 6635 -1489
rect 6638 -1500 6647 -1484
rect 6663 -1500 6672 -1484
rect 6679 -1489 6689 -1469
rect 6699 -1489 6713 -1469
rect 6714 -1482 6725 -1469
rect 6679 -1500 6713 -1489
rect 6714 -1500 6725 -1484
rect 6771 -1493 6787 -1477
rect 6794 -1479 6824 -1427
rect 6858 -1431 6859 -1424
rect 6843 -1439 6859 -1431
rect 6830 -1471 6843 -1452
rect 6858 -1471 6888 -1455
rect 6830 -1487 6904 -1471
rect 6830 -1489 6843 -1487
rect 6858 -1489 6892 -1487
rect 6495 -1511 6508 -1509
rect 6523 -1511 6557 -1509
rect 6495 -1527 6557 -1511
rect 6601 -1516 6617 -1509
rect 6679 -1516 6709 -1505
rect 6757 -1509 6803 -1493
rect 6830 -1505 6904 -1489
rect 6757 -1511 6791 -1509
rect 6756 -1527 6803 -1511
rect 6830 -1527 6843 -1505
rect 6858 -1527 6888 -1505
rect 6915 -1527 6916 -1511
rect 6931 -1527 6944 -1367
rect 4595 -1560 4596 -1534
rect 4603 -1560 4630 -1534
rect 4538 -1578 4568 -1564
rect 4595 -1568 4630 -1560
rect 4632 -1535 4673 -1527
rect 4632 -1561 4647 -1535
rect 4654 -1561 4673 -1535
rect 4737 -1539 4799 -1527
rect 4811 -1539 4886 -1527
rect 4944 -1539 5019 -1527
rect 5031 -1539 5062 -1527
rect 5068 -1539 5103 -1527
rect 4737 -1541 4899 -1539
rect 4755 -1559 4768 -1541
rect 4783 -1543 4798 -1541
rect 4595 -1578 4596 -1568
rect 4611 -1578 4624 -1568
rect 4632 -1569 4673 -1561
rect 4756 -1565 4768 -1559
rect 3379 -1579 4624 -1578
rect 4638 -1579 4639 -1569
rect 4654 -1579 4667 -1569
rect 4682 -1579 4712 -1565
rect 4756 -1579 4798 -1565
rect 4822 -1568 4829 -1561
rect 4832 -1565 4899 -1541
rect 4931 -1541 5103 -1539
rect 4901 -1563 4929 -1559
rect 4931 -1563 5011 -1541
rect 5032 -1543 5047 -1541
rect 4901 -1565 5011 -1563
rect 4832 -1569 5011 -1565
rect 4805 -1579 4835 -1569
rect 4837 -1579 4990 -1569
rect 4998 -1579 5028 -1569
rect 5032 -1579 5062 -1565
rect 5090 -1579 5103 -1541
rect 5175 -1535 5210 -1527
rect 5175 -1561 5176 -1535
rect 5183 -1561 5210 -1535
rect 5118 -1579 5148 -1565
rect 5175 -1569 5210 -1561
rect 5212 -1535 5253 -1527
rect 5212 -1561 5227 -1535
rect 5234 -1561 5253 -1535
rect 5317 -1539 5379 -1527
rect 5391 -1539 5466 -1527
rect 5524 -1539 5599 -1527
rect 5611 -1539 5642 -1527
rect 5648 -1539 5683 -1527
rect 5317 -1541 5479 -1539
rect 5335 -1559 5348 -1541
rect 5363 -1543 5378 -1541
rect 5212 -1569 5253 -1561
rect 5336 -1565 5348 -1559
rect 5175 -1579 5176 -1569
rect 5191 -1579 5204 -1569
rect 5218 -1579 5219 -1569
rect 5234 -1579 5247 -1569
rect 5262 -1579 5292 -1565
rect 5336 -1579 5378 -1565
rect 5402 -1568 5409 -1561
rect 5412 -1565 5479 -1541
rect 5511 -1541 5683 -1539
rect 5481 -1563 5509 -1559
rect 5511 -1563 5591 -1541
rect 5612 -1543 5627 -1541
rect 5481 -1565 5591 -1563
rect 5412 -1569 5591 -1565
rect 5385 -1579 5415 -1569
rect 5417 -1579 5570 -1569
rect 5578 -1579 5608 -1569
rect 5612 -1579 5642 -1565
rect 5670 -1579 5683 -1541
rect 5755 -1535 5790 -1527
rect 5755 -1561 5756 -1535
rect 5763 -1561 5790 -1535
rect 5698 -1579 5728 -1565
rect 5755 -1569 5790 -1561
rect 5792 -1535 5833 -1527
rect 5792 -1561 5807 -1535
rect 5814 -1561 5833 -1535
rect 5897 -1539 5959 -1527
rect 5971 -1539 6046 -1527
rect 6104 -1539 6179 -1527
rect 6191 -1539 6222 -1527
rect 6228 -1539 6263 -1527
rect 5897 -1541 6059 -1539
rect 5915 -1559 5928 -1541
rect 5943 -1543 5958 -1541
rect 5792 -1569 5833 -1561
rect 5916 -1565 5928 -1559
rect 5755 -1579 5756 -1569
rect 5771 -1579 5784 -1569
rect 5798 -1579 5799 -1569
rect 5814 -1579 5827 -1569
rect 5842 -1579 5872 -1565
rect 5916 -1579 5958 -1565
rect 5982 -1568 5989 -1561
rect 5992 -1565 6059 -1541
rect 6091 -1541 6263 -1539
rect 6061 -1563 6089 -1559
rect 6091 -1563 6171 -1541
rect 6192 -1543 6207 -1541
rect 6061 -1565 6171 -1563
rect 5992 -1569 6171 -1565
rect 5965 -1579 5995 -1569
rect 5997 -1579 6150 -1569
rect 6158 -1579 6188 -1569
rect 6192 -1579 6222 -1565
rect 6250 -1579 6263 -1541
rect 6335 -1535 6370 -1527
rect 6335 -1561 6336 -1535
rect 6343 -1561 6370 -1535
rect 6278 -1579 6308 -1565
rect 6335 -1569 6370 -1561
rect 6372 -1535 6413 -1527
rect 6372 -1561 6387 -1535
rect 6394 -1561 6413 -1535
rect 6477 -1539 6539 -1527
rect 6551 -1539 6626 -1527
rect 6684 -1539 6759 -1527
rect 6771 -1539 6802 -1527
rect 6808 -1539 6843 -1527
rect 6477 -1541 6639 -1539
rect 6495 -1559 6508 -1541
rect 6523 -1543 6538 -1541
rect 6372 -1569 6413 -1561
rect 6496 -1565 6508 -1559
rect 6335 -1579 6336 -1569
rect 6351 -1579 6364 -1569
rect 6378 -1579 6379 -1569
rect 6394 -1579 6407 -1569
rect 6422 -1579 6452 -1565
rect 6496 -1579 6538 -1565
rect 6562 -1568 6569 -1561
rect 6572 -1565 6639 -1541
rect 6671 -1541 6843 -1539
rect 6641 -1563 6669 -1559
rect 6671 -1563 6751 -1541
rect 6772 -1543 6787 -1541
rect 6641 -1565 6751 -1563
rect 6572 -1569 6751 -1565
rect 6545 -1579 6575 -1569
rect 6577 -1579 6730 -1569
rect 6738 -1579 6768 -1569
rect 6772 -1579 6802 -1565
rect 6830 -1579 6843 -1541
rect 6915 -1535 6950 -1527
rect 6915 -1561 6916 -1535
rect 6923 -1561 6950 -1535
rect 6858 -1579 6888 -1565
rect 6915 -1569 6950 -1561
rect 6915 -1579 6916 -1569
rect 6931 -1579 6944 -1569
rect 3379 -1592 6944 -1579
rect 3379 -1610 3408 -1592
rect 3451 -1622 3464 -1592
rect 3494 -1622 3507 -1592
rect 3522 -1610 3552 -1592
rect 3595 -1606 3609 -1592
rect 3645 -1606 3865 -1592
rect 3596 -1608 3609 -1606
rect 3562 -1620 3577 -1608
rect 3559 -1622 3581 -1620
rect 3586 -1622 3616 -1608
rect 3677 -1610 3830 -1606
rect 3659 -1622 3851 -1610
rect 3894 -1622 3924 -1608
rect 3930 -1622 3943 -1592
rect 3958 -1610 3988 -1592
rect 4031 -1622 4044 -1592
rect 4074 -1622 4087 -1592
rect 4102 -1610 4132 -1592
rect 4175 -1606 4189 -1592
rect 4225 -1606 4445 -1592
rect 4176 -1608 4189 -1606
rect 4142 -1620 4157 -1608
rect 4139 -1622 4161 -1620
rect 4166 -1622 4196 -1608
rect 4257 -1610 4410 -1606
rect 4239 -1622 4431 -1610
rect 4474 -1622 4504 -1608
rect 4510 -1622 4523 -1592
rect 4538 -1610 4568 -1592
rect 4611 -1593 6944 -1592
rect 4611 -1622 4624 -1593
rect 3379 -1623 4624 -1622
rect 4654 -1623 4667 -1593
rect 4682 -1611 4712 -1593
rect 4756 -1609 4769 -1593
rect 4805 -1607 5025 -1593
rect 4722 -1621 4737 -1609
rect 4719 -1623 4741 -1621
rect 4746 -1623 4776 -1609
rect 4837 -1611 4990 -1607
rect 4819 -1623 5011 -1611
rect 5054 -1623 5084 -1609
rect 5090 -1623 5103 -1593
rect 5118 -1611 5148 -1593
rect 5191 -1623 5204 -1593
rect 5234 -1623 5247 -1593
rect 5262 -1611 5292 -1593
rect 5336 -1609 5349 -1593
rect 5385 -1607 5605 -1593
rect 5302 -1621 5317 -1609
rect 5299 -1623 5321 -1621
rect 5326 -1623 5356 -1609
rect 5417 -1611 5570 -1607
rect 5399 -1623 5591 -1611
rect 5634 -1623 5664 -1609
rect 5670 -1623 5683 -1593
rect 5698 -1611 5728 -1593
rect 5771 -1623 5784 -1593
rect 5814 -1623 5827 -1593
rect 5842 -1611 5872 -1593
rect 5916 -1609 5929 -1593
rect 5965 -1607 6185 -1593
rect 5882 -1621 5897 -1609
rect 5879 -1623 5901 -1621
rect 5906 -1623 5936 -1609
rect 5997 -1611 6150 -1607
rect 5979 -1623 6171 -1611
rect 6214 -1623 6244 -1609
rect 6250 -1623 6263 -1593
rect 6278 -1611 6308 -1593
rect 6351 -1623 6364 -1593
rect 6394 -1623 6407 -1593
rect 6422 -1611 6452 -1593
rect 6496 -1609 6509 -1593
rect 6545 -1607 6765 -1593
rect 6462 -1621 6477 -1609
rect 6459 -1623 6481 -1621
rect 6486 -1623 6516 -1609
rect 6577 -1611 6730 -1607
rect 6559 -1623 6751 -1611
rect 6794 -1623 6824 -1609
rect 6830 -1623 6843 -1593
rect 6858 -1611 6888 -1593
rect 6931 -1623 6944 -1593
rect 3379 -1636 6944 -1623
rect 3379 -1663 3391 -1655
rect 3379 -1692 3397 -1663
rect 3379 -1693 3391 -1692
rect 3379 -1740 3408 -1724
rect 3379 -1756 3424 -1740
rect 3379 -1758 3412 -1756
rect 3379 -1774 3424 -1758
rect 3379 -1796 3408 -1774
rect 3435 -1796 3436 -1780
rect 3451 -1796 3464 -1636
rect 3494 -1740 3507 -1636
rect 3552 -1658 3553 -1648
rect 3568 -1658 3581 -1648
rect 3552 -1662 3581 -1658
rect 3586 -1662 3616 -1636
rect 3634 -1650 3650 -1648
rect 3722 -1650 3775 -1636
rect 3723 -1652 3787 -1650
rect 3830 -1652 3845 -1636
rect 3894 -1639 3924 -1636
rect 3894 -1642 3930 -1639
rect 3860 -1650 3876 -1648
rect 3634 -1662 3649 -1658
rect 3552 -1664 3649 -1662
rect 3677 -1664 3845 -1652
rect 3861 -1662 3876 -1658
rect 3894 -1661 3933 -1642
rect 3952 -1648 3959 -1647
rect 3958 -1655 3959 -1648
rect 3942 -1658 3943 -1655
rect 3958 -1658 3971 -1655
rect 3894 -1662 3924 -1661
rect 3933 -1662 3939 -1661
rect 3942 -1662 3971 -1658
rect 3861 -1663 3971 -1662
rect 3861 -1664 3977 -1663
rect 3536 -1672 3587 -1664
rect 3536 -1684 3561 -1672
rect 3568 -1684 3587 -1672
rect 3618 -1672 3668 -1664
rect 3618 -1680 3634 -1672
rect 3641 -1674 3668 -1672
rect 3677 -1674 3898 -1664
rect 3641 -1684 3898 -1674
rect 3927 -1672 3977 -1664
rect 3927 -1681 3943 -1672
rect 3536 -1692 3587 -1684
rect 3634 -1692 3898 -1684
rect 3924 -1684 3943 -1681
rect 3950 -1684 3977 -1672
rect 3924 -1692 3977 -1684
rect 3552 -1700 3553 -1692
rect 3568 -1700 3581 -1692
rect 3552 -1708 3568 -1700
rect 3549 -1715 3568 -1712
rect 3549 -1724 3571 -1715
rect 3522 -1734 3571 -1724
rect 3522 -1740 3552 -1734
rect 3571 -1739 3576 -1734
rect 3494 -1756 3568 -1740
rect 3586 -1748 3616 -1692
rect 3651 -1702 3859 -1692
rect 3894 -1696 3939 -1692
rect 3942 -1693 3943 -1692
rect 3958 -1693 3971 -1692
rect 3677 -1732 3866 -1702
rect 3692 -1735 3866 -1732
rect 3685 -1738 3866 -1735
rect 3494 -1758 3507 -1756
rect 3522 -1758 3556 -1756
rect 3494 -1774 3568 -1758
rect 3595 -1762 3608 -1748
rect 3623 -1762 3639 -1746
rect 3685 -1751 3696 -1738
rect 3478 -1796 3479 -1780
rect 3494 -1796 3507 -1774
rect 3522 -1796 3552 -1774
rect 3595 -1778 3657 -1762
rect 3685 -1769 3696 -1753
rect 3701 -1758 3711 -1738
rect 3721 -1758 3735 -1738
rect 3738 -1751 3747 -1738
rect 3763 -1751 3772 -1738
rect 3701 -1769 3735 -1758
rect 3738 -1769 3747 -1753
rect 3763 -1769 3772 -1753
rect 3779 -1758 3789 -1738
rect 3799 -1758 3813 -1738
rect 3814 -1751 3825 -1738
rect 3779 -1769 3813 -1758
rect 3814 -1769 3825 -1753
rect 3871 -1762 3887 -1746
rect 3894 -1748 3924 -1696
rect 3958 -1700 3959 -1693
rect 3943 -1708 3959 -1700
rect 3930 -1740 3943 -1721
rect 3958 -1740 3988 -1724
rect 3930 -1756 4004 -1740
rect 3930 -1758 3943 -1756
rect 3958 -1758 3992 -1756
rect 3595 -1780 3608 -1778
rect 3623 -1780 3657 -1778
rect 3595 -1796 3657 -1780
rect 3701 -1785 3717 -1778
rect 3779 -1785 3809 -1774
rect 3857 -1778 3903 -1762
rect 3930 -1774 4004 -1758
rect 3857 -1780 3891 -1778
rect 3856 -1796 3903 -1780
rect 3930 -1796 3943 -1774
rect 3958 -1796 3988 -1774
rect 4015 -1796 4016 -1780
rect 4031 -1796 4044 -1636
rect 4074 -1740 4087 -1636
rect 4132 -1658 4133 -1648
rect 4148 -1658 4161 -1648
rect 4132 -1662 4161 -1658
rect 4166 -1662 4196 -1636
rect 4214 -1650 4230 -1648
rect 4302 -1650 4355 -1636
rect 4303 -1652 4367 -1650
rect 4410 -1652 4425 -1636
rect 4474 -1639 4504 -1636
rect 4611 -1637 6944 -1636
rect 4474 -1642 4510 -1639
rect 4440 -1650 4456 -1648
rect 4214 -1662 4229 -1658
rect 4132 -1664 4229 -1662
rect 4257 -1664 4425 -1652
rect 4441 -1662 4456 -1658
rect 4474 -1661 4513 -1642
rect 4532 -1648 4539 -1647
rect 4538 -1655 4539 -1648
rect 4522 -1658 4523 -1655
rect 4538 -1658 4551 -1655
rect 4474 -1662 4504 -1661
rect 4513 -1662 4519 -1661
rect 4522 -1662 4551 -1658
rect 4441 -1663 4551 -1662
rect 4441 -1664 4557 -1663
rect 4116 -1672 4167 -1664
rect 4116 -1684 4141 -1672
rect 4148 -1684 4167 -1672
rect 4198 -1672 4248 -1664
rect 4198 -1680 4214 -1672
rect 4221 -1674 4248 -1672
rect 4257 -1674 4478 -1664
rect 4221 -1684 4478 -1674
rect 4507 -1672 4557 -1664
rect 4507 -1681 4523 -1672
rect 4116 -1692 4167 -1684
rect 4214 -1692 4478 -1684
rect 4504 -1684 4523 -1681
rect 4530 -1684 4557 -1672
rect 4504 -1692 4557 -1684
rect 4132 -1700 4133 -1692
rect 4148 -1700 4161 -1692
rect 4132 -1708 4148 -1700
rect 4129 -1715 4148 -1712
rect 4129 -1724 4151 -1715
rect 4102 -1734 4151 -1724
rect 4102 -1740 4132 -1734
rect 4151 -1739 4156 -1734
rect 4074 -1756 4148 -1740
rect 4166 -1748 4196 -1692
rect 4231 -1702 4439 -1692
rect 4474 -1696 4519 -1692
rect 4522 -1693 4523 -1692
rect 4538 -1693 4551 -1692
rect 4257 -1732 4446 -1702
rect 4272 -1735 4446 -1732
rect 4265 -1738 4446 -1735
rect 4074 -1758 4087 -1756
rect 4102 -1758 4136 -1756
rect 4074 -1774 4148 -1758
rect 4175 -1762 4188 -1748
rect 4203 -1762 4219 -1746
rect 4265 -1751 4276 -1738
rect 4058 -1796 4059 -1780
rect 4074 -1796 4087 -1774
rect 4102 -1796 4132 -1774
rect 4175 -1778 4237 -1762
rect 4265 -1769 4276 -1753
rect 4281 -1758 4291 -1738
rect 4301 -1758 4315 -1738
rect 4318 -1751 4327 -1738
rect 4343 -1751 4352 -1738
rect 4281 -1769 4315 -1758
rect 4318 -1769 4327 -1753
rect 4343 -1769 4352 -1753
rect 4359 -1758 4369 -1738
rect 4379 -1758 4393 -1738
rect 4394 -1751 4405 -1738
rect 4359 -1769 4393 -1758
rect 4394 -1769 4405 -1753
rect 4451 -1762 4467 -1746
rect 4474 -1748 4504 -1696
rect 4538 -1700 4539 -1693
rect 4523 -1708 4539 -1700
rect 4510 -1740 4523 -1721
rect 4538 -1740 4568 -1724
rect 4510 -1756 4584 -1740
rect 4510 -1758 4523 -1756
rect 4538 -1758 4572 -1756
rect 4175 -1780 4188 -1778
rect 4203 -1780 4237 -1778
rect 4175 -1796 4237 -1780
rect 4281 -1785 4297 -1778
rect 4359 -1785 4389 -1774
rect 4437 -1778 4483 -1762
rect 4510 -1774 4584 -1758
rect 4437 -1780 4471 -1778
rect 4436 -1796 4483 -1780
rect 4510 -1796 4523 -1774
rect 4538 -1796 4568 -1774
rect 4595 -1796 4596 -1780
rect 4611 -1796 4624 -1637
rect 4654 -1741 4667 -1637
rect 4712 -1659 4713 -1649
rect 4728 -1659 4741 -1649
rect 4712 -1663 4741 -1659
rect 4746 -1663 4776 -1637
rect 4794 -1651 4810 -1649
rect 4882 -1651 4935 -1637
rect 4883 -1653 4947 -1651
rect 4990 -1653 5005 -1637
rect 5054 -1640 5084 -1637
rect 5054 -1643 5090 -1640
rect 5020 -1651 5036 -1649
rect 4794 -1663 4809 -1659
rect 4712 -1665 4809 -1663
rect 4837 -1665 5005 -1653
rect 5021 -1663 5036 -1659
rect 5054 -1662 5093 -1643
rect 5112 -1649 5119 -1648
rect 5118 -1656 5119 -1649
rect 5102 -1659 5103 -1656
rect 5118 -1659 5131 -1656
rect 5054 -1663 5084 -1662
rect 5093 -1663 5099 -1662
rect 5102 -1663 5131 -1659
rect 5021 -1664 5131 -1663
rect 5021 -1665 5137 -1664
rect 4696 -1673 4747 -1665
rect 4696 -1685 4721 -1673
rect 4728 -1685 4747 -1673
rect 4778 -1673 4828 -1665
rect 4778 -1681 4794 -1673
rect 4801 -1675 4828 -1673
rect 4837 -1675 5058 -1665
rect 4801 -1685 5058 -1675
rect 5087 -1673 5137 -1665
rect 5087 -1682 5103 -1673
rect 4696 -1693 4747 -1685
rect 4794 -1693 5058 -1685
rect 5084 -1685 5103 -1682
rect 5110 -1685 5137 -1673
rect 5084 -1693 5137 -1685
rect 4712 -1701 4713 -1693
rect 4728 -1701 4741 -1693
rect 4712 -1709 4728 -1701
rect 4709 -1716 4728 -1713
rect 4709 -1725 4731 -1716
rect 4682 -1735 4731 -1725
rect 4682 -1741 4712 -1735
rect 4731 -1740 4736 -1735
rect 4654 -1757 4728 -1741
rect 4746 -1749 4776 -1693
rect 4811 -1703 5019 -1693
rect 5054 -1697 5099 -1693
rect 5102 -1694 5103 -1693
rect 5118 -1694 5131 -1693
rect 4837 -1733 5026 -1703
rect 4852 -1736 5026 -1733
rect 4845 -1739 5026 -1736
rect 4654 -1759 4667 -1757
rect 4682 -1759 4716 -1757
rect 4654 -1775 4728 -1759
rect 4755 -1763 4768 -1749
rect 4783 -1763 4799 -1747
rect 4845 -1752 4856 -1739
rect 3435 -1804 3470 -1796
rect 3435 -1830 3436 -1804
rect 3443 -1830 3470 -1804
rect 3379 -1848 3408 -1834
rect 3435 -1838 3470 -1830
rect 3472 -1804 3513 -1796
rect 3472 -1830 3487 -1804
rect 3494 -1830 3513 -1804
rect 3577 -1808 3639 -1796
rect 3651 -1808 3726 -1796
rect 3784 -1808 3859 -1796
rect 3871 -1808 3902 -1796
rect 3908 -1808 3943 -1796
rect 3577 -1810 3739 -1808
rect 3472 -1838 3513 -1830
rect 3595 -1834 3608 -1810
rect 3623 -1812 3638 -1810
rect 3435 -1848 3436 -1838
rect 3451 -1848 3464 -1838
rect 3478 -1848 3479 -1838
rect 3494 -1848 3507 -1838
rect 3522 -1848 3552 -1834
rect 3595 -1848 3638 -1834
rect 3662 -1837 3669 -1830
rect 3672 -1834 3739 -1810
rect 3771 -1810 3943 -1808
rect 3741 -1832 3769 -1828
rect 3771 -1832 3851 -1810
rect 3872 -1812 3887 -1810
rect 3741 -1834 3851 -1832
rect 3672 -1838 3851 -1834
rect 3645 -1848 3675 -1838
rect 3677 -1848 3830 -1838
rect 3838 -1848 3868 -1838
rect 3872 -1848 3902 -1834
rect 3930 -1848 3943 -1810
rect 4015 -1804 4050 -1796
rect 4015 -1830 4016 -1804
rect 4023 -1830 4050 -1804
rect 3958 -1848 3988 -1834
rect 4015 -1838 4050 -1830
rect 4052 -1804 4093 -1796
rect 4052 -1830 4067 -1804
rect 4074 -1830 4093 -1804
rect 4157 -1808 4219 -1796
rect 4231 -1808 4306 -1796
rect 4364 -1808 4439 -1796
rect 4451 -1808 4482 -1796
rect 4488 -1808 4523 -1796
rect 4157 -1810 4319 -1808
rect 4052 -1838 4093 -1830
rect 4175 -1834 4188 -1810
rect 4203 -1812 4218 -1810
rect 4015 -1848 4016 -1838
rect 4031 -1848 4044 -1838
rect 4058 -1848 4059 -1838
rect 4074 -1848 4087 -1838
rect 4102 -1848 4132 -1834
rect 4175 -1848 4218 -1834
rect 4242 -1837 4249 -1830
rect 4252 -1834 4319 -1810
rect 4351 -1810 4523 -1808
rect 4321 -1832 4349 -1828
rect 4351 -1832 4431 -1810
rect 4452 -1812 4467 -1810
rect 4321 -1834 4431 -1832
rect 4252 -1838 4431 -1834
rect 4225 -1848 4255 -1838
rect 4257 -1848 4410 -1838
rect 4418 -1848 4448 -1838
rect 4452 -1848 4482 -1834
rect 4510 -1848 4523 -1810
rect 4595 -1804 4630 -1796
rect 4638 -1797 4639 -1781
rect 4654 -1797 4667 -1775
rect 4682 -1797 4712 -1775
rect 4755 -1779 4817 -1763
rect 4845 -1770 4856 -1754
rect 4861 -1759 4871 -1739
rect 4881 -1759 4895 -1739
rect 4898 -1752 4907 -1739
rect 4923 -1752 4932 -1739
rect 4861 -1770 4895 -1759
rect 4898 -1770 4907 -1754
rect 4923 -1770 4932 -1754
rect 4939 -1759 4949 -1739
rect 4959 -1759 4973 -1739
rect 4974 -1752 4985 -1739
rect 4939 -1770 4973 -1759
rect 4974 -1770 4985 -1754
rect 5031 -1763 5047 -1747
rect 5054 -1749 5084 -1697
rect 5118 -1701 5119 -1694
rect 5103 -1709 5119 -1701
rect 5090 -1741 5103 -1722
rect 5118 -1741 5148 -1725
rect 5090 -1757 5164 -1741
rect 5090 -1759 5103 -1757
rect 5118 -1759 5152 -1757
rect 4755 -1781 4768 -1779
rect 4783 -1781 4817 -1779
rect 4755 -1797 4817 -1781
rect 4861 -1786 4877 -1779
rect 4939 -1786 4969 -1775
rect 5017 -1779 5063 -1763
rect 5090 -1775 5164 -1759
rect 5017 -1781 5051 -1779
rect 5016 -1797 5063 -1781
rect 5090 -1797 5103 -1775
rect 5118 -1797 5148 -1775
rect 5175 -1797 5176 -1781
rect 5191 -1797 5204 -1637
rect 5234 -1741 5247 -1637
rect 5292 -1659 5293 -1649
rect 5308 -1659 5321 -1649
rect 5292 -1663 5321 -1659
rect 5326 -1663 5356 -1637
rect 5374 -1651 5390 -1649
rect 5462 -1651 5515 -1637
rect 5463 -1653 5527 -1651
rect 5570 -1653 5585 -1637
rect 5634 -1640 5664 -1637
rect 5634 -1643 5670 -1640
rect 5600 -1651 5616 -1649
rect 5374 -1663 5389 -1659
rect 5292 -1665 5389 -1663
rect 5417 -1665 5585 -1653
rect 5601 -1663 5616 -1659
rect 5634 -1662 5673 -1643
rect 5692 -1649 5699 -1648
rect 5698 -1656 5699 -1649
rect 5682 -1659 5683 -1656
rect 5698 -1659 5711 -1656
rect 5634 -1663 5664 -1662
rect 5673 -1663 5679 -1662
rect 5682 -1663 5711 -1659
rect 5601 -1664 5711 -1663
rect 5601 -1665 5717 -1664
rect 5276 -1673 5327 -1665
rect 5276 -1685 5301 -1673
rect 5308 -1685 5327 -1673
rect 5358 -1673 5408 -1665
rect 5358 -1681 5374 -1673
rect 5381 -1675 5408 -1673
rect 5417 -1675 5638 -1665
rect 5381 -1685 5638 -1675
rect 5667 -1673 5717 -1665
rect 5667 -1682 5683 -1673
rect 5276 -1693 5327 -1685
rect 5374 -1693 5638 -1685
rect 5664 -1685 5683 -1682
rect 5690 -1685 5717 -1673
rect 5664 -1693 5717 -1685
rect 5292 -1701 5293 -1693
rect 5308 -1701 5321 -1693
rect 5292 -1709 5308 -1701
rect 5289 -1716 5308 -1713
rect 5289 -1725 5311 -1716
rect 5262 -1735 5311 -1725
rect 5262 -1741 5292 -1735
rect 5311 -1740 5316 -1735
rect 5234 -1757 5308 -1741
rect 5326 -1749 5356 -1693
rect 5391 -1703 5599 -1693
rect 5634 -1697 5679 -1693
rect 5682 -1694 5683 -1693
rect 5698 -1694 5711 -1693
rect 5417 -1733 5606 -1703
rect 5432 -1736 5606 -1733
rect 5425 -1739 5606 -1736
rect 5234 -1759 5247 -1757
rect 5262 -1759 5296 -1757
rect 5234 -1775 5308 -1759
rect 5335 -1763 5348 -1749
rect 5363 -1763 5379 -1747
rect 5425 -1752 5436 -1739
rect 5218 -1797 5219 -1781
rect 5234 -1797 5247 -1775
rect 5262 -1797 5292 -1775
rect 5335 -1779 5397 -1763
rect 5425 -1770 5436 -1754
rect 5441 -1759 5451 -1739
rect 5461 -1759 5475 -1739
rect 5478 -1752 5487 -1739
rect 5503 -1752 5512 -1739
rect 5441 -1770 5475 -1759
rect 5478 -1770 5487 -1754
rect 5503 -1770 5512 -1754
rect 5519 -1759 5529 -1739
rect 5539 -1759 5553 -1739
rect 5554 -1752 5565 -1739
rect 5519 -1770 5553 -1759
rect 5554 -1770 5565 -1754
rect 5611 -1763 5627 -1747
rect 5634 -1749 5664 -1697
rect 5698 -1701 5699 -1694
rect 5683 -1709 5699 -1701
rect 5670 -1741 5683 -1722
rect 5698 -1741 5728 -1725
rect 5670 -1757 5744 -1741
rect 5670 -1759 5683 -1757
rect 5698 -1759 5732 -1757
rect 5335 -1781 5348 -1779
rect 5363 -1781 5397 -1779
rect 5335 -1797 5397 -1781
rect 5441 -1786 5457 -1779
rect 5519 -1786 5549 -1775
rect 5597 -1779 5643 -1763
rect 5670 -1775 5744 -1759
rect 5597 -1781 5631 -1779
rect 5596 -1797 5643 -1781
rect 5670 -1797 5683 -1775
rect 5698 -1797 5728 -1775
rect 5755 -1797 5756 -1781
rect 5771 -1797 5784 -1637
rect 5814 -1741 5827 -1637
rect 5872 -1659 5873 -1649
rect 5888 -1659 5901 -1649
rect 5872 -1663 5901 -1659
rect 5906 -1663 5936 -1637
rect 5954 -1651 5970 -1649
rect 6042 -1651 6095 -1637
rect 6043 -1653 6107 -1651
rect 6150 -1653 6165 -1637
rect 6214 -1640 6244 -1637
rect 6214 -1643 6250 -1640
rect 6180 -1651 6196 -1649
rect 5954 -1663 5969 -1659
rect 5872 -1665 5969 -1663
rect 5997 -1665 6165 -1653
rect 6181 -1663 6196 -1659
rect 6214 -1662 6253 -1643
rect 6272 -1649 6279 -1648
rect 6278 -1656 6279 -1649
rect 6262 -1659 6263 -1656
rect 6278 -1659 6291 -1656
rect 6214 -1663 6244 -1662
rect 6253 -1663 6259 -1662
rect 6262 -1663 6291 -1659
rect 6181 -1664 6291 -1663
rect 6181 -1665 6297 -1664
rect 5856 -1673 5907 -1665
rect 5856 -1685 5881 -1673
rect 5888 -1685 5907 -1673
rect 5938 -1673 5988 -1665
rect 5938 -1681 5954 -1673
rect 5961 -1675 5988 -1673
rect 5997 -1675 6218 -1665
rect 5961 -1685 6218 -1675
rect 6247 -1673 6297 -1665
rect 6247 -1682 6263 -1673
rect 5856 -1693 5907 -1685
rect 5954 -1693 6218 -1685
rect 6244 -1685 6263 -1682
rect 6270 -1685 6297 -1673
rect 6244 -1693 6297 -1685
rect 5872 -1701 5873 -1693
rect 5888 -1701 5901 -1693
rect 5872 -1709 5888 -1701
rect 5869 -1716 5888 -1713
rect 5869 -1725 5891 -1716
rect 5842 -1735 5891 -1725
rect 5842 -1741 5872 -1735
rect 5891 -1740 5896 -1735
rect 5814 -1757 5888 -1741
rect 5906 -1749 5936 -1693
rect 5971 -1703 6179 -1693
rect 6214 -1697 6259 -1693
rect 6262 -1694 6263 -1693
rect 6278 -1694 6291 -1693
rect 5997 -1733 6186 -1703
rect 6012 -1736 6186 -1733
rect 6005 -1739 6186 -1736
rect 5814 -1759 5827 -1757
rect 5842 -1759 5876 -1757
rect 5814 -1775 5888 -1759
rect 5915 -1763 5928 -1749
rect 5943 -1763 5959 -1747
rect 6005 -1752 6016 -1739
rect 5798 -1797 5799 -1781
rect 5814 -1797 5827 -1775
rect 5842 -1797 5872 -1775
rect 5915 -1779 5977 -1763
rect 6005 -1770 6016 -1754
rect 6021 -1759 6031 -1739
rect 6041 -1759 6055 -1739
rect 6058 -1752 6067 -1739
rect 6083 -1752 6092 -1739
rect 6021 -1770 6055 -1759
rect 6058 -1770 6067 -1754
rect 6083 -1770 6092 -1754
rect 6099 -1759 6109 -1739
rect 6119 -1759 6133 -1739
rect 6134 -1752 6145 -1739
rect 6099 -1770 6133 -1759
rect 6134 -1770 6145 -1754
rect 6191 -1763 6207 -1747
rect 6214 -1749 6244 -1697
rect 6278 -1701 6279 -1694
rect 6263 -1709 6279 -1701
rect 6250 -1741 6263 -1722
rect 6278 -1741 6308 -1725
rect 6250 -1757 6324 -1741
rect 6250 -1759 6263 -1757
rect 6278 -1759 6312 -1757
rect 5915 -1781 5928 -1779
rect 5943 -1781 5977 -1779
rect 5915 -1797 5977 -1781
rect 6021 -1786 6037 -1779
rect 6099 -1786 6129 -1775
rect 6177 -1779 6223 -1763
rect 6250 -1775 6324 -1759
rect 6177 -1781 6211 -1779
rect 6176 -1797 6223 -1781
rect 6250 -1797 6263 -1775
rect 6278 -1797 6308 -1775
rect 6335 -1797 6336 -1781
rect 6351 -1797 6364 -1637
rect 6394 -1741 6407 -1637
rect 6452 -1659 6453 -1649
rect 6468 -1659 6481 -1649
rect 6452 -1663 6481 -1659
rect 6486 -1663 6516 -1637
rect 6534 -1651 6550 -1649
rect 6622 -1651 6675 -1637
rect 6623 -1653 6687 -1651
rect 6730 -1653 6745 -1637
rect 6794 -1640 6824 -1637
rect 6794 -1643 6830 -1640
rect 6760 -1651 6776 -1649
rect 6534 -1663 6549 -1659
rect 6452 -1665 6549 -1663
rect 6577 -1665 6745 -1653
rect 6761 -1663 6776 -1659
rect 6794 -1662 6833 -1643
rect 6852 -1649 6859 -1648
rect 6858 -1656 6859 -1649
rect 6842 -1659 6843 -1656
rect 6858 -1659 6871 -1656
rect 6794 -1663 6824 -1662
rect 6833 -1663 6839 -1662
rect 6842 -1663 6871 -1659
rect 6761 -1664 6871 -1663
rect 6761 -1665 6877 -1664
rect 6436 -1673 6487 -1665
rect 6436 -1685 6461 -1673
rect 6468 -1685 6487 -1673
rect 6518 -1673 6568 -1665
rect 6518 -1681 6534 -1673
rect 6541 -1675 6568 -1673
rect 6577 -1675 6798 -1665
rect 6541 -1685 6798 -1675
rect 6827 -1673 6877 -1665
rect 6827 -1682 6843 -1673
rect 6436 -1693 6487 -1685
rect 6534 -1693 6798 -1685
rect 6824 -1685 6843 -1682
rect 6850 -1685 6877 -1673
rect 6824 -1693 6877 -1685
rect 6452 -1701 6453 -1693
rect 6468 -1701 6481 -1693
rect 6452 -1709 6468 -1701
rect 6449 -1716 6468 -1713
rect 6449 -1725 6471 -1716
rect 6422 -1735 6471 -1725
rect 6422 -1741 6452 -1735
rect 6471 -1740 6476 -1735
rect 6394 -1757 6468 -1741
rect 6486 -1749 6516 -1693
rect 6551 -1703 6759 -1693
rect 6794 -1697 6839 -1693
rect 6842 -1694 6843 -1693
rect 6858 -1694 6871 -1693
rect 6577 -1733 6766 -1703
rect 6592 -1736 6766 -1733
rect 6585 -1739 6766 -1736
rect 6394 -1759 6407 -1757
rect 6422 -1759 6456 -1757
rect 6394 -1775 6468 -1759
rect 6495 -1763 6508 -1749
rect 6523 -1763 6539 -1747
rect 6585 -1752 6596 -1739
rect 6378 -1797 6379 -1781
rect 6394 -1797 6407 -1775
rect 6422 -1797 6452 -1775
rect 6495 -1779 6557 -1763
rect 6585 -1770 6596 -1754
rect 6601 -1759 6611 -1739
rect 6621 -1759 6635 -1739
rect 6638 -1752 6647 -1739
rect 6663 -1752 6672 -1739
rect 6601 -1770 6635 -1759
rect 6638 -1770 6647 -1754
rect 6663 -1770 6672 -1754
rect 6679 -1759 6689 -1739
rect 6699 -1759 6713 -1739
rect 6714 -1752 6725 -1739
rect 6679 -1770 6713 -1759
rect 6714 -1770 6725 -1754
rect 6771 -1763 6787 -1747
rect 6794 -1749 6824 -1697
rect 6858 -1701 6859 -1694
rect 6843 -1709 6859 -1701
rect 6830 -1741 6843 -1722
rect 6858 -1741 6888 -1725
rect 6830 -1757 6904 -1741
rect 6830 -1759 6843 -1757
rect 6858 -1759 6892 -1757
rect 6495 -1781 6508 -1779
rect 6523 -1781 6557 -1779
rect 6495 -1797 6557 -1781
rect 6601 -1786 6617 -1779
rect 6679 -1786 6709 -1775
rect 6757 -1779 6803 -1763
rect 6830 -1775 6904 -1759
rect 6757 -1781 6791 -1779
rect 6756 -1797 6803 -1781
rect 6830 -1797 6843 -1775
rect 6858 -1797 6888 -1775
rect 6915 -1797 6916 -1781
rect 6931 -1797 6944 -1637
rect 4595 -1830 4596 -1804
rect 4603 -1830 4630 -1804
rect 4538 -1848 4568 -1834
rect 4595 -1838 4630 -1830
rect 4632 -1805 4673 -1797
rect 4632 -1831 4647 -1805
rect 4654 -1831 4673 -1805
rect 4737 -1809 4799 -1797
rect 4811 -1809 4886 -1797
rect 4944 -1809 5019 -1797
rect 5031 -1809 5062 -1797
rect 5068 -1809 5103 -1797
rect 4737 -1811 4899 -1809
rect 4595 -1848 4596 -1838
rect 4611 -1848 4624 -1838
rect 4632 -1839 4673 -1831
rect 4755 -1835 4768 -1811
rect 4783 -1813 4798 -1811
rect 3379 -1849 4624 -1848
rect 4638 -1849 4639 -1839
rect 4654 -1849 4667 -1839
rect 4682 -1849 4712 -1835
rect 4755 -1849 4798 -1835
rect 4822 -1838 4829 -1831
rect 4832 -1835 4899 -1811
rect 4931 -1811 5103 -1809
rect 4901 -1833 4929 -1829
rect 4931 -1833 5011 -1811
rect 5032 -1813 5047 -1811
rect 4901 -1835 5011 -1833
rect 4832 -1839 5011 -1835
rect 4805 -1849 4835 -1839
rect 4837 -1849 4990 -1839
rect 4998 -1849 5028 -1839
rect 5032 -1849 5062 -1835
rect 5090 -1849 5103 -1811
rect 5175 -1805 5210 -1797
rect 5175 -1831 5176 -1805
rect 5183 -1831 5210 -1805
rect 5118 -1849 5148 -1835
rect 5175 -1839 5210 -1831
rect 5212 -1805 5253 -1797
rect 5212 -1831 5227 -1805
rect 5234 -1831 5253 -1805
rect 5317 -1809 5379 -1797
rect 5391 -1809 5466 -1797
rect 5524 -1809 5599 -1797
rect 5611 -1809 5642 -1797
rect 5648 -1809 5683 -1797
rect 5317 -1811 5479 -1809
rect 5212 -1839 5253 -1831
rect 5335 -1835 5348 -1811
rect 5363 -1813 5378 -1811
rect 5175 -1849 5176 -1839
rect 5191 -1849 5204 -1839
rect 5218 -1849 5219 -1839
rect 5234 -1849 5247 -1839
rect 5262 -1849 5292 -1835
rect 5335 -1849 5378 -1835
rect 5402 -1838 5409 -1831
rect 5412 -1835 5479 -1811
rect 5511 -1811 5683 -1809
rect 5481 -1833 5509 -1829
rect 5511 -1833 5591 -1811
rect 5612 -1813 5627 -1811
rect 5481 -1835 5591 -1833
rect 5412 -1839 5591 -1835
rect 5385 -1849 5415 -1839
rect 5417 -1849 5570 -1839
rect 5578 -1849 5608 -1839
rect 5612 -1849 5642 -1835
rect 5670 -1849 5683 -1811
rect 5755 -1805 5790 -1797
rect 5755 -1831 5756 -1805
rect 5763 -1831 5790 -1805
rect 5698 -1849 5728 -1835
rect 5755 -1839 5790 -1831
rect 5792 -1805 5833 -1797
rect 5792 -1831 5807 -1805
rect 5814 -1831 5833 -1805
rect 5897 -1809 5959 -1797
rect 5971 -1809 6046 -1797
rect 6104 -1809 6179 -1797
rect 6191 -1809 6222 -1797
rect 6228 -1809 6263 -1797
rect 5897 -1811 6059 -1809
rect 5792 -1839 5833 -1831
rect 5915 -1835 5928 -1811
rect 5943 -1813 5958 -1811
rect 5755 -1849 5756 -1839
rect 5771 -1849 5784 -1839
rect 5798 -1849 5799 -1839
rect 5814 -1849 5827 -1839
rect 5842 -1849 5872 -1835
rect 5915 -1849 5958 -1835
rect 5982 -1838 5989 -1831
rect 5992 -1835 6059 -1811
rect 6091 -1811 6263 -1809
rect 6061 -1833 6089 -1829
rect 6091 -1833 6171 -1811
rect 6192 -1813 6207 -1811
rect 6061 -1835 6171 -1833
rect 5992 -1839 6171 -1835
rect 5965 -1849 5995 -1839
rect 5997 -1849 6150 -1839
rect 6158 -1849 6188 -1839
rect 6192 -1849 6222 -1835
rect 6250 -1849 6263 -1811
rect 6335 -1805 6370 -1797
rect 6335 -1831 6336 -1805
rect 6343 -1831 6370 -1805
rect 6278 -1849 6308 -1835
rect 6335 -1839 6370 -1831
rect 6372 -1805 6413 -1797
rect 6372 -1831 6387 -1805
rect 6394 -1831 6413 -1805
rect 6477 -1809 6539 -1797
rect 6551 -1809 6626 -1797
rect 6684 -1809 6759 -1797
rect 6771 -1809 6802 -1797
rect 6808 -1809 6843 -1797
rect 6477 -1811 6639 -1809
rect 6372 -1839 6413 -1831
rect 6495 -1835 6508 -1811
rect 6523 -1813 6538 -1811
rect 6335 -1849 6336 -1839
rect 6351 -1849 6364 -1839
rect 6378 -1849 6379 -1839
rect 6394 -1849 6407 -1839
rect 6422 -1849 6452 -1835
rect 6495 -1849 6538 -1835
rect 6562 -1838 6569 -1831
rect 6572 -1835 6639 -1811
rect 6671 -1811 6843 -1809
rect 6641 -1833 6669 -1829
rect 6671 -1833 6751 -1811
rect 6772 -1813 6787 -1811
rect 6641 -1835 6751 -1833
rect 6572 -1839 6751 -1835
rect 6545 -1849 6575 -1839
rect 6577 -1849 6730 -1839
rect 6738 -1849 6768 -1839
rect 6772 -1849 6802 -1835
rect 6830 -1849 6843 -1811
rect 6915 -1805 6950 -1797
rect 6915 -1831 6916 -1805
rect 6923 -1831 6950 -1805
rect 6858 -1849 6888 -1835
rect 6915 -1839 6950 -1831
rect 6915 -1849 6916 -1839
rect 6931 -1849 6944 -1839
rect 3379 -1862 6944 -1849
rect 3379 -1880 3408 -1862
rect 3451 -1892 3464 -1862
rect 3494 -1892 3507 -1862
rect 3522 -1880 3552 -1862
rect 3595 -1876 3609 -1862
rect 3645 -1876 3865 -1862
rect 3596 -1878 3609 -1876
rect 3562 -1890 3577 -1878
rect 3559 -1892 3581 -1890
rect 3586 -1892 3616 -1878
rect 3677 -1880 3830 -1876
rect 3659 -1892 3851 -1880
rect 3894 -1892 3924 -1878
rect 3930 -1892 3943 -1862
rect 3958 -1880 3988 -1862
rect 4031 -1892 4044 -1862
rect 4074 -1892 4087 -1862
rect 4102 -1880 4132 -1862
rect 4175 -1876 4189 -1862
rect 4225 -1876 4445 -1862
rect 4176 -1878 4189 -1876
rect 4142 -1890 4157 -1878
rect 4139 -1892 4161 -1890
rect 4166 -1892 4196 -1878
rect 4257 -1880 4410 -1876
rect 4239 -1892 4431 -1880
rect 4474 -1892 4504 -1878
rect 4510 -1892 4523 -1862
rect 4538 -1880 4568 -1862
rect 4611 -1863 6944 -1862
rect 4611 -1892 4624 -1863
rect 3379 -1893 4624 -1892
rect 4654 -1893 4667 -1863
rect 4682 -1881 4712 -1863
rect 4755 -1877 4769 -1863
rect 4805 -1877 5025 -1863
rect 4756 -1879 4769 -1877
rect 4722 -1891 4737 -1879
rect 4719 -1893 4741 -1891
rect 4746 -1893 4776 -1879
rect 4837 -1881 4990 -1877
rect 4819 -1893 5011 -1881
rect 5054 -1893 5084 -1879
rect 5090 -1893 5103 -1863
rect 5118 -1881 5148 -1863
rect 5191 -1893 5204 -1863
rect 5234 -1893 5247 -1863
rect 5262 -1881 5292 -1863
rect 5335 -1877 5349 -1863
rect 5385 -1877 5605 -1863
rect 5336 -1879 5349 -1877
rect 5302 -1891 5317 -1879
rect 5299 -1893 5321 -1891
rect 5326 -1893 5356 -1879
rect 5417 -1881 5570 -1877
rect 5399 -1893 5591 -1881
rect 5634 -1893 5664 -1879
rect 5670 -1893 5683 -1863
rect 5698 -1881 5728 -1863
rect 5771 -1893 5784 -1863
rect 5814 -1893 5827 -1863
rect 5842 -1881 5872 -1863
rect 5915 -1877 5929 -1863
rect 5965 -1877 6185 -1863
rect 5916 -1879 5929 -1877
rect 5882 -1891 5897 -1879
rect 5879 -1893 5901 -1891
rect 5906 -1893 5936 -1879
rect 5997 -1881 6150 -1877
rect 5979 -1893 6171 -1881
rect 6214 -1893 6244 -1879
rect 6250 -1893 6263 -1863
rect 6278 -1881 6308 -1863
rect 6351 -1893 6364 -1863
rect 6394 -1893 6407 -1863
rect 6422 -1881 6452 -1863
rect 6495 -1877 6509 -1863
rect 6545 -1877 6765 -1863
rect 6496 -1879 6509 -1877
rect 6462 -1891 6477 -1879
rect 6459 -1893 6481 -1891
rect 6486 -1893 6516 -1879
rect 6577 -1881 6730 -1877
rect 6559 -1893 6751 -1881
rect 6794 -1893 6824 -1879
rect 6830 -1893 6843 -1863
rect 6858 -1881 6888 -1863
rect 6931 -1893 6944 -1863
rect 3379 -1906 6944 -1893
rect 3379 -1933 3391 -1925
rect 3379 -1962 3397 -1933
rect 3379 -1963 3391 -1962
rect 3379 -2010 3408 -1994
rect 3379 -2026 3424 -2010
rect 3379 -2028 3412 -2026
rect 3379 -2044 3424 -2028
rect 3379 -2066 3408 -2044
rect 3435 -2066 3436 -2050
rect 3451 -2066 3464 -1906
rect 3494 -2010 3507 -1906
rect 3552 -1928 3553 -1918
rect 3568 -1928 3581 -1918
rect 3552 -1932 3581 -1928
rect 3586 -1932 3616 -1906
rect 3634 -1920 3650 -1918
rect 3722 -1920 3775 -1906
rect 3723 -1922 3787 -1920
rect 3634 -1932 3649 -1928
rect 3552 -1934 3649 -1932
rect 3536 -1942 3587 -1934
rect 3536 -1954 3561 -1942
rect 3568 -1954 3587 -1942
rect 3618 -1942 3668 -1934
rect 3618 -1950 3634 -1942
rect 3641 -1944 3668 -1942
rect 3677 -1942 3692 -1938
rect 3739 -1942 3771 -1922
rect 3830 -1934 3845 -1906
rect 3894 -1909 3924 -1906
rect 3894 -1912 3930 -1909
rect 3860 -1920 3876 -1918
rect 3861 -1932 3876 -1928
rect 3894 -1931 3933 -1912
rect 3952 -1918 3959 -1917
rect 3958 -1925 3959 -1918
rect 3942 -1928 3943 -1925
rect 3958 -1928 3971 -1925
rect 3894 -1932 3924 -1931
rect 3933 -1932 3939 -1931
rect 3942 -1932 3971 -1928
rect 3861 -1933 3971 -1932
rect 3861 -1934 3977 -1933
rect 3830 -1942 3898 -1934
rect 3677 -1944 3746 -1942
rect 3764 -1944 3898 -1942
rect 3641 -1948 3713 -1944
rect 3641 -1950 3766 -1948
rect 3641 -1954 3713 -1950
rect 3536 -1962 3587 -1954
rect 3634 -1958 3713 -1954
rect 3794 -1958 3898 -1944
rect 3927 -1942 3977 -1934
rect 3927 -1951 3943 -1942
rect 3634 -1962 3898 -1958
rect 3924 -1954 3943 -1951
rect 3950 -1954 3977 -1942
rect 3924 -1962 3977 -1954
rect 3552 -1970 3553 -1962
rect 3568 -1970 3581 -1962
rect 3552 -1978 3568 -1970
rect 3549 -1985 3568 -1982
rect 3549 -1994 3571 -1985
rect 3522 -2004 3571 -1994
rect 3522 -2010 3552 -2004
rect 3571 -2009 3576 -2004
rect 3494 -2026 3568 -2010
rect 3586 -2018 3616 -1962
rect 3651 -1972 3859 -1962
rect 3894 -1966 3939 -1962
rect 3942 -1963 3943 -1962
rect 3958 -1963 3971 -1962
rect 3818 -1976 3866 -1972
rect 3701 -1998 3731 -1989
rect 3794 -1996 3809 -1989
rect 3830 -1998 3866 -1976
rect 3677 -2002 3866 -1998
rect 3692 -2005 3866 -2002
rect 3685 -2008 3866 -2005
rect 3494 -2028 3507 -2026
rect 3522 -2028 3556 -2026
rect 3494 -2044 3568 -2028
rect 3595 -2032 3608 -2018
rect 3623 -2032 3639 -2016
rect 3685 -2021 3696 -2008
rect 3478 -2066 3479 -2050
rect 3494 -2066 3507 -2044
rect 3522 -2066 3552 -2044
rect 3595 -2048 3657 -2032
rect 3685 -2039 3696 -2023
rect 3701 -2028 3711 -2008
rect 3721 -2028 3735 -2008
rect 3738 -2021 3747 -2008
rect 3763 -2021 3772 -2008
rect 3701 -2039 3735 -2028
rect 3738 -2039 3747 -2023
rect 3763 -2039 3772 -2023
rect 3779 -2028 3789 -2008
rect 3799 -2028 3813 -2008
rect 3814 -2021 3825 -2008
rect 3779 -2039 3813 -2028
rect 3814 -2039 3825 -2023
rect 3871 -2032 3887 -2016
rect 3894 -2018 3924 -1966
rect 3958 -1970 3959 -1963
rect 3943 -1978 3959 -1970
rect 3930 -2010 3943 -1991
rect 3958 -2010 3988 -1994
rect 3930 -2026 4004 -2010
rect 3930 -2028 3943 -2026
rect 3958 -2028 3992 -2026
rect 3595 -2050 3608 -2048
rect 3623 -2050 3657 -2048
rect 3595 -2066 3657 -2050
rect 3701 -2055 3717 -2048
rect 3779 -2055 3809 -2044
rect 3857 -2048 3903 -2032
rect 3930 -2044 4004 -2028
rect 3857 -2050 3891 -2048
rect 3856 -2066 3903 -2050
rect 3930 -2066 3943 -2044
rect 3958 -2066 3988 -2044
rect 4015 -2066 4016 -2050
rect 4031 -2066 4044 -1906
rect 4074 -2010 4087 -1906
rect 4132 -1928 4133 -1918
rect 4148 -1928 4161 -1918
rect 4132 -1932 4161 -1928
rect 4166 -1932 4196 -1906
rect 4214 -1920 4230 -1918
rect 4302 -1920 4355 -1906
rect 4303 -1922 4367 -1920
rect 4214 -1932 4229 -1928
rect 4132 -1934 4229 -1932
rect 4116 -1942 4167 -1934
rect 4116 -1954 4141 -1942
rect 4148 -1954 4167 -1942
rect 4198 -1942 4248 -1934
rect 4198 -1950 4214 -1942
rect 4221 -1944 4248 -1942
rect 4257 -1942 4272 -1938
rect 4319 -1942 4351 -1922
rect 4410 -1934 4425 -1906
rect 4474 -1909 4504 -1906
rect 4611 -1907 6944 -1906
rect 4474 -1912 4510 -1909
rect 4440 -1920 4456 -1918
rect 4441 -1932 4456 -1928
rect 4474 -1931 4513 -1912
rect 4532 -1918 4539 -1917
rect 4538 -1925 4539 -1918
rect 4522 -1928 4523 -1925
rect 4538 -1928 4551 -1925
rect 4474 -1932 4504 -1931
rect 4513 -1932 4519 -1931
rect 4522 -1932 4551 -1928
rect 4441 -1933 4551 -1932
rect 4441 -1934 4557 -1933
rect 4410 -1942 4478 -1934
rect 4257 -1944 4326 -1942
rect 4344 -1944 4478 -1942
rect 4221 -1948 4293 -1944
rect 4221 -1950 4346 -1948
rect 4221 -1954 4293 -1950
rect 4116 -1962 4167 -1954
rect 4214 -1958 4293 -1954
rect 4374 -1958 4478 -1944
rect 4507 -1942 4557 -1934
rect 4507 -1951 4523 -1942
rect 4214 -1962 4478 -1958
rect 4504 -1954 4523 -1951
rect 4530 -1954 4557 -1942
rect 4504 -1962 4557 -1954
rect 4132 -1970 4133 -1962
rect 4148 -1970 4161 -1962
rect 4132 -1978 4148 -1970
rect 4129 -1985 4148 -1982
rect 4129 -1994 4151 -1985
rect 4102 -2004 4151 -1994
rect 4102 -2010 4132 -2004
rect 4151 -2009 4156 -2004
rect 4074 -2026 4148 -2010
rect 4166 -2018 4196 -1962
rect 4231 -1972 4439 -1962
rect 4474 -1966 4519 -1962
rect 4522 -1963 4523 -1962
rect 4538 -1963 4551 -1962
rect 4398 -1976 4446 -1972
rect 4281 -1998 4311 -1989
rect 4374 -1996 4389 -1989
rect 4410 -1998 4446 -1976
rect 4257 -2002 4446 -1998
rect 4272 -2005 4446 -2002
rect 4265 -2008 4446 -2005
rect 4074 -2028 4087 -2026
rect 4102 -2028 4136 -2026
rect 4074 -2044 4148 -2028
rect 4175 -2032 4188 -2018
rect 4203 -2032 4219 -2016
rect 4265 -2021 4276 -2008
rect 4058 -2066 4059 -2050
rect 4074 -2066 4087 -2044
rect 4102 -2066 4132 -2044
rect 4175 -2048 4237 -2032
rect 4265 -2039 4276 -2023
rect 4281 -2028 4291 -2008
rect 4301 -2028 4315 -2008
rect 4318 -2021 4327 -2008
rect 4343 -2021 4352 -2008
rect 4281 -2039 4315 -2028
rect 4318 -2039 4327 -2023
rect 4343 -2039 4352 -2023
rect 4359 -2028 4369 -2008
rect 4379 -2028 4393 -2008
rect 4394 -2021 4405 -2008
rect 4359 -2039 4393 -2028
rect 4394 -2039 4405 -2023
rect 4451 -2032 4467 -2016
rect 4474 -2018 4504 -1966
rect 4538 -1970 4539 -1963
rect 4523 -1978 4539 -1970
rect 4510 -2010 4523 -1991
rect 4538 -2010 4568 -1994
rect 4510 -2026 4584 -2010
rect 4510 -2028 4523 -2026
rect 4538 -2028 4572 -2026
rect 4175 -2050 4188 -2048
rect 4203 -2050 4237 -2048
rect 4175 -2066 4237 -2050
rect 4281 -2055 4297 -2048
rect 4359 -2055 4389 -2044
rect 4437 -2048 4483 -2032
rect 4510 -2044 4584 -2028
rect 4437 -2050 4471 -2048
rect 4436 -2066 4483 -2050
rect 4510 -2066 4523 -2044
rect 4538 -2066 4568 -2044
rect 4595 -2066 4596 -2050
rect 4611 -2066 4624 -1907
rect 4654 -2011 4667 -1907
rect 4712 -1929 4713 -1919
rect 4728 -1929 4741 -1919
rect 4712 -1933 4741 -1929
rect 4746 -1933 4776 -1907
rect 4794 -1921 4810 -1919
rect 4882 -1921 4935 -1907
rect 4883 -1923 4947 -1921
rect 4794 -1933 4809 -1929
rect 4712 -1935 4809 -1933
rect 4696 -1943 4747 -1935
rect 4696 -1955 4721 -1943
rect 4728 -1955 4747 -1943
rect 4778 -1943 4828 -1935
rect 4778 -1951 4794 -1943
rect 4801 -1945 4828 -1943
rect 4837 -1943 4852 -1939
rect 4899 -1943 4931 -1923
rect 4990 -1935 5005 -1907
rect 5054 -1910 5084 -1907
rect 5054 -1913 5090 -1910
rect 5020 -1921 5036 -1919
rect 5021 -1933 5036 -1929
rect 5054 -1932 5093 -1913
rect 5112 -1919 5119 -1918
rect 5118 -1926 5119 -1919
rect 5102 -1929 5103 -1926
rect 5118 -1929 5131 -1926
rect 5054 -1933 5084 -1932
rect 5093 -1933 5099 -1932
rect 5102 -1933 5131 -1929
rect 5021 -1934 5131 -1933
rect 5021 -1935 5137 -1934
rect 4990 -1943 5058 -1935
rect 4837 -1945 4906 -1943
rect 4924 -1945 5058 -1943
rect 4801 -1949 4873 -1945
rect 4801 -1951 4926 -1949
rect 4801 -1955 4873 -1951
rect 4696 -1963 4747 -1955
rect 4794 -1959 4873 -1955
rect 4954 -1959 5058 -1945
rect 5087 -1943 5137 -1935
rect 5087 -1952 5103 -1943
rect 4794 -1963 5058 -1959
rect 5084 -1955 5103 -1952
rect 5110 -1955 5137 -1943
rect 5084 -1963 5137 -1955
rect 4712 -1971 4713 -1963
rect 4728 -1971 4741 -1963
rect 4712 -1979 4728 -1971
rect 4709 -1986 4728 -1983
rect 4709 -1995 4731 -1986
rect 4682 -2005 4731 -1995
rect 4682 -2011 4712 -2005
rect 4731 -2010 4736 -2005
rect 4654 -2027 4728 -2011
rect 4746 -2019 4776 -1963
rect 4811 -1973 5019 -1963
rect 5054 -1967 5099 -1963
rect 5102 -1964 5103 -1963
rect 5118 -1964 5131 -1963
rect 4978 -1977 5026 -1973
rect 4861 -1999 4891 -1990
rect 4954 -1997 4969 -1990
rect 4990 -1999 5026 -1977
rect 4837 -2003 5026 -1999
rect 4852 -2006 5026 -2003
rect 4845 -2009 5026 -2006
rect 4654 -2029 4667 -2027
rect 4682 -2029 4716 -2027
rect 4654 -2045 4728 -2029
rect 4755 -2033 4768 -2019
rect 4783 -2033 4799 -2017
rect 4845 -2022 4856 -2009
rect 3435 -2074 3470 -2066
rect 3435 -2100 3436 -2074
rect 3443 -2100 3470 -2074
rect 3435 -2108 3470 -2100
rect 3472 -2074 3513 -2066
rect 3472 -2100 3487 -2074
rect 3494 -2100 3513 -2074
rect 3577 -2078 3639 -2066
rect 3651 -2078 3726 -2066
rect 3784 -2078 3859 -2066
rect 3871 -2078 3902 -2066
rect 3908 -2078 3943 -2066
rect 3577 -2080 3739 -2078
rect 3472 -2108 3513 -2100
rect 3595 -2108 3608 -2080
rect 3623 -2082 3638 -2080
rect 3662 -2107 3669 -2100
rect 3672 -2108 3739 -2080
rect 3771 -2080 3943 -2078
rect 3741 -2102 3769 -2098
rect 3771 -2102 3851 -2080
rect 3872 -2082 3887 -2080
rect 3741 -2104 3851 -2102
rect 3741 -2108 3769 -2104
rect 3771 -2108 3851 -2104
rect 3379 -2118 3408 -2108
rect 3435 -2118 3436 -2108
rect 3451 -2118 3464 -2108
rect 3478 -2118 3479 -2108
rect 3494 -2118 3507 -2108
rect 3522 -2118 3552 -2108
rect 3595 -2118 3638 -2108
rect 3645 -2118 3653 -2108
rect 3672 -2116 3675 -2108
rect 3739 -2116 3771 -2108
rect 3672 -2118 3838 -2116
rect 3857 -2118 3868 -2108
rect 3872 -2118 3902 -2108
rect 3930 -2118 3943 -2080
rect 4015 -2074 4050 -2066
rect 4015 -2100 4016 -2074
rect 4023 -2100 4050 -2074
rect 4015 -2108 4050 -2100
rect 4052 -2074 4093 -2066
rect 4052 -2100 4067 -2074
rect 4074 -2100 4093 -2074
rect 4157 -2078 4219 -2066
rect 4231 -2078 4306 -2066
rect 4364 -2078 4439 -2066
rect 4451 -2078 4482 -2066
rect 4488 -2078 4523 -2066
rect 4157 -2080 4319 -2078
rect 4052 -2108 4093 -2100
rect 4175 -2108 4188 -2080
rect 4203 -2082 4218 -2080
rect 4242 -2107 4249 -2100
rect 4252 -2108 4319 -2080
rect 4351 -2080 4523 -2078
rect 4321 -2102 4349 -2098
rect 4351 -2102 4431 -2080
rect 4452 -2082 4467 -2080
rect 4321 -2104 4431 -2102
rect 4321 -2108 4349 -2104
rect 4351 -2108 4431 -2104
rect 3958 -2118 3988 -2108
rect 4015 -2118 4016 -2108
rect 4031 -2118 4044 -2108
rect 4058 -2118 4059 -2108
rect 4074 -2118 4087 -2108
rect 4102 -2118 4132 -2108
rect 4175 -2118 4218 -2108
rect 4225 -2118 4233 -2108
rect 4252 -2116 4255 -2108
rect 4319 -2116 4351 -2108
rect 4252 -2118 4418 -2116
rect 4437 -2118 4448 -2108
rect 4452 -2118 4482 -2108
rect 4510 -2118 4523 -2080
rect 4595 -2074 4630 -2066
rect 4638 -2067 4639 -2051
rect 4654 -2067 4667 -2045
rect 4682 -2067 4712 -2045
rect 4755 -2049 4817 -2033
rect 4845 -2040 4856 -2024
rect 4861 -2029 4871 -2009
rect 4881 -2029 4895 -2009
rect 4898 -2022 4907 -2009
rect 4923 -2022 4932 -2009
rect 4861 -2040 4895 -2029
rect 4898 -2040 4907 -2024
rect 4923 -2040 4932 -2024
rect 4939 -2029 4949 -2009
rect 4959 -2029 4973 -2009
rect 4974 -2022 4985 -2009
rect 4939 -2040 4973 -2029
rect 4974 -2040 4985 -2024
rect 5031 -2033 5047 -2017
rect 5054 -2019 5084 -1967
rect 5118 -1971 5119 -1964
rect 5103 -1979 5119 -1971
rect 5090 -2011 5103 -1992
rect 5118 -2011 5148 -1995
rect 5090 -2027 5164 -2011
rect 5090 -2029 5103 -2027
rect 5118 -2029 5152 -2027
rect 4755 -2051 4768 -2049
rect 4783 -2051 4817 -2049
rect 4755 -2067 4817 -2051
rect 4861 -2056 4877 -2049
rect 4939 -2056 4969 -2045
rect 5017 -2049 5063 -2033
rect 5090 -2045 5164 -2029
rect 5017 -2051 5051 -2049
rect 5016 -2067 5063 -2051
rect 5090 -2067 5103 -2045
rect 5118 -2067 5148 -2045
rect 5175 -2067 5176 -2051
rect 5191 -2067 5204 -1907
rect 5234 -2011 5247 -1907
rect 5292 -1929 5293 -1919
rect 5308 -1929 5321 -1919
rect 5292 -1933 5321 -1929
rect 5326 -1933 5356 -1907
rect 5374 -1921 5390 -1919
rect 5462 -1921 5515 -1907
rect 5463 -1923 5527 -1921
rect 5374 -1933 5389 -1929
rect 5292 -1935 5389 -1933
rect 5276 -1943 5327 -1935
rect 5276 -1955 5301 -1943
rect 5308 -1955 5327 -1943
rect 5358 -1943 5408 -1935
rect 5358 -1951 5374 -1943
rect 5381 -1945 5408 -1943
rect 5417 -1943 5432 -1939
rect 5479 -1943 5511 -1923
rect 5570 -1935 5585 -1907
rect 5634 -1910 5664 -1907
rect 5634 -1913 5670 -1910
rect 5600 -1921 5616 -1919
rect 5601 -1933 5616 -1929
rect 5634 -1932 5673 -1913
rect 5692 -1919 5699 -1918
rect 5698 -1926 5699 -1919
rect 5682 -1929 5683 -1926
rect 5698 -1929 5711 -1926
rect 5634 -1933 5664 -1932
rect 5673 -1933 5679 -1932
rect 5682 -1933 5711 -1929
rect 5601 -1934 5711 -1933
rect 5601 -1935 5717 -1934
rect 5570 -1943 5638 -1935
rect 5417 -1945 5486 -1943
rect 5504 -1945 5638 -1943
rect 5381 -1949 5453 -1945
rect 5381 -1951 5506 -1949
rect 5381 -1955 5453 -1951
rect 5276 -1963 5327 -1955
rect 5374 -1959 5453 -1955
rect 5534 -1959 5638 -1945
rect 5667 -1943 5717 -1935
rect 5667 -1952 5683 -1943
rect 5374 -1963 5638 -1959
rect 5664 -1955 5683 -1952
rect 5690 -1955 5717 -1943
rect 5664 -1963 5717 -1955
rect 5292 -1971 5293 -1963
rect 5308 -1971 5321 -1963
rect 5292 -1979 5308 -1971
rect 5289 -1986 5308 -1983
rect 5289 -1995 5311 -1986
rect 5262 -2005 5311 -1995
rect 5262 -2011 5292 -2005
rect 5311 -2010 5316 -2005
rect 5234 -2027 5308 -2011
rect 5326 -2019 5356 -1963
rect 5391 -1973 5599 -1963
rect 5634 -1967 5679 -1963
rect 5682 -1964 5683 -1963
rect 5698 -1964 5711 -1963
rect 5558 -1977 5606 -1973
rect 5441 -1999 5471 -1990
rect 5534 -1997 5549 -1990
rect 5570 -1999 5606 -1977
rect 5417 -2003 5606 -1999
rect 5432 -2006 5606 -2003
rect 5425 -2009 5606 -2006
rect 5234 -2029 5247 -2027
rect 5262 -2029 5296 -2027
rect 5234 -2045 5308 -2029
rect 5335 -2033 5348 -2019
rect 5363 -2033 5379 -2017
rect 5425 -2022 5436 -2009
rect 5218 -2067 5219 -2051
rect 5234 -2067 5247 -2045
rect 5262 -2067 5292 -2045
rect 5335 -2049 5397 -2033
rect 5425 -2040 5436 -2024
rect 5441 -2029 5451 -2009
rect 5461 -2029 5475 -2009
rect 5478 -2022 5487 -2009
rect 5503 -2022 5512 -2009
rect 5441 -2040 5475 -2029
rect 5478 -2040 5487 -2024
rect 5503 -2040 5512 -2024
rect 5519 -2029 5529 -2009
rect 5539 -2029 5553 -2009
rect 5554 -2022 5565 -2009
rect 5519 -2040 5553 -2029
rect 5554 -2040 5565 -2024
rect 5611 -2033 5627 -2017
rect 5634 -2019 5664 -1967
rect 5698 -1971 5699 -1964
rect 5683 -1979 5699 -1971
rect 5670 -2011 5683 -1992
rect 5698 -2011 5728 -1995
rect 5670 -2027 5744 -2011
rect 5670 -2029 5683 -2027
rect 5698 -2029 5732 -2027
rect 5335 -2051 5348 -2049
rect 5363 -2051 5397 -2049
rect 5335 -2067 5397 -2051
rect 5441 -2056 5457 -2049
rect 5519 -2056 5549 -2045
rect 5597 -2049 5643 -2033
rect 5670 -2045 5744 -2029
rect 5597 -2051 5631 -2049
rect 5596 -2067 5643 -2051
rect 5670 -2067 5683 -2045
rect 5698 -2067 5728 -2045
rect 5755 -2067 5756 -2051
rect 5771 -2067 5784 -1907
rect 5814 -2011 5827 -1907
rect 5872 -1929 5873 -1919
rect 5888 -1929 5901 -1919
rect 5872 -1933 5901 -1929
rect 5906 -1933 5936 -1907
rect 5954 -1921 5970 -1919
rect 6042 -1921 6095 -1907
rect 6043 -1923 6107 -1921
rect 5954 -1933 5969 -1929
rect 5872 -1935 5969 -1933
rect 5856 -1943 5907 -1935
rect 5856 -1955 5881 -1943
rect 5888 -1955 5907 -1943
rect 5938 -1943 5988 -1935
rect 5938 -1951 5954 -1943
rect 5961 -1945 5988 -1943
rect 5997 -1943 6012 -1939
rect 6059 -1943 6091 -1923
rect 6150 -1935 6165 -1907
rect 6214 -1910 6244 -1907
rect 6214 -1913 6250 -1910
rect 6180 -1921 6196 -1919
rect 6181 -1933 6196 -1929
rect 6214 -1932 6253 -1913
rect 6272 -1919 6279 -1918
rect 6278 -1926 6279 -1919
rect 6262 -1929 6263 -1926
rect 6278 -1929 6291 -1926
rect 6214 -1933 6244 -1932
rect 6253 -1933 6259 -1932
rect 6262 -1933 6291 -1929
rect 6181 -1934 6291 -1933
rect 6181 -1935 6297 -1934
rect 6150 -1943 6218 -1935
rect 5997 -1945 6066 -1943
rect 6084 -1945 6218 -1943
rect 5961 -1949 6033 -1945
rect 5961 -1951 6086 -1949
rect 5961 -1955 6033 -1951
rect 5856 -1963 5907 -1955
rect 5954 -1959 6033 -1955
rect 6114 -1959 6218 -1945
rect 6247 -1943 6297 -1935
rect 6247 -1952 6263 -1943
rect 5954 -1963 6218 -1959
rect 6244 -1955 6263 -1952
rect 6270 -1955 6297 -1943
rect 6244 -1963 6297 -1955
rect 5872 -1971 5873 -1963
rect 5888 -1971 5901 -1963
rect 5872 -1979 5888 -1971
rect 5869 -1986 5888 -1983
rect 5869 -1995 5891 -1986
rect 5842 -2005 5891 -1995
rect 5842 -2011 5872 -2005
rect 5891 -2010 5896 -2005
rect 5814 -2027 5888 -2011
rect 5906 -2019 5936 -1963
rect 5971 -1973 6179 -1963
rect 6214 -1967 6259 -1963
rect 6262 -1964 6263 -1963
rect 6278 -1964 6291 -1963
rect 6138 -1977 6186 -1973
rect 6021 -1999 6051 -1990
rect 6114 -1997 6129 -1990
rect 6150 -1999 6186 -1977
rect 5997 -2003 6186 -1999
rect 6012 -2006 6186 -2003
rect 6005 -2009 6186 -2006
rect 5814 -2029 5827 -2027
rect 5842 -2029 5876 -2027
rect 5814 -2045 5888 -2029
rect 5915 -2033 5928 -2019
rect 5943 -2033 5959 -2017
rect 6005 -2022 6016 -2009
rect 5798 -2067 5799 -2051
rect 5814 -2067 5827 -2045
rect 5842 -2067 5872 -2045
rect 5915 -2049 5977 -2033
rect 6005 -2040 6016 -2024
rect 6021 -2029 6031 -2009
rect 6041 -2029 6055 -2009
rect 6058 -2022 6067 -2009
rect 6083 -2022 6092 -2009
rect 6021 -2040 6055 -2029
rect 6058 -2040 6067 -2024
rect 6083 -2040 6092 -2024
rect 6099 -2029 6109 -2009
rect 6119 -2029 6133 -2009
rect 6134 -2022 6145 -2009
rect 6099 -2040 6133 -2029
rect 6134 -2040 6145 -2024
rect 6191 -2033 6207 -2017
rect 6214 -2019 6244 -1967
rect 6278 -1971 6279 -1964
rect 6263 -1979 6279 -1971
rect 6250 -2011 6263 -1992
rect 6278 -2011 6308 -1995
rect 6250 -2027 6324 -2011
rect 6250 -2029 6263 -2027
rect 6278 -2029 6312 -2027
rect 5915 -2051 5928 -2049
rect 5943 -2051 5977 -2049
rect 5915 -2067 5977 -2051
rect 6021 -2056 6037 -2049
rect 6099 -2056 6129 -2045
rect 6177 -2049 6223 -2033
rect 6250 -2045 6324 -2029
rect 6177 -2051 6211 -2049
rect 6176 -2067 6223 -2051
rect 6250 -2067 6263 -2045
rect 6278 -2067 6308 -2045
rect 6335 -2067 6336 -2051
rect 6351 -2067 6364 -1907
rect 6394 -2011 6407 -1907
rect 6452 -1929 6453 -1919
rect 6468 -1929 6481 -1919
rect 6452 -1933 6481 -1929
rect 6486 -1933 6516 -1907
rect 6534 -1921 6550 -1919
rect 6622 -1921 6675 -1907
rect 6623 -1923 6687 -1921
rect 6534 -1933 6549 -1929
rect 6452 -1935 6549 -1933
rect 6436 -1943 6487 -1935
rect 6436 -1955 6461 -1943
rect 6468 -1955 6487 -1943
rect 6518 -1943 6568 -1935
rect 6518 -1951 6534 -1943
rect 6541 -1945 6568 -1943
rect 6577 -1943 6592 -1939
rect 6639 -1943 6671 -1923
rect 6730 -1935 6745 -1907
rect 6794 -1910 6824 -1907
rect 6794 -1913 6830 -1910
rect 6760 -1921 6776 -1919
rect 6761 -1933 6776 -1929
rect 6794 -1932 6833 -1913
rect 6852 -1919 6859 -1918
rect 6858 -1926 6859 -1919
rect 6842 -1929 6843 -1926
rect 6858 -1929 6871 -1926
rect 6794 -1933 6824 -1932
rect 6833 -1933 6839 -1932
rect 6842 -1933 6871 -1929
rect 6761 -1934 6871 -1933
rect 6761 -1935 6877 -1934
rect 6730 -1943 6798 -1935
rect 6577 -1945 6646 -1943
rect 6664 -1945 6798 -1943
rect 6541 -1949 6613 -1945
rect 6541 -1951 6666 -1949
rect 6541 -1955 6613 -1951
rect 6436 -1963 6487 -1955
rect 6534 -1959 6613 -1955
rect 6694 -1959 6798 -1945
rect 6827 -1943 6877 -1935
rect 6827 -1952 6843 -1943
rect 6534 -1963 6798 -1959
rect 6824 -1955 6843 -1952
rect 6850 -1955 6877 -1943
rect 6824 -1963 6877 -1955
rect 6452 -1971 6453 -1963
rect 6468 -1971 6481 -1963
rect 6452 -1979 6468 -1971
rect 6449 -1986 6468 -1983
rect 6449 -1995 6471 -1986
rect 6422 -2005 6471 -1995
rect 6422 -2011 6452 -2005
rect 6471 -2010 6476 -2005
rect 6394 -2027 6468 -2011
rect 6486 -2019 6516 -1963
rect 6551 -1973 6759 -1963
rect 6794 -1967 6839 -1963
rect 6842 -1964 6843 -1963
rect 6858 -1964 6871 -1963
rect 6718 -1977 6766 -1973
rect 6601 -1999 6631 -1990
rect 6694 -1997 6709 -1990
rect 6730 -1999 6766 -1977
rect 6577 -2003 6766 -1999
rect 6592 -2006 6766 -2003
rect 6585 -2009 6766 -2006
rect 6394 -2029 6407 -2027
rect 6422 -2029 6456 -2027
rect 6394 -2045 6468 -2029
rect 6495 -2033 6508 -2019
rect 6523 -2033 6539 -2017
rect 6585 -2022 6596 -2009
rect 6378 -2067 6379 -2051
rect 6394 -2067 6407 -2045
rect 6422 -2067 6452 -2045
rect 6495 -2049 6557 -2033
rect 6585 -2040 6596 -2024
rect 6601 -2029 6611 -2009
rect 6621 -2029 6635 -2009
rect 6638 -2022 6647 -2009
rect 6663 -2022 6672 -2009
rect 6601 -2040 6635 -2029
rect 6638 -2040 6647 -2024
rect 6663 -2040 6672 -2024
rect 6679 -2029 6689 -2009
rect 6699 -2029 6713 -2009
rect 6714 -2022 6725 -2009
rect 6679 -2040 6713 -2029
rect 6714 -2040 6725 -2024
rect 6771 -2033 6787 -2017
rect 6794 -2019 6824 -1967
rect 6858 -1971 6859 -1964
rect 6843 -1979 6859 -1971
rect 6830 -2011 6843 -1992
rect 6858 -2011 6888 -1995
rect 6830 -2027 6904 -2011
rect 6830 -2029 6843 -2027
rect 6858 -2029 6892 -2027
rect 6495 -2051 6508 -2049
rect 6523 -2051 6557 -2049
rect 6495 -2067 6557 -2051
rect 6601 -2056 6617 -2049
rect 6679 -2056 6709 -2045
rect 6757 -2049 6803 -2033
rect 6830 -2045 6904 -2029
rect 6757 -2051 6791 -2049
rect 6756 -2067 6803 -2051
rect 6830 -2067 6843 -2045
rect 6858 -2067 6888 -2045
rect 6915 -2067 6916 -2051
rect 6931 -2067 6944 -1907
rect 4595 -2100 4596 -2074
rect 4603 -2100 4630 -2074
rect 4595 -2108 4630 -2100
rect 4632 -2075 4673 -2067
rect 4632 -2101 4647 -2075
rect 4654 -2101 4673 -2075
rect 4737 -2079 4799 -2067
rect 4811 -2079 4886 -2067
rect 4944 -2079 5019 -2067
rect 5031 -2079 5062 -2067
rect 5068 -2079 5103 -2067
rect 4737 -2081 4899 -2079
rect 4538 -2118 4568 -2108
rect 4595 -2118 4596 -2108
rect 4611 -2118 4624 -2108
rect 4632 -2109 4673 -2101
rect 4755 -2109 4768 -2081
rect 4783 -2083 4798 -2081
rect 4822 -2108 4829 -2101
rect 4832 -2109 4899 -2081
rect 4931 -2081 5103 -2079
rect 4901 -2103 4929 -2099
rect 4931 -2103 5011 -2081
rect 5032 -2083 5047 -2081
rect 4901 -2105 5011 -2103
rect 4901 -2109 4929 -2105
rect 4931 -2109 5011 -2105
rect 3379 -2119 4624 -2118
rect 4638 -2119 4639 -2109
rect 4654 -2119 4667 -2109
rect 4682 -2119 4712 -2109
rect 4755 -2119 4798 -2109
rect 4805 -2119 4813 -2109
rect 4832 -2117 4835 -2109
rect 4899 -2117 4931 -2109
rect 4832 -2119 4998 -2117
rect 5017 -2119 5028 -2109
rect 5032 -2119 5062 -2109
rect 5090 -2119 5103 -2081
rect 5175 -2075 5210 -2067
rect 5175 -2101 5176 -2075
rect 5183 -2101 5210 -2075
rect 5175 -2109 5210 -2101
rect 5212 -2075 5253 -2067
rect 5212 -2101 5227 -2075
rect 5234 -2101 5253 -2075
rect 5317 -2079 5379 -2067
rect 5391 -2079 5466 -2067
rect 5524 -2079 5599 -2067
rect 5611 -2079 5642 -2067
rect 5648 -2079 5683 -2067
rect 5317 -2081 5479 -2079
rect 5212 -2109 5253 -2101
rect 5335 -2109 5348 -2081
rect 5363 -2083 5378 -2081
rect 5402 -2108 5409 -2101
rect 5412 -2109 5479 -2081
rect 5511 -2081 5683 -2079
rect 5481 -2103 5509 -2099
rect 5511 -2103 5591 -2081
rect 5612 -2083 5627 -2081
rect 5481 -2105 5591 -2103
rect 5481 -2109 5509 -2105
rect 5511 -2109 5591 -2105
rect 5118 -2119 5148 -2109
rect 5175 -2119 5176 -2109
rect 5191 -2119 5204 -2109
rect 5218 -2119 5219 -2109
rect 5234 -2119 5247 -2109
rect 5262 -2119 5292 -2109
rect 5335 -2119 5378 -2109
rect 5385 -2119 5393 -2109
rect 5412 -2117 5415 -2109
rect 5479 -2117 5511 -2109
rect 5412 -2119 5578 -2117
rect 5597 -2119 5608 -2109
rect 5612 -2119 5642 -2109
rect 5670 -2119 5683 -2081
rect 5755 -2075 5790 -2067
rect 5755 -2101 5756 -2075
rect 5763 -2101 5790 -2075
rect 5755 -2109 5790 -2101
rect 5792 -2075 5833 -2067
rect 5792 -2101 5807 -2075
rect 5814 -2101 5833 -2075
rect 5897 -2079 5959 -2067
rect 5971 -2079 6046 -2067
rect 6104 -2079 6179 -2067
rect 6191 -2079 6222 -2067
rect 6228 -2079 6263 -2067
rect 5897 -2081 6059 -2079
rect 5792 -2109 5833 -2101
rect 5915 -2109 5928 -2081
rect 5943 -2083 5958 -2081
rect 5982 -2108 5989 -2101
rect 5992 -2109 6059 -2081
rect 6091 -2081 6263 -2079
rect 6061 -2103 6089 -2099
rect 6091 -2103 6171 -2081
rect 6192 -2083 6207 -2081
rect 6061 -2105 6171 -2103
rect 6061 -2109 6089 -2105
rect 6091 -2109 6171 -2105
rect 5698 -2119 5728 -2109
rect 5755 -2119 5756 -2109
rect 5771 -2119 5784 -2109
rect 5798 -2119 5799 -2109
rect 5814 -2119 5827 -2109
rect 5842 -2119 5872 -2109
rect 5915 -2119 5958 -2109
rect 5965 -2119 5973 -2109
rect 5992 -2117 5995 -2109
rect 6059 -2117 6091 -2109
rect 5992 -2119 6158 -2117
rect 6177 -2119 6188 -2109
rect 6192 -2119 6222 -2109
rect 6250 -2119 6263 -2081
rect 6335 -2075 6370 -2067
rect 6335 -2101 6336 -2075
rect 6343 -2101 6370 -2075
rect 6335 -2109 6370 -2101
rect 6372 -2075 6413 -2067
rect 6372 -2101 6387 -2075
rect 6394 -2101 6413 -2075
rect 6477 -2079 6539 -2067
rect 6551 -2079 6626 -2067
rect 6684 -2079 6759 -2067
rect 6771 -2079 6802 -2067
rect 6808 -2079 6843 -2067
rect 6477 -2081 6639 -2079
rect 6372 -2109 6413 -2101
rect 6495 -2109 6508 -2081
rect 6523 -2083 6538 -2081
rect 6562 -2108 6569 -2101
rect 6572 -2109 6639 -2081
rect 6671 -2081 6843 -2079
rect 6641 -2103 6669 -2099
rect 6671 -2103 6751 -2081
rect 6772 -2083 6787 -2081
rect 6641 -2105 6751 -2103
rect 6641 -2109 6669 -2105
rect 6671 -2109 6751 -2105
rect 6278 -2119 6308 -2109
rect 6335 -2119 6336 -2109
rect 6351 -2119 6364 -2109
rect 6378 -2119 6379 -2109
rect 6394 -2119 6407 -2109
rect 6422 -2119 6452 -2109
rect 6495 -2119 6538 -2109
rect 6545 -2119 6553 -2109
rect 6572 -2117 6575 -2109
rect 6639 -2117 6671 -2109
rect 6572 -2119 6738 -2117
rect 6757 -2119 6768 -2109
rect 6772 -2119 6802 -2109
rect 6830 -2119 6843 -2081
rect 6915 -2075 6950 -2067
rect 6915 -2101 6916 -2075
rect 6923 -2101 6950 -2075
rect 6915 -2109 6950 -2101
rect 6858 -2119 6888 -2109
rect 6915 -2119 6916 -2109
rect 6931 -2119 6944 -2109
rect 3379 -2132 6944 -2119
rect 3379 -2150 3408 -2132
rect 3451 -2146 3464 -2132
rect 3494 -2146 3507 -2132
rect 3522 -2150 3552 -2132
rect 3595 -2146 3608 -2132
rect 3645 -2145 3653 -2132
rect 3686 -2145 3824 -2132
rect 3857 -2145 3865 -2132
rect 3722 -2146 3773 -2145
rect 3930 -2146 3943 -2132
rect 3723 -2148 3787 -2146
rect 3958 -2150 3988 -2132
rect 4031 -2146 4044 -2132
rect 4074 -2146 4087 -2132
rect 4102 -2150 4132 -2132
rect 4175 -2146 4188 -2132
rect 4225 -2145 4233 -2132
rect 4266 -2145 4404 -2132
rect 4437 -2145 4445 -2132
rect 4302 -2146 4353 -2145
rect 4510 -2146 4523 -2132
rect 4303 -2148 4367 -2146
rect 4538 -2150 4568 -2132
rect 4611 -2133 6944 -2132
rect 4611 -2146 4624 -2133
rect 4654 -2147 4667 -2133
rect 4682 -2151 4712 -2133
rect 4755 -2147 4768 -2133
rect 4805 -2146 4813 -2133
rect 4846 -2146 4984 -2133
rect 5017 -2146 5025 -2133
rect 4882 -2147 4933 -2146
rect 5090 -2147 5103 -2133
rect 4883 -2149 4947 -2147
rect 5118 -2151 5148 -2133
rect 5191 -2147 5204 -2133
rect 5234 -2147 5247 -2133
rect 5262 -2151 5292 -2133
rect 5335 -2147 5348 -2133
rect 5385 -2146 5393 -2133
rect 5426 -2146 5564 -2133
rect 5597 -2146 5605 -2133
rect 5462 -2147 5513 -2146
rect 5670 -2147 5683 -2133
rect 5463 -2149 5527 -2147
rect 5698 -2151 5728 -2133
rect 5771 -2147 5784 -2133
rect 5814 -2147 5827 -2133
rect 5842 -2151 5872 -2133
rect 5915 -2147 5928 -2133
rect 5965 -2146 5973 -2133
rect 6006 -2146 6144 -2133
rect 6177 -2146 6185 -2133
rect 6042 -2147 6093 -2146
rect 6250 -2147 6263 -2133
rect 6043 -2149 6107 -2147
rect 6278 -2151 6308 -2133
rect 6351 -2147 6364 -2133
rect 6394 -2147 6407 -2133
rect 6422 -2151 6452 -2133
rect 6495 -2147 6508 -2133
rect 6545 -2146 6553 -2133
rect 6586 -2146 6724 -2133
rect 6757 -2146 6765 -2133
rect 6622 -2147 6673 -2146
rect 6830 -2147 6843 -2133
rect 6623 -2149 6687 -2147
rect 6858 -2151 6888 -2133
rect 6931 -2147 6944 -2133
<< nwell >>
rect 197 2048 350 2144
rect 777 2048 930 2144
rect 1357 2048 1510 2144
rect 1937 2048 2090 2144
rect 2517 2048 2670 2144
rect 3097 2048 3250 2144
rect 3677 2048 3830 2144
rect 4257 2048 4410 2144
rect 197 1778 350 1874
rect 777 1778 930 1874
rect 1357 1778 1510 1874
rect 1937 1778 2090 1874
rect 2517 1778 2670 1874
rect 3097 1778 3250 1874
rect 3677 1778 3830 1874
rect 4257 1778 4410 1874
rect 197 1508 350 1604
rect 777 1508 930 1604
rect 1357 1508 1510 1604
rect 1937 1508 2090 1604
rect 2517 1508 2670 1604
rect 3097 1508 3250 1604
rect 3677 1508 3830 1604
rect 4257 1508 4410 1604
rect 197 1238 350 1334
rect 777 1238 930 1334
rect 1357 1238 1510 1334
rect 1937 1238 2090 1334
rect 2517 1238 2670 1334
rect 3097 1238 3250 1334
rect 3677 1238 3830 1334
rect 4257 1238 4410 1334
rect 4837 2048 4990 2144
rect 5417 2048 5570 2144
rect 4837 1778 4990 1874
rect 5417 1778 5570 1874
rect 4837 1508 4990 1604
rect 5417 1508 5570 1604
rect 4837 1238 4990 1334
rect 5417 1238 5570 1334
rect 5997 2048 6150 2144
rect 6577 2048 6730 2144
rect 5997 1778 6150 1874
rect 6577 1778 6730 1874
rect 5997 1508 6150 1604
rect 6577 1508 6730 1604
rect 5997 1238 6150 1334
rect 6577 1238 6730 1334
rect 197 968 350 1064
rect 777 968 930 1064
rect 1357 968 1510 1064
rect 1937 968 2090 1064
rect 2517 968 2670 1064
rect 3097 968 3250 1064
rect 3677 968 3830 1064
rect 4257 968 4410 1064
rect 197 698 350 794
rect 777 698 930 794
rect 1357 698 1510 794
rect 1937 698 2090 794
rect 2517 698 2670 794
rect 3097 698 3250 794
rect 3677 698 3830 794
rect 4257 698 4410 794
rect 197 428 350 524
rect 777 428 930 524
rect 1357 428 1510 524
rect 1937 428 2090 524
rect 2517 428 2670 524
rect 3097 428 3250 524
rect 3677 428 3830 524
rect 4257 428 4410 524
rect 197 158 350 254
rect 777 158 930 254
rect 1357 158 1510 254
rect 1937 158 2090 254
rect 2517 158 2670 254
rect 3097 158 3250 254
rect 3677 158 3830 254
rect 4257 158 4410 254
rect 197 -112 350 -16
rect 777 -112 930 -16
rect 1357 -112 1510 -16
rect 1937 -112 2090 -16
rect 2517 -112 2670 -16
rect 3097 -112 3250 -16
rect 3677 -112 3830 -16
rect 4257 -112 4410 -16
rect 197 -382 350 -286
rect 777 -382 930 -286
rect 1357 -382 1510 -286
rect 1937 -382 2090 -286
rect 2517 -382 2670 -286
rect 3097 -382 3250 -286
rect 3677 -382 3830 -286
rect 4257 -382 4410 -286
rect 197 -652 350 -556
rect 777 -652 930 -556
rect 1357 -652 1510 -556
rect 1937 -652 2090 -556
rect 2517 -652 2670 -556
rect 3097 -652 3250 -556
rect 3677 -652 3830 -556
rect 4257 -652 4410 -556
rect 197 -922 350 -826
rect 777 -922 930 -826
rect 1357 -922 1510 -826
rect 1937 -922 2090 -826
rect 2517 -922 2670 -826
rect 3097 -922 3250 -826
rect 3677 -922 3830 -826
rect 4257 -922 4410 -826
rect 197 -1192 350 -1096
rect 777 -1192 930 -1096
rect 1357 -1192 1510 -1096
rect 1937 -1192 2090 -1096
rect 2517 -1192 2670 -1096
rect 3097 -1192 3250 -1096
rect 3677 -1192 3830 -1096
rect 4257 -1192 4410 -1096
rect 197 -1462 350 -1366
rect 777 -1462 930 -1366
rect 1357 -1462 1510 -1366
rect 1937 -1462 2090 -1366
rect 2517 -1462 2670 -1366
rect 3097 -1462 3250 -1366
rect 3677 -1462 3830 -1366
rect 4257 -1462 4410 -1366
rect 197 -1732 350 -1636
rect 777 -1732 930 -1636
rect 1357 -1732 1510 -1636
rect 1937 -1732 2090 -1636
rect 2517 -1732 2670 -1636
rect 3097 -1732 3250 -1636
rect 3677 -1732 3830 -1636
rect 4257 -1732 4410 -1636
rect 197 -2002 350 -1906
rect 777 -2002 930 -1906
rect 1357 -2002 1510 -1906
rect 1937 -2002 2090 -1906
rect 2517 -2002 2670 -1906
rect 3097 -2002 3250 -1906
rect 3677 -2002 3830 -1906
rect 4257 -2002 4410 -1906
rect 4837 967 4990 1063
rect 5417 967 5570 1063
rect 4837 697 4990 793
rect 5417 697 5570 793
rect 4837 427 4990 523
rect 5417 427 5570 523
rect 4837 157 4990 253
rect 5417 157 5570 253
rect 4837 -113 4990 -17
rect 5417 -113 5570 -17
rect 4837 -383 4990 -287
rect 5417 -383 5570 -287
rect 4837 -653 4990 -557
rect 5417 -653 5570 -557
rect 4837 -923 4990 -827
rect 5417 -923 5570 -827
rect 4837 -1193 4990 -1097
rect 5417 -1193 5570 -1097
rect 4837 -1463 4990 -1367
rect 5417 -1463 5570 -1367
rect 4837 -1733 4990 -1637
rect 5417 -1733 5570 -1637
rect 4837 -2003 4990 -1907
rect 5417 -2003 5570 -1907
rect 5997 967 6150 1063
rect 6577 967 6730 1063
rect 5997 697 6150 793
rect 6577 697 6730 793
rect 5997 427 6150 523
rect 6577 427 6730 523
rect 5997 157 6150 253
rect 6577 157 6730 253
rect 5997 -113 6150 -17
rect 6577 -113 6730 -17
rect 5997 -383 6150 -287
rect 6577 -383 6730 -287
rect 5997 -653 6150 -557
rect 6577 -653 6730 -557
rect 5997 -923 6150 -827
rect 6577 -923 6730 -827
rect 5997 -1193 6150 -1097
rect 6577 -1193 6730 -1097
rect 5997 -1463 6150 -1367
rect 6577 -1463 6730 -1367
rect 5997 -1733 6150 -1637
rect 6577 -1733 6730 -1637
rect 5997 -2003 6150 -1907
rect 6577 -2003 6730 -1907
<< pwell >>
rect -1 2002 169 2174
rect 381 2002 749 2174
rect 961 2002 1329 2174
rect 1541 2002 1909 2174
rect 2121 2002 2489 2174
rect 2701 2002 3069 2174
rect 3281 2002 3649 2174
rect 3861 2002 4229 2174
rect 4441 2002 4611 2174
rect -1 1904 4611 2002
rect -1 1732 169 1904
rect 381 1732 749 1904
rect 961 1732 1329 1904
rect 1541 1732 1909 1904
rect 2121 1732 2489 1904
rect 2701 1732 3069 1904
rect 3281 1732 3649 1904
rect 3861 1732 4229 1904
rect 4441 1732 4611 1904
rect -1 1634 4611 1732
rect -1 1462 169 1634
rect 381 1462 749 1634
rect 961 1462 1329 1634
rect 1541 1462 1909 1634
rect 2121 1462 2489 1634
rect 2701 1462 3069 1634
rect 3281 1462 3649 1634
rect 3861 1462 4229 1634
rect 4441 1462 4611 1634
rect -1 1364 4611 1462
rect -1 1192 169 1364
rect 381 1192 749 1364
rect 961 1192 1329 1364
rect 1541 1192 1909 1364
rect 2121 1192 2489 1364
rect 2701 1192 3069 1364
rect 3281 1192 3649 1364
rect 3861 1192 4229 1364
rect 4441 1192 4611 1364
rect -1 1094 4611 1192
rect 4639 2002 4809 2174
rect 5021 2002 5389 2174
rect 5601 2002 5771 2174
rect 4639 1904 5771 2002
rect 4639 1732 4809 1904
rect 5021 1732 5389 1904
rect 5601 1732 5771 1904
rect 4639 1634 5771 1732
rect 4639 1462 4809 1634
rect 5021 1462 5389 1634
rect 5601 1462 5771 1634
rect 4639 1364 5771 1462
rect 4639 1192 4809 1364
rect 5021 1192 5389 1364
rect 5601 1192 5771 1364
rect 4639 1094 5771 1192
rect 5799 2002 5969 2174
rect 6181 2002 6549 2174
rect 6761 2002 6931 2174
rect 5799 1904 6931 2002
rect 5799 1732 5969 1904
rect 6181 1732 6549 1904
rect 6761 1732 6931 1904
rect 5799 1634 6931 1732
rect 5799 1462 5969 1634
rect 6181 1462 6549 1634
rect 6761 1462 6931 1634
rect 5799 1364 6931 1462
rect 5799 1192 5969 1364
rect 6181 1192 6549 1364
rect 6761 1192 6931 1364
rect 5799 1094 6931 1192
rect -1 922 169 1094
rect 381 922 749 1094
rect 961 922 1329 1094
rect 1541 922 1909 1094
rect 2121 922 2489 1094
rect 2701 922 3069 1094
rect 3281 922 3649 1094
rect 3861 922 4229 1094
rect 4441 922 4611 1094
rect -1 824 4611 922
rect -1 652 169 824
rect 381 652 749 824
rect 961 652 1329 824
rect 1541 652 1909 824
rect 2121 652 2489 824
rect 2701 652 3069 824
rect 3281 652 3649 824
rect 3861 652 4229 824
rect 4441 652 4611 824
rect -1 554 4611 652
rect -1 382 169 554
rect 381 382 749 554
rect 961 382 1329 554
rect 1541 382 1909 554
rect 2121 382 2489 554
rect 2701 382 3069 554
rect 3281 382 3649 554
rect 3861 382 4229 554
rect 4441 382 4611 554
rect -1 284 4611 382
rect -1 112 169 284
rect 381 112 749 284
rect 961 112 1329 284
rect 1541 112 1909 284
rect 2121 112 2489 284
rect 2701 112 3069 284
rect 3281 112 3649 284
rect 3861 112 4229 284
rect 4441 112 4611 284
rect -1 14 4611 112
rect -1 -158 169 14
rect 381 -158 749 14
rect 961 -158 1329 14
rect 1541 -158 1909 14
rect 2121 -158 2489 14
rect 2701 -158 3069 14
rect 3281 -158 3649 14
rect 3861 -158 4229 14
rect 4441 -158 4611 14
rect -1 -256 4611 -158
rect -1 -428 169 -256
rect 381 -428 749 -256
rect 961 -428 1329 -256
rect 1541 -428 1909 -256
rect 2121 -428 2489 -256
rect 2701 -428 3069 -256
rect 3281 -428 3649 -256
rect 3861 -428 4229 -256
rect 4441 -428 4611 -256
rect -1 -526 4611 -428
rect -1 -698 169 -526
rect 381 -698 749 -526
rect 961 -698 1329 -526
rect 1541 -698 1909 -526
rect 2121 -698 2489 -526
rect 2701 -698 3069 -526
rect 3281 -698 3649 -526
rect 3861 -698 4229 -526
rect 4441 -698 4611 -526
rect -1 -796 4611 -698
rect -1 -968 169 -796
rect 381 -968 749 -796
rect 961 -968 1329 -796
rect 1541 -968 1909 -796
rect 2121 -968 2489 -796
rect 2701 -968 3069 -796
rect 3281 -968 3649 -796
rect 3861 -968 4229 -796
rect 4441 -968 4611 -796
rect -1 -1066 4611 -968
rect -1 -1238 169 -1066
rect 381 -1238 749 -1066
rect 961 -1238 1329 -1066
rect 1541 -1238 1909 -1066
rect 2121 -1238 2489 -1066
rect 2701 -1238 3069 -1066
rect 3281 -1238 3649 -1066
rect 3861 -1238 4229 -1066
rect 4441 -1238 4611 -1066
rect -1 -1336 4611 -1238
rect -1 -1508 169 -1336
rect 381 -1508 749 -1336
rect 961 -1508 1329 -1336
rect 1541 -1508 1909 -1336
rect 2121 -1508 2489 -1336
rect 2701 -1508 3069 -1336
rect 3281 -1508 3649 -1336
rect 3861 -1508 4229 -1336
rect 4441 -1508 4611 -1336
rect -1 -1606 4611 -1508
rect -1 -1778 169 -1606
rect 381 -1778 749 -1606
rect 961 -1778 1329 -1606
rect 1541 -1778 1909 -1606
rect 2121 -1778 2489 -1606
rect 2701 -1778 3069 -1606
rect 3281 -1778 3649 -1606
rect 3861 -1778 4229 -1606
rect 4441 -1778 4611 -1606
rect -1 -1876 4611 -1778
rect -1 -2048 169 -1876
rect 381 -2048 749 -1876
rect 961 -2048 1329 -1876
rect 1541 -2048 1909 -1876
rect 2121 -2048 2489 -1876
rect 2701 -2048 3069 -1876
rect 3281 -2048 3649 -1876
rect 3861 -2048 4229 -1876
rect 4441 -2048 4611 -1876
rect -1 -2146 4611 -2048
rect 4639 921 4809 1093
rect 5021 921 5389 1093
rect 5601 921 5771 1093
rect 4639 823 5771 921
rect 4639 651 4809 823
rect 5021 651 5389 823
rect 5601 651 5771 823
rect 4639 553 5771 651
rect 4639 381 4809 553
rect 5021 381 5389 553
rect 5601 381 5771 553
rect 4639 283 5771 381
rect 4639 111 4809 283
rect 5021 111 5389 283
rect 5601 111 5771 283
rect 4639 13 5771 111
rect 4639 -159 4809 13
rect 5021 -159 5389 13
rect 5601 -159 5771 13
rect 4639 -257 5771 -159
rect 4639 -429 4809 -257
rect 5021 -429 5389 -257
rect 5601 -429 5771 -257
rect 4639 -527 5771 -429
rect 4639 -699 4809 -527
rect 5021 -699 5389 -527
rect 5601 -699 5771 -527
rect 4639 -797 5771 -699
rect 4639 -969 4809 -797
rect 5021 -969 5389 -797
rect 5601 -969 5771 -797
rect 4639 -1067 5771 -969
rect 4639 -1239 4809 -1067
rect 5021 -1239 5389 -1067
rect 5601 -1239 5771 -1067
rect 4639 -1337 5771 -1239
rect 4639 -1509 4809 -1337
rect 5021 -1509 5389 -1337
rect 5601 -1509 5771 -1337
rect 4639 -1607 5771 -1509
rect 4639 -1779 4809 -1607
rect 5021 -1779 5389 -1607
rect 5601 -1779 5771 -1607
rect 4639 -1877 5771 -1779
rect 4639 -2049 4809 -1877
rect 5021 -2049 5389 -1877
rect 5601 -2049 5771 -1877
rect 4639 -2147 5771 -2049
rect 5799 921 5969 1093
rect 6181 921 6549 1093
rect 6761 921 6931 1093
rect 5799 823 6931 921
rect 5799 651 5969 823
rect 6181 651 6549 823
rect 6761 651 6931 823
rect 5799 553 6931 651
rect 5799 381 5969 553
rect 6181 381 6549 553
rect 6761 381 6931 553
rect 5799 283 6931 381
rect 5799 111 5969 283
rect 6181 111 6549 283
rect 6761 111 6931 283
rect 5799 13 6931 111
rect 5799 -159 5969 13
rect 6181 -159 6549 13
rect 6761 -159 6931 13
rect 5799 -257 6931 -159
rect 5799 -429 5969 -257
rect 6181 -429 6549 -257
rect 6761 -429 6931 -257
rect 5799 -527 6931 -429
rect 5799 -699 5969 -527
rect 6181 -699 6549 -527
rect 6761 -699 6931 -527
rect 5799 -797 6931 -699
rect 5799 -969 5969 -797
rect 6181 -969 6549 -797
rect 6761 -969 6931 -797
rect 5799 -1067 6931 -969
rect 5799 -1239 5969 -1067
rect 6181 -1239 6549 -1067
rect 6761 -1239 6931 -1067
rect 5799 -1337 6931 -1239
rect 5799 -1509 5969 -1337
rect 6181 -1509 6549 -1337
rect 6761 -1509 6931 -1337
rect 5799 -1607 6931 -1509
rect 5799 -1779 5969 -1607
rect 6181 -1779 6549 -1607
rect 6761 -1779 6931 -1607
rect 5799 -1877 6931 -1779
rect 5799 -2049 5969 -1877
rect 6181 -2049 6549 -1877
rect 6761 -2049 6931 -1877
rect 5799 -2147 6931 -2049
<< nmos >>
rect 106 2088 136 2116
rect 414 2088 444 2116
rect 686 2088 716 2116
rect 994 2088 1024 2116
rect 1266 2088 1296 2116
rect 1574 2088 1604 2116
rect 1846 2088 1876 2116
rect 2154 2088 2184 2116
rect 2426 2088 2456 2116
rect 2734 2088 2764 2116
rect 3006 2088 3036 2116
rect 3314 2088 3344 2116
rect 3586 2088 3616 2116
rect 3894 2088 3924 2116
rect 4166 2088 4196 2116
rect 4474 2088 4504 2116
rect 4746 2088 4776 2116
rect 5054 2088 5084 2116
rect 5326 2088 5356 2116
rect 5634 2088 5664 2116
rect 5906 2088 5936 2116
rect 6214 2088 6244 2116
rect 6486 2088 6516 2116
rect 6794 2088 6824 2116
rect 42 1942 72 1984
rect 478 1942 508 1984
rect 622 1942 652 1984
rect 1058 1942 1088 1984
rect 1202 1942 1232 1984
rect 1638 1942 1668 1984
rect 1782 1942 1812 1984
rect 2218 1942 2248 1984
rect 2362 1942 2392 1984
rect 2798 1942 2828 1984
rect 2942 1942 2972 1984
rect 3378 1942 3408 1984
rect 3522 1942 3552 1984
rect 3958 1942 3988 1984
rect 4102 1942 4132 1984
rect 4538 1942 4568 1984
rect 4682 1942 4712 1984
rect 5118 1942 5148 1984
rect 5262 1942 5292 1984
rect 5698 1942 5728 1984
rect 5842 1942 5872 1984
rect 6278 1942 6308 1984
rect 6422 1942 6452 1984
rect 6858 1942 6888 1984
rect 106 1818 136 1846
rect 414 1818 444 1846
rect 686 1818 716 1846
rect 994 1818 1024 1846
rect 1266 1818 1296 1846
rect 1574 1818 1604 1846
rect 1846 1818 1876 1846
rect 2154 1818 2184 1846
rect 2426 1818 2456 1846
rect 2734 1818 2764 1846
rect 3006 1818 3036 1846
rect 3314 1818 3344 1846
rect 3586 1818 3616 1846
rect 3894 1818 3924 1846
rect 4166 1818 4196 1846
rect 4474 1818 4504 1846
rect 4746 1818 4776 1846
rect 5054 1818 5084 1846
rect 5326 1818 5356 1846
rect 5634 1818 5664 1846
rect 5906 1818 5936 1846
rect 6214 1818 6244 1846
rect 6486 1818 6516 1846
rect 6794 1818 6824 1846
rect 42 1672 72 1714
rect 478 1672 508 1714
rect 622 1672 652 1714
rect 1058 1672 1088 1714
rect 1202 1672 1232 1714
rect 1638 1672 1668 1714
rect 1782 1672 1812 1714
rect 2218 1672 2248 1714
rect 2362 1672 2392 1714
rect 2798 1672 2828 1714
rect 2942 1672 2972 1714
rect 3378 1672 3408 1714
rect 3522 1672 3552 1714
rect 3958 1672 3988 1714
rect 4102 1672 4132 1714
rect 4538 1672 4568 1714
rect 4682 1672 4712 1714
rect 5118 1672 5148 1714
rect 5262 1672 5292 1714
rect 5698 1672 5728 1714
rect 5842 1672 5872 1714
rect 6278 1672 6308 1714
rect 6422 1672 6452 1714
rect 6858 1672 6888 1714
rect 106 1548 136 1576
rect 414 1548 444 1576
rect 686 1548 716 1576
rect 994 1548 1024 1576
rect 1266 1548 1296 1576
rect 1574 1548 1604 1576
rect 1846 1548 1876 1576
rect 2154 1548 2184 1576
rect 2426 1548 2456 1576
rect 2734 1548 2764 1576
rect 3006 1548 3036 1576
rect 3314 1548 3344 1576
rect 3586 1548 3616 1576
rect 3894 1548 3924 1576
rect 4166 1548 4196 1576
rect 4474 1548 4504 1576
rect 4746 1548 4776 1576
rect 5054 1548 5084 1576
rect 5326 1548 5356 1576
rect 5634 1548 5664 1576
rect 5906 1548 5936 1576
rect 6214 1548 6244 1576
rect 6486 1548 6516 1576
rect 6794 1548 6824 1576
rect 42 1402 72 1444
rect 478 1402 508 1444
rect 622 1402 652 1444
rect 1058 1402 1088 1444
rect 1202 1402 1232 1444
rect 1638 1402 1668 1444
rect 1782 1402 1812 1444
rect 2218 1402 2248 1444
rect 2362 1402 2392 1444
rect 2798 1402 2828 1444
rect 2942 1402 2972 1444
rect 3378 1402 3408 1444
rect 3522 1402 3552 1444
rect 3958 1402 3988 1444
rect 4102 1402 4132 1444
rect 4538 1402 4568 1444
rect 4682 1402 4712 1444
rect 5118 1402 5148 1444
rect 5262 1402 5292 1444
rect 5698 1402 5728 1444
rect 5842 1402 5872 1444
rect 6278 1402 6308 1444
rect 6422 1402 6452 1444
rect 6858 1402 6888 1444
rect 106 1278 136 1306
rect 414 1278 444 1306
rect 686 1278 716 1306
rect 994 1278 1024 1306
rect 1266 1278 1296 1306
rect 1574 1278 1604 1306
rect 1846 1278 1876 1306
rect 2154 1278 2184 1306
rect 2426 1278 2456 1306
rect 2734 1278 2764 1306
rect 3006 1278 3036 1306
rect 3314 1278 3344 1306
rect 3586 1278 3616 1306
rect 3894 1278 3924 1306
rect 4166 1278 4196 1306
rect 4474 1278 4504 1306
rect 4746 1278 4776 1306
rect 5054 1278 5084 1306
rect 5326 1278 5356 1306
rect 5634 1278 5664 1306
rect 5906 1278 5936 1306
rect 6214 1278 6244 1306
rect 6486 1278 6516 1306
rect 6794 1278 6824 1306
rect 42 1132 72 1174
rect 478 1132 508 1174
rect 622 1132 652 1174
rect 1058 1132 1088 1174
rect 1202 1132 1232 1174
rect 1638 1132 1668 1174
rect 1782 1132 1812 1174
rect 2218 1132 2248 1174
rect 2362 1132 2392 1174
rect 2798 1132 2828 1174
rect 2942 1132 2972 1174
rect 3378 1132 3408 1174
rect 3522 1132 3552 1174
rect 3958 1132 3988 1174
rect 4102 1132 4132 1174
rect 4538 1132 4568 1174
rect 4682 1132 4712 1174
rect 5118 1132 5148 1174
rect 5262 1132 5292 1174
rect 5698 1132 5728 1174
rect 5842 1132 5872 1174
rect 6278 1132 6308 1174
rect 6422 1132 6452 1174
rect 6858 1132 6888 1174
rect 106 1008 136 1036
rect 414 1008 444 1036
rect 686 1008 716 1036
rect 994 1008 1024 1036
rect 1266 1008 1296 1036
rect 1574 1008 1604 1036
rect 1846 1008 1876 1036
rect 2154 1008 2184 1036
rect 2426 1008 2456 1036
rect 2734 1008 2764 1036
rect 3006 1008 3036 1036
rect 3314 1008 3344 1036
rect 3586 1008 3616 1036
rect 3894 1008 3924 1036
rect 4166 1008 4196 1036
rect 4474 1008 4504 1036
rect 4746 1007 4776 1035
rect 5054 1007 5084 1035
rect 5326 1007 5356 1035
rect 42 862 72 904
rect 478 862 508 904
rect 622 862 652 904
rect 1058 862 1088 904
rect 1202 862 1232 904
rect 1638 862 1668 904
rect 1782 862 1812 904
rect 2218 862 2248 904
rect 2362 862 2392 904
rect 2798 862 2828 904
rect 2942 862 2972 904
rect 3378 862 3408 904
rect 3522 862 3552 904
rect 3958 862 3988 904
rect 4102 862 4132 904
rect 4538 862 4568 904
rect 5634 1007 5664 1035
rect 5906 1007 5936 1035
rect 6214 1007 6244 1035
rect 6486 1007 6516 1035
rect 6794 1007 6824 1035
rect 4682 861 4712 903
rect 5118 861 5148 903
rect 5262 861 5292 903
rect 5698 861 5728 903
rect 5842 861 5872 903
rect 6278 861 6308 903
rect 6422 861 6452 903
rect 6858 861 6888 903
rect 106 738 136 766
rect 414 738 444 766
rect 686 738 716 766
rect 994 738 1024 766
rect 1266 738 1296 766
rect 1574 738 1604 766
rect 1846 738 1876 766
rect 2154 738 2184 766
rect 2426 738 2456 766
rect 2734 738 2764 766
rect 3006 738 3036 766
rect 3314 738 3344 766
rect 3586 738 3616 766
rect 3894 738 3924 766
rect 4166 738 4196 766
rect 4474 738 4504 766
rect 4746 737 4776 765
rect 5054 737 5084 765
rect 5326 737 5356 765
rect 42 592 72 634
rect 478 592 508 634
rect 622 592 652 634
rect 1058 592 1088 634
rect 1202 592 1232 634
rect 1638 592 1668 634
rect 1782 592 1812 634
rect 2218 592 2248 634
rect 2362 592 2392 634
rect 2798 592 2828 634
rect 2942 592 2972 634
rect 3378 592 3408 634
rect 3522 592 3552 634
rect 3958 592 3988 634
rect 4102 592 4132 634
rect 4538 592 4568 634
rect 5634 737 5664 765
rect 5906 737 5936 765
rect 6214 737 6244 765
rect 6486 737 6516 765
rect 6794 737 6824 765
rect 4682 591 4712 633
rect 5118 591 5148 633
rect 5262 591 5292 633
rect 5698 591 5728 633
rect 5842 591 5872 633
rect 6278 591 6308 633
rect 6422 591 6452 633
rect 6858 591 6888 633
rect 106 468 136 496
rect 414 468 444 496
rect 686 468 716 496
rect 994 468 1024 496
rect 1266 468 1296 496
rect 1574 468 1604 496
rect 1846 468 1876 496
rect 2154 468 2184 496
rect 2426 468 2456 496
rect 2734 468 2764 496
rect 3006 468 3036 496
rect 3314 468 3344 496
rect 3586 468 3616 496
rect 3894 468 3924 496
rect 4166 468 4196 496
rect 4474 468 4504 496
rect 4746 467 4776 495
rect 5054 467 5084 495
rect 5326 467 5356 495
rect 42 322 72 364
rect 478 322 508 364
rect 622 322 652 364
rect 1058 322 1088 364
rect 1202 322 1232 364
rect 1638 322 1668 364
rect 1782 322 1812 364
rect 2218 322 2248 364
rect 2362 322 2392 364
rect 2798 322 2828 364
rect 2942 322 2972 364
rect 3378 322 3408 364
rect 3522 322 3552 364
rect 3958 322 3988 364
rect 4102 322 4132 364
rect 4538 322 4568 364
rect 5634 467 5664 495
rect 5906 467 5936 495
rect 6214 467 6244 495
rect 6486 467 6516 495
rect 6794 467 6824 495
rect 4682 321 4712 363
rect 5118 321 5148 363
rect 5262 321 5292 363
rect 5698 321 5728 363
rect 5842 321 5872 363
rect 6278 321 6308 363
rect 6422 321 6452 363
rect 6858 321 6888 363
rect 106 198 136 226
rect 414 198 444 226
rect 686 198 716 226
rect 994 198 1024 226
rect 1266 198 1296 226
rect 1574 198 1604 226
rect 1846 198 1876 226
rect 2154 198 2184 226
rect 2426 198 2456 226
rect 2734 198 2764 226
rect 3006 198 3036 226
rect 3314 198 3344 226
rect 3586 198 3616 226
rect 3894 198 3924 226
rect 4166 198 4196 226
rect 4474 198 4504 226
rect 4746 197 4776 225
rect 5054 197 5084 225
rect 5326 197 5356 225
rect 42 52 72 94
rect 478 52 508 94
rect 622 52 652 94
rect 1058 52 1088 94
rect 1202 52 1232 94
rect 1638 52 1668 94
rect 1782 52 1812 94
rect 2218 52 2248 94
rect 2362 52 2392 94
rect 2798 52 2828 94
rect 2942 52 2972 94
rect 3378 52 3408 94
rect 3522 52 3552 94
rect 3958 52 3988 94
rect 4102 52 4132 94
rect 4538 52 4568 94
rect 5634 197 5664 225
rect 5906 197 5936 225
rect 6214 197 6244 225
rect 6486 197 6516 225
rect 6794 197 6824 225
rect 4682 51 4712 93
rect 5118 51 5148 93
rect 5262 51 5292 93
rect 5698 51 5728 93
rect 5842 51 5872 93
rect 6278 51 6308 93
rect 6422 51 6452 93
rect 6858 51 6888 93
rect 106 -72 136 -44
rect 414 -72 444 -44
rect 686 -72 716 -44
rect 994 -72 1024 -44
rect 1266 -72 1296 -44
rect 1574 -72 1604 -44
rect 1846 -72 1876 -44
rect 2154 -72 2184 -44
rect 2426 -72 2456 -44
rect 2734 -72 2764 -44
rect 3006 -72 3036 -44
rect 3314 -72 3344 -44
rect 3586 -72 3616 -44
rect 3894 -72 3924 -44
rect 4166 -72 4196 -44
rect 4474 -72 4504 -44
rect 4746 -73 4776 -45
rect 5054 -73 5084 -45
rect 5326 -73 5356 -45
rect 42 -218 72 -176
rect 478 -218 508 -176
rect 622 -218 652 -176
rect 1058 -218 1088 -176
rect 1202 -218 1232 -176
rect 1638 -218 1668 -176
rect 1782 -218 1812 -176
rect 2218 -218 2248 -176
rect 2362 -218 2392 -176
rect 2798 -218 2828 -176
rect 2942 -218 2972 -176
rect 3378 -218 3408 -176
rect 3522 -218 3552 -176
rect 3958 -218 3988 -176
rect 4102 -218 4132 -176
rect 4538 -218 4568 -176
rect 5634 -73 5664 -45
rect 5906 -73 5936 -45
rect 6214 -73 6244 -45
rect 6486 -73 6516 -45
rect 6794 -73 6824 -45
rect 4682 -219 4712 -177
rect 5118 -219 5148 -177
rect 5262 -219 5292 -177
rect 5698 -219 5728 -177
rect 5842 -219 5872 -177
rect 6278 -219 6308 -177
rect 6422 -219 6452 -177
rect 6858 -219 6888 -177
rect 106 -342 136 -314
rect 414 -342 444 -314
rect 686 -342 716 -314
rect 994 -342 1024 -314
rect 1266 -342 1296 -314
rect 1574 -342 1604 -314
rect 1846 -342 1876 -314
rect 2154 -342 2184 -314
rect 2426 -342 2456 -314
rect 2734 -342 2764 -314
rect 3006 -342 3036 -314
rect 3314 -342 3344 -314
rect 3586 -342 3616 -314
rect 3894 -342 3924 -314
rect 4166 -342 4196 -314
rect 4474 -342 4504 -314
rect 4746 -343 4776 -315
rect 5054 -343 5084 -315
rect 5326 -343 5356 -315
rect 42 -488 72 -446
rect 478 -488 508 -446
rect 622 -488 652 -446
rect 1058 -488 1088 -446
rect 1202 -488 1232 -446
rect 1638 -488 1668 -446
rect 1782 -488 1812 -446
rect 2218 -488 2248 -446
rect 2362 -488 2392 -446
rect 2798 -488 2828 -446
rect 2942 -488 2972 -446
rect 3378 -488 3408 -446
rect 3522 -488 3552 -446
rect 3958 -488 3988 -446
rect 4102 -488 4132 -446
rect 4538 -488 4568 -446
rect 5634 -343 5664 -315
rect 5906 -343 5936 -315
rect 6214 -343 6244 -315
rect 6486 -343 6516 -315
rect 6794 -343 6824 -315
rect 4682 -489 4712 -447
rect 5118 -489 5148 -447
rect 5262 -489 5292 -447
rect 5698 -489 5728 -447
rect 5842 -489 5872 -447
rect 6278 -489 6308 -447
rect 6422 -489 6452 -447
rect 6858 -489 6888 -447
rect 106 -612 136 -584
rect 414 -612 444 -584
rect 686 -612 716 -584
rect 994 -612 1024 -584
rect 1266 -612 1296 -584
rect 1574 -612 1604 -584
rect 1846 -612 1876 -584
rect 2154 -612 2184 -584
rect 2426 -612 2456 -584
rect 2734 -612 2764 -584
rect 3006 -612 3036 -584
rect 3314 -612 3344 -584
rect 3586 -612 3616 -584
rect 3894 -612 3924 -584
rect 4166 -612 4196 -584
rect 4474 -612 4504 -584
rect 4746 -613 4776 -585
rect 5054 -613 5084 -585
rect 5326 -613 5356 -585
rect 42 -758 72 -716
rect 478 -758 508 -716
rect 622 -758 652 -716
rect 1058 -758 1088 -716
rect 1202 -758 1232 -716
rect 1638 -758 1668 -716
rect 1782 -758 1812 -716
rect 2218 -758 2248 -716
rect 2362 -758 2392 -716
rect 2798 -758 2828 -716
rect 2942 -758 2972 -716
rect 3378 -758 3408 -716
rect 3522 -758 3552 -716
rect 3958 -758 3988 -716
rect 4102 -758 4132 -716
rect 4538 -758 4568 -716
rect 5634 -613 5664 -585
rect 5906 -613 5936 -585
rect 6214 -613 6244 -585
rect 6486 -613 6516 -585
rect 6794 -613 6824 -585
rect 4682 -759 4712 -717
rect 5118 -759 5148 -717
rect 5262 -759 5292 -717
rect 5698 -759 5728 -717
rect 5842 -759 5872 -717
rect 6278 -759 6308 -717
rect 6422 -759 6452 -717
rect 6858 -759 6888 -717
rect 106 -882 136 -854
rect 414 -882 444 -854
rect 686 -882 716 -854
rect 994 -882 1024 -854
rect 1266 -882 1296 -854
rect 1574 -882 1604 -854
rect 1846 -882 1876 -854
rect 2154 -882 2184 -854
rect 2426 -882 2456 -854
rect 2734 -882 2764 -854
rect 3006 -882 3036 -854
rect 3314 -882 3344 -854
rect 3586 -882 3616 -854
rect 3894 -882 3924 -854
rect 4166 -882 4196 -854
rect 4474 -882 4504 -854
rect 4746 -883 4776 -855
rect 5054 -883 5084 -855
rect 5326 -883 5356 -855
rect 42 -1028 72 -986
rect 478 -1028 508 -986
rect 622 -1028 652 -986
rect 1058 -1028 1088 -986
rect 1202 -1028 1232 -986
rect 1638 -1028 1668 -986
rect 1782 -1028 1812 -986
rect 2218 -1028 2248 -986
rect 2362 -1028 2392 -986
rect 2798 -1028 2828 -986
rect 2942 -1028 2972 -986
rect 3378 -1028 3408 -986
rect 3522 -1028 3552 -986
rect 3958 -1028 3988 -986
rect 4102 -1028 4132 -986
rect 4538 -1028 4568 -986
rect 5634 -883 5664 -855
rect 5906 -883 5936 -855
rect 6214 -883 6244 -855
rect 6486 -883 6516 -855
rect 6794 -883 6824 -855
rect 4682 -1029 4712 -987
rect 5118 -1029 5148 -987
rect 5262 -1029 5292 -987
rect 5698 -1029 5728 -987
rect 5842 -1029 5872 -987
rect 6278 -1029 6308 -987
rect 6422 -1029 6452 -987
rect 6858 -1029 6888 -987
rect 106 -1152 136 -1124
rect 414 -1152 444 -1124
rect 686 -1152 716 -1124
rect 994 -1152 1024 -1124
rect 1266 -1152 1296 -1124
rect 1574 -1152 1604 -1124
rect 1846 -1152 1876 -1124
rect 2154 -1152 2184 -1124
rect 2426 -1152 2456 -1124
rect 2734 -1152 2764 -1124
rect 3006 -1152 3036 -1124
rect 3314 -1152 3344 -1124
rect 3586 -1152 3616 -1124
rect 3894 -1152 3924 -1124
rect 4166 -1152 4196 -1124
rect 4474 -1152 4504 -1124
rect 4746 -1153 4776 -1125
rect 5054 -1153 5084 -1125
rect 5326 -1153 5356 -1125
rect 42 -1298 72 -1256
rect 478 -1298 508 -1256
rect 622 -1298 652 -1256
rect 1058 -1298 1088 -1256
rect 1202 -1298 1232 -1256
rect 1638 -1298 1668 -1256
rect 1782 -1298 1812 -1256
rect 2218 -1298 2248 -1256
rect 2362 -1298 2392 -1256
rect 2798 -1298 2828 -1256
rect 2942 -1298 2972 -1256
rect 3378 -1298 3408 -1256
rect 3522 -1298 3552 -1256
rect 3958 -1298 3988 -1256
rect 4102 -1298 4132 -1256
rect 4538 -1298 4568 -1256
rect 5634 -1153 5664 -1125
rect 5906 -1153 5936 -1125
rect 6214 -1153 6244 -1125
rect 6486 -1153 6516 -1125
rect 6794 -1153 6824 -1125
rect 4682 -1299 4712 -1257
rect 5118 -1299 5148 -1257
rect 5262 -1299 5292 -1257
rect 5698 -1299 5728 -1257
rect 5842 -1299 5872 -1257
rect 6278 -1299 6308 -1257
rect 6422 -1299 6452 -1257
rect 6858 -1299 6888 -1257
rect 106 -1422 136 -1394
rect 414 -1422 444 -1394
rect 686 -1422 716 -1394
rect 994 -1422 1024 -1394
rect 1266 -1422 1296 -1394
rect 1574 -1422 1604 -1394
rect 1846 -1422 1876 -1394
rect 2154 -1422 2184 -1394
rect 2426 -1422 2456 -1394
rect 2734 -1422 2764 -1394
rect 3006 -1422 3036 -1394
rect 3314 -1422 3344 -1394
rect 3586 -1422 3616 -1394
rect 3894 -1422 3924 -1394
rect 4166 -1422 4196 -1394
rect 4474 -1422 4504 -1394
rect 4746 -1423 4776 -1395
rect 5054 -1423 5084 -1395
rect 5326 -1423 5356 -1395
rect 42 -1568 72 -1526
rect 478 -1568 508 -1526
rect 622 -1568 652 -1526
rect 1058 -1568 1088 -1526
rect 1202 -1568 1232 -1526
rect 1638 -1568 1668 -1526
rect 1782 -1568 1812 -1526
rect 2218 -1568 2248 -1526
rect 2362 -1568 2392 -1526
rect 2798 -1568 2828 -1526
rect 2942 -1568 2972 -1526
rect 3378 -1568 3408 -1526
rect 3522 -1568 3552 -1526
rect 3958 -1568 3988 -1526
rect 4102 -1568 4132 -1526
rect 4538 -1568 4568 -1526
rect 5634 -1423 5664 -1395
rect 5906 -1423 5936 -1395
rect 6214 -1423 6244 -1395
rect 6486 -1423 6516 -1395
rect 6794 -1423 6824 -1395
rect 4682 -1569 4712 -1527
rect 5118 -1569 5148 -1527
rect 5262 -1569 5292 -1527
rect 5698 -1569 5728 -1527
rect 5842 -1569 5872 -1527
rect 6278 -1569 6308 -1527
rect 6422 -1569 6452 -1527
rect 6858 -1569 6888 -1527
rect 106 -1692 136 -1664
rect 414 -1692 444 -1664
rect 686 -1692 716 -1664
rect 994 -1692 1024 -1664
rect 1266 -1692 1296 -1664
rect 1574 -1692 1604 -1664
rect 1846 -1692 1876 -1664
rect 2154 -1692 2184 -1664
rect 2426 -1692 2456 -1664
rect 2734 -1692 2764 -1664
rect 3006 -1692 3036 -1664
rect 3314 -1692 3344 -1664
rect 3586 -1692 3616 -1664
rect 3894 -1692 3924 -1664
rect 4166 -1692 4196 -1664
rect 4474 -1692 4504 -1664
rect 4746 -1693 4776 -1665
rect 5054 -1693 5084 -1665
rect 5326 -1693 5356 -1665
rect 42 -1838 72 -1796
rect 478 -1838 508 -1796
rect 622 -1838 652 -1796
rect 1058 -1838 1088 -1796
rect 1202 -1838 1232 -1796
rect 1638 -1838 1668 -1796
rect 1782 -1838 1812 -1796
rect 2218 -1838 2248 -1796
rect 2362 -1838 2392 -1796
rect 2798 -1838 2828 -1796
rect 2942 -1838 2972 -1796
rect 3378 -1838 3408 -1796
rect 3522 -1838 3552 -1796
rect 3958 -1838 3988 -1796
rect 4102 -1838 4132 -1796
rect 4538 -1838 4568 -1796
rect 5634 -1693 5664 -1665
rect 5906 -1693 5936 -1665
rect 6214 -1693 6244 -1665
rect 6486 -1693 6516 -1665
rect 6794 -1693 6824 -1665
rect 4682 -1839 4712 -1797
rect 5118 -1839 5148 -1797
rect 5262 -1839 5292 -1797
rect 5698 -1839 5728 -1797
rect 5842 -1839 5872 -1797
rect 6278 -1839 6308 -1797
rect 6422 -1839 6452 -1797
rect 6858 -1839 6888 -1797
rect 106 -1962 136 -1934
rect 414 -1962 444 -1934
rect 686 -1962 716 -1934
rect 994 -1962 1024 -1934
rect 1266 -1962 1296 -1934
rect 1574 -1962 1604 -1934
rect 1846 -1962 1876 -1934
rect 2154 -1962 2184 -1934
rect 2426 -1962 2456 -1934
rect 2734 -1962 2764 -1934
rect 3006 -1962 3036 -1934
rect 3314 -1962 3344 -1934
rect 3586 -1962 3616 -1934
rect 3894 -1962 3924 -1934
rect 4166 -1962 4196 -1934
rect 4474 -1962 4504 -1934
rect 4746 -1963 4776 -1935
rect 5054 -1963 5084 -1935
rect 5326 -1963 5356 -1935
rect 42 -2108 72 -2066
rect 478 -2108 508 -2066
rect 622 -2108 652 -2066
rect 1058 -2108 1088 -2066
rect 1202 -2108 1232 -2066
rect 1638 -2108 1668 -2066
rect 1782 -2108 1812 -2066
rect 2218 -2108 2248 -2066
rect 2362 -2108 2392 -2066
rect 2798 -2108 2828 -2066
rect 2942 -2108 2972 -2066
rect 3378 -2108 3408 -2066
rect 3522 -2108 3552 -2066
rect 3958 -2108 3988 -2066
rect 4102 -2108 4132 -2066
rect 4538 -2108 4568 -2066
rect 5634 -1963 5664 -1935
rect 5906 -1963 5936 -1935
rect 6214 -1963 6244 -1935
rect 6486 -1963 6516 -1935
rect 6794 -1963 6824 -1935
rect 4682 -2109 4712 -2067
rect 5118 -2109 5148 -2067
rect 5262 -2109 5292 -2067
rect 5698 -2109 5728 -2067
rect 5842 -2109 5872 -2067
rect 6278 -2109 6308 -2067
rect 6422 -2109 6452 -2067
rect 6858 -2109 6888 -2067
<< npd >>
rect 221 1942 251 1984
rect 299 1942 329 1984
rect 801 1942 831 1984
rect 879 1942 909 1984
rect 1381 1942 1411 1984
rect 1459 1942 1489 1984
rect 1961 1942 1991 1984
rect 2039 1942 2069 1984
rect 2541 1942 2571 1984
rect 2619 1942 2649 1984
rect 3121 1942 3151 1984
rect 3199 1942 3229 1984
rect 3701 1942 3731 1984
rect 3779 1942 3809 1984
rect 4281 1942 4311 1984
rect 4359 1942 4389 1984
rect 4861 1942 4891 1984
rect 4939 1942 4969 1984
rect 5441 1942 5471 1984
rect 5519 1942 5549 1984
rect 6021 1942 6051 1984
rect 6099 1942 6129 1984
rect 6601 1942 6631 1984
rect 6679 1942 6709 1984
rect 221 1672 251 1714
rect 299 1672 329 1714
rect 801 1672 831 1714
rect 879 1672 909 1714
rect 1381 1672 1411 1714
rect 1459 1672 1489 1714
rect 1961 1672 1991 1714
rect 2039 1672 2069 1714
rect 2541 1672 2571 1714
rect 2619 1672 2649 1714
rect 3121 1672 3151 1714
rect 3199 1672 3229 1714
rect 3701 1672 3731 1714
rect 3779 1672 3809 1714
rect 4281 1672 4311 1714
rect 4359 1672 4389 1714
rect 4861 1672 4891 1714
rect 4939 1672 4969 1714
rect 5441 1672 5471 1714
rect 5519 1672 5549 1714
rect 6021 1672 6051 1714
rect 6099 1672 6129 1714
rect 6601 1672 6631 1714
rect 6679 1672 6709 1714
rect 221 1402 251 1444
rect 299 1402 329 1444
rect 801 1402 831 1444
rect 879 1402 909 1444
rect 1381 1402 1411 1444
rect 1459 1402 1489 1444
rect 1961 1402 1991 1444
rect 2039 1402 2069 1444
rect 2541 1402 2571 1444
rect 2619 1402 2649 1444
rect 3121 1402 3151 1444
rect 3199 1402 3229 1444
rect 3701 1402 3731 1444
rect 3779 1402 3809 1444
rect 4281 1402 4311 1444
rect 4359 1402 4389 1444
rect 4861 1402 4891 1444
rect 4939 1402 4969 1444
rect 5441 1402 5471 1444
rect 5519 1402 5549 1444
rect 6021 1402 6051 1444
rect 6099 1402 6129 1444
rect 6601 1402 6631 1444
rect 6679 1402 6709 1444
rect 221 1132 251 1174
rect 299 1132 329 1174
rect 801 1132 831 1174
rect 879 1132 909 1174
rect 1381 1132 1411 1174
rect 1459 1132 1489 1174
rect 1961 1132 1991 1174
rect 2039 1132 2069 1174
rect 2541 1132 2571 1174
rect 2619 1132 2649 1174
rect 3121 1132 3151 1174
rect 3199 1132 3229 1174
rect 3701 1132 3731 1174
rect 3779 1132 3809 1174
rect 4281 1132 4311 1174
rect 4359 1132 4389 1174
rect 4861 1132 4891 1174
rect 4939 1132 4969 1174
rect 5441 1132 5471 1174
rect 5519 1132 5549 1174
rect 6021 1132 6051 1174
rect 6099 1132 6129 1174
rect 6601 1132 6631 1174
rect 6679 1132 6709 1174
rect 221 862 251 904
rect 299 862 329 904
rect 801 862 831 904
rect 879 862 909 904
rect 1381 862 1411 904
rect 1459 862 1489 904
rect 1961 862 1991 904
rect 2039 862 2069 904
rect 2541 862 2571 904
rect 2619 862 2649 904
rect 3121 862 3151 904
rect 3199 862 3229 904
rect 3701 862 3731 904
rect 3779 862 3809 904
rect 4281 862 4311 904
rect 4359 862 4389 904
rect 4861 861 4891 903
rect 4939 861 4969 903
rect 5441 861 5471 903
rect 5519 861 5549 903
rect 6021 861 6051 903
rect 6099 861 6129 903
rect 6601 861 6631 903
rect 6679 861 6709 903
rect 221 592 251 634
rect 299 592 329 634
rect 801 592 831 634
rect 879 592 909 634
rect 1381 592 1411 634
rect 1459 592 1489 634
rect 1961 592 1991 634
rect 2039 592 2069 634
rect 2541 592 2571 634
rect 2619 592 2649 634
rect 3121 592 3151 634
rect 3199 592 3229 634
rect 3701 592 3731 634
rect 3779 592 3809 634
rect 4281 592 4311 634
rect 4359 592 4389 634
rect 4861 591 4891 633
rect 4939 591 4969 633
rect 5441 591 5471 633
rect 5519 591 5549 633
rect 6021 591 6051 633
rect 6099 591 6129 633
rect 6601 591 6631 633
rect 6679 591 6709 633
rect 221 322 251 364
rect 299 322 329 364
rect 801 322 831 364
rect 879 322 909 364
rect 1381 322 1411 364
rect 1459 322 1489 364
rect 1961 322 1991 364
rect 2039 322 2069 364
rect 2541 322 2571 364
rect 2619 322 2649 364
rect 3121 322 3151 364
rect 3199 322 3229 364
rect 3701 322 3731 364
rect 3779 322 3809 364
rect 4281 322 4311 364
rect 4359 322 4389 364
rect 4861 321 4891 363
rect 4939 321 4969 363
rect 5441 321 5471 363
rect 5519 321 5549 363
rect 6021 321 6051 363
rect 6099 321 6129 363
rect 6601 321 6631 363
rect 6679 321 6709 363
rect 221 52 251 94
rect 299 52 329 94
rect 801 52 831 94
rect 879 52 909 94
rect 1381 52 1411 94
rect 1459 52 1489 94
rect 1961 52 1991 94
rect 2039 52 2069 94
rect 2541 52 2571 94
rect 2619 52 2649 94
rect 3121 52 3151 94
rect 3199 52 3229 94
rect 3701 52 3731 94
rect 3779 52 3809 94
rect 4281 52 4311 94
rect 4359 52 4389 94
rect 4861 51 4891 93
rect 4939 51 4969 93
rect 5441 51 5471 93
rect 5519 51 5549 93
rect 6021 51 6051 93
rect 6099 51 6129 93
rect 6601 51 6631 93
rect 6679 51 6709 93
rect 221 -218 251 -176
rect 299 -218 329 -176
rect 801 -218 831 -176
rect 879 -218 909 -176
rect 1381 -218 1411 -176
rect 1459 -218 1489 -176
rect 1961 -218 1991 -176
rect 2039 -218 2069 -176
rect 2541 -218 2571 -176
rect 2619 -218 2649 -176
rect 3121 -218 3151 -176
rect 3199 -218 3229 -176
rect 3701 -218 3731 -176
rect 3779 -218 3809 -176
rect 4281 -218 4311 -176
rect 4359 -218 4389 -176
rect 4861 -219 4891 -177
rect 4939 -219 4969 -177
rect 5441 -219 5471 -177
rect 5519 -219 5549 -177
rect 6021 -219 6051 -177
rect 6099 -219 6129 -177
rect 6601 -219 6631 -177
rect 6679 -219 6709 -177
rect 221 -488 251 -446
rect 299 -488 329 -446
rect 801 -488 831 -446
rect 879 -488 909 -446
rect 1381 -488 1411 -446
rect 1459 -488 1489 -446
rect 1961 -488 1991 -446
rect 2039 -488 2069 -446
rect 2541 -488 2571 -446
rect 2619 -488 2649 -446
rect 3121 -488 3151 -446
rect 3199 -488 3229 -446
rect 3701 -488 3731 -446
rect 3779 -488 3809 -446
rect 4281 -488 4311 -446
rect 4359 -488 4389 -446
rect 4861 -489 4891 -447
rect 4939 -489 4969 -447
rect 5441 -489 5471 -447
rect 5519 -489 5549 -447
rect 6021 -489 6051 -447
rect 6099 -489 6129 -447
rect 6601 -489 6631 -447
rect 6679 -489 6709 -447
rect 221 -758 251 -716
rect 299 -758 329 -716
rect 801 -758 831 -716
rect 879 -758 909 -716
rect 1381 -758 1411 -716
rect 1459 -758 1489 -716
rect 1961 -758 1991 -716
rect 2039 -758 2069 -716
rect 2541 -758 2571 -716
rect 2619 -758 2649 -716
rect 3121 -758 3151 -716
rect 3199 -758 3229 -716
rect 3701 -758 3731 -716
rect 3779 -758 3809 -716
rect 4281 -758 4311 -716
rect 4359 -758 4389 -716
rect 4861 -759 4891 -717
rect 4939 -759 4969 -717
rect 5441 -759 5471 -717
rect 5519 -759 5549 -717
rect 6021 -759 6051 -717
rect 6099 -759 6129 -717
rect 6601 -759 6631 -717
rect 6679 -759 6709 -717
rect 221 -1028 251 -986
rect 299 -1028 329 -986
rect 801 -1028 831 -986
rect 879 -1028 909 -986
rect 1381 -1028 1411 -986
rect 1459 -1028 1489 -986
rect 1961 -1028 1991 -986
rect 2039 -1028 2069 -986
rect 2541 -1028 2571 -986
rect 2619 -1028 2649 -986
rect 3121 -1028 3151 -986
rect 3199 -1028 3229 -986
rect 3701 -1028 3731 -986
rect 3779 -1028 3809 -986
rect 4281 -1028 4311 -986
rect 4359 -1028 4389 -986
rect 4861 -1029 4891 -987
rect 4939 -1029 4969 -987
rect 5441 -1029 5471 -987
rect 5519 -1029 5549 -987
rect 6021 -1029 6051 -987
rect 6099 -1029 6129 -987
rect 6601 -1029 6631 -987
rect 6679 -1029 6709 -987
rect 221 -1298 251 -1256
rect 299 -1298 329 -1256
rect 801 -1298 831 -1256
rect 879 -1298 909 -1256
rect 1381 -1298 1411 -1256
rect 1459 -1298 1489 -1256
rect 1961 -1298 1991 -1256
rect 2039 -1298 2069 -1256
rect 2541 -1298 2571 -1256
rect 2619 -1298 2649 -1256
rect 3121 -1298 3151 -1256
rect 3199 -1298 3229 -1256
rect 3701 -1298 3731 -1256
rect 3779 -1298 3809 -1256
rect 4281 -1298 4311 -1256
rect 4359 -1298 4389 -1256
rect 4861 -1299 4891 -1257
rect 4939 -1299 4969 -1257
rect 5441 -1299 5471 -1257
rect 5519 -1299 5549 -1257
rect 6021 -1299 6051 -1257
rect 6099 -1299 6129 -1257
rect 6601 -1299 6631 -1257
rect 6679 -1299 6709 -1257
rect 221 -1568 251 -1526
rect 299 -1568 329 -1526
rect 801 -1568 831 -1526
rect 879 -1568 909 -1526
rect 1381 -1568 1411 -1526
rect 1459 -1568 1489 -1526
rect 1961 -1568 1991 -1526
rect 2039 -1568 2069 -1526
rect 2541 -1568 2571 -1526
rect 2619 -1568 2649 -1526
rect 3121 -1568 3151 -1526
rect 3199 -1568 3229 -1526
rect 3701 -1568 3731 -1526
rect 3779 -1568 3809 -1526
rect 4281 -1568 4311 -1526
rect 4359 -1568 4389 -1526
rect 4861 -1569 4891 -1527
rect 4939 -1569 4969 -1527
rect 5441 -1569 5471 -1527
rect 5519 -1569 5549 -1527
rect 6021 -1569 6051 -1527
rect 6099 -1569 6129 -1527
rect 6601 -1569 6631 -1527
rect 6679 -1569 6709 -1527
rect 221 -1838 251 -1796
rect 299 -1838 329 -1796
rect 801 -1838 831 -1796
rect 879 -1838 909 -1796
rect 1381 -1838 1411 -1796
rect 1459 -1838 1489 -1796
rect 1961 -1838 1991 -1796
rect 2039 -1838 2069 -1796
rect 2541 -1838 2571 -1796
rect 2619 -1838 2649 -1796
rect 3121 -1838 3151 -1796
rect 3199 -1838 3229 -1796
rect 3701 -1838 3731 -1796
rect 3779 -1838 3809 -1796
rect 4281 -1838 4311 -1796
rect 4359 -1838 4389 -1796
rect 4861 -1839 4891 -1797
rect 4939 -1839 4969 -1797
rect 5441 -1839 5471 -1797
rect 5519 -1839 5549 -1797
rect 6021 -1839 6051 -1797
rect 6099 -1839 6129 -1797
rect 6601 -1839 6631 -1797
rect 6679 -1839 6709 -1797
rect 221 -2108 251 -2066
rect 299 -2108 329 -2066
rect 801 -2108 831 -2066
rect 879 -2108 909 -2066
rect 1381 -2108 1411 -2066
rect 1459 -2108 1489 -2066
rect 1961 -2108 1991 -2066
rect 2039 -2108 2069 -2066
rect 2541 -2108 2571 -2066
rect 2619 -2108 2649 -2066
rect 3121 -2108 3151 -2066
rect 3199 -2108 3229 -2066
rect 3701 -2108 3731 -2066
rect 3779 -2108 3809 -2066
rect 4281 -2108 4311 -2066
rect 4359 -2108 4389 -2066
rect 4861 -2109 4891 -2067
rect 4939 -2109 4969 -2067
rect 5441 -2109 5471 -2067
rect 5519 -2109 5549 -2067
rect 6021 -2109 6051 -2067
rect 6099 -2109 6129 -2067
rect 6601 -2109 6631 -2067
rect 6679 -2109 6709 -2067
<< npass >>
rect 128 1942 158 1970
rect 392 1942 422 1970
rect 708 1942 738 1970
rect 972 1942 1002 1970
rect 1288 1942 1318 1970
rect 1552 1942 1582 1970
rect 1868 1942 1898 1970
rect 2132 1942 2162 1970
rect 2448 1942 2478 1970
rect 2712 1942 2742 1970
rect 3028 1942 3058 1970
rect 3292 1942 3322 1970
rect 3608 1942 3638 1970
rect 3872 1942 3902 1970
rect 4188 1942 4218 1970
rect 4452 1942 4482 1970
rect 4768 1942 4798 1970
rect 5032 1942 5062 1970
rect 5348 1942 5378 1970
rect 5612 1942 5642 1970
rect 5928 1942 5958 1970
rect 6192 1942 6222 1970
rect 6508 1942 6538 1970
rect 6772 1942 6802 1970
rect 128 1672 158 1700
rect 392 1672 422 1700
rect 708 1672 738 1700
rect 972 1672 1002 1700
rect 1288 1672 1318 1700
rect 1552 1672 1582 1700
rect 1868 1672 1898 1700
rect 2132 1672 2162 1700
rect 2448 1672 2478 1700
rect 2712 1672 2742 1700
rect 3028 1672 3058 1700
rect 3292 1672 3322 1700
rect 3608 1672 3638 1700
rect 3872 1672 3902 1700
rect 4188 1672 4218 1700
rect 4452 1672 4482 1700
rect 4768 1672 4798 1700
rect 5032 1672 5062 1700
rect 5348 1672 5378 1700
rect 5612 1672 5642 1700
rect 5928 1672 5958 1700
rect 6192 1672 6222 1700
rect 6508 1672 6538 1700
rect 6772 1672 6802 1700
rect 128 1402 158 1430
rect 392 1402 422 1430
rect 708 1402 738 1430
rect 972 1402 1002 1430
rect 1288 1402 1318 1430
rect 1552 1402 1582 1430
rect 1868 1402 1898 1430
rect 2132 1402 2162 1430
rect 2448 1402 2478 1430
rect 2712 1402 2742 1430
rect 3028 1402 3058 1430
rect 3292 1402 3322 1430
rect 3608 1402 3638 1430
rect 3872 1402 3902 1430
rect 4188 1402 4218 1430
rect 4452 1402 4482 1430
rect 4768 1402 4798 1430
rect 5032 1402 5062 1430
rect 5348 1402 5378 1430
rect 5612 1402 5642 1430
rect 5928 1402 5958 1430
rect 6192 1402 6222 1430
rect 6508 1402 6538 1430
rect 6772 1402 6802 1430
rect 128 1132 158 1160
rect 392 1132 422 1160
rect 708 1132 738 1160
rect 972 1132 1002 1160
rect 1288 1132 1318 1160
rect 1552 1132 1582 1160
rect 1868 1132 1898 1160
rect 2132 1132 2162 1160
rect 2448 1132 2478 1160
rect 2712 1132 2742 1160
rect 3028 1132 3058 1160
rect 3292 1132 3322 1160
rect 3608 1132 3638 1160
rect 3872 1132 3902 1160
rect 4188 1132 4218 1160
rect 4452 1132 4482 1160
rect 4768 1132 4798 1160
rect 5032 1132 5062 1160
rect 5348 1132 5378 1160
rect 5612 1132 5642 1160
rect 5928 1132 5958 1160
rect 6192 1132 6222 1160
rect 6508 1132 6538 1160
rect 6772 1132 6802 1160
rect 128 862 158 890
rect 392 862 422 890
rect 708 862 738 890
rect 972 862 1002 890
rect 1288 862 1318 890
rect 1552 862 1582 890
rect 1868 862 1898 890
rect 2132 862 2162 890
rect 2448 862 2478 890
rect 2712 862 2742 890
rect 3028 862 3058 890
rect 3292 862 3322 890
rect 3608 862 3638 890
rect 3872 862 3902 890
rect 4188 862 4218 890
rect 4452 862 4482 890
rect 4768 861 4798 889
rect 5032 861 5062 889
rect 5348 861 5378 889
rect 5612 861 5642 889
rect 5928 861 5958 889
rect 6192 861 6222 889
rect 6508 861 6538 889
rect 6772 861 6802 889
rect 128 592 158 620
rect 392 592 422 620
rect 708 592 738 620
rect 972 592 1002 620
rect 1288 592 1318 620
rect 1552 592 1582 620
rect 1868 592 1898 620
rect 2132 592 2162 620
rect 2448 592 2478 620
rect 2712 592 2742 620
rect 3028 592 3058 620
rect 3292 592 3322 620
rect 3608 592 3638 620
rect 3872 592 3902 620
rect 4188 592 4218 620
rect 4452 592 4482 620
rect 4768 591 4798 619
rect 5032 591 5062 619
rect 5348 591 5378 619
rect 5612 591 5642 619
rect 5928 591 5958 619
rect 6192 591 6222 619
rect 6508 591 6538 619
rect 6772 591 6802 619
rect 128 322 158 350
rect 392 322 422 350
rect 708 322 738 350
rect 972 322 1002 350
rect 1288 322 1318 350
rect 1552 322 1582 350
rect 1868 322 1898 350
rect 2132 322 2162 350
rect 2448 322 2478 350
rect 2712 322 2742 350
rect 3028 322 3058 350
rect 3292 322 3322 350
rect 3608 322 3638 350
rect 3872 322 3902 350
rect 4188 322 4218 350
rect 4452 322 4482 350
rect 4768 321 4798 349
rect 5032 321 5062 349
rect 5348 321 5378 349
rect 5612 321 5642 349
rect 5928 321 5958 349
rect 6192 321 6222 349
rect 6508 321 6538 349
rect 6772 321 6802 349
rect 128 52 158 80
rect 392 52 422 80
rect 708 52 738 80
rect 972 52 1002 80
rect 1288 52 1318 80
rect 1552 52 1582 80
rect 1868 52 1898 80
rect 2132 52 2162 80
rect 2448 52 2478 80
rect 2712 52 2742 80
rect 3028 52 3058 80
rect 3292 52 3322 80
rect 3608 52 3638 80
rect 3872 52 3902 80
rect 4188 52 4218 80
rect 4452 52 4482 80
rect 4768 51 4798 79
rect 5032 51 5062 79
rect 5348 51 5378 79
rect 5612 51 5642 79
rect 5928 51 5958 79
rect 6192 51 6222 79
rect 6508 51 6538 79
rect 6772 51 6802 79
rect 128 -218 158 -190
rect 392 -218 422 -190
rect 708 -218 738 -190
rect 972 -218 1002 -190
rect 1288 -218 1318 -190
rect 1552 -218 1582 -190
rect 1868 -218 1898 -190
rect 2132 -218 2162 -190
rect 2448 -218 2478 -190
rect 2712 -218 2742 -190
rect 3028 -218 3058 -190
rect 3292 -218 3322 -190
rect 3608 -218 3638 -190
rect 3872 -218 3902 -190
rect 4188 -218 4218 -190
rect 4452 -218 4482 -190
rect 4768 -219 4798 -191
rect 5032 -219 5062 -191
rect 5348 -219 5378 -191
rect 5612 -219 5642 -191
rect 5928 -219 5958 -191
rect 6192 -219 6222 -191
rect 6508 -219 6538 -191
rect 6772 -219 6802 -191
rect 128 -488 158 -460
rect 392 -488 422 -460
rect 708 -488 738 -460
rect 972 -488 1002 -460
rect 1288 -488 1318 -460
rect 1552 -488 1582 -460
rect 1868 -488 1898 -460
rect 2132 -488 2162 -460
rect 2448 -488 2478 -460
rect 2712 -488 2742 -460
rect 3028 -488 3058 -460
rect 3292 -488 3322 -460
rect 3608 -488 3638 -460
rect 3872 -488 3902 -460
rect 4188 -488 4218 -460
rect 4452 -488 4482 -460
rect 4768 -489 4798 -461
rect 5032 -489 5062 -461
rect 5348 -489 5378 -461
rect 5612 -489 5642 -461
rect 5928 -489 5958 -461
rect 6192 -489 6222 -461
rect 6508 -489 6538 -461
rect 6772 -489 6802 -461
rect 128 -758 158 -730
rect 392 -758 422 -730
rect 708 -758 738 -730
rect 972 -758 1002 -730
rect 1288 -758 1318 -730
rect 1552 -758 1582 -730
rect 1868 -758 1898 -730
rect 2132 -758 2162 -730
rect 2448 -758 2478 -730
rect 2712 -758 2742 -730
rect 3028 -758 3058 -730
rect 3292 -758 3322 -730
rect 3608 -758 3638 -730
rect 3872 -758 3902 -730
rect 4188 -758 4218 -730
rect 4452 -758 4482 -730
rect 4768 -759 4798 -731
rect 5032 -759 5062 -731
rect 5348 -759 5378 -731
rect 5612 -759 5642 -731
rect 5928 -759 5958 -731
rect 6192 -759 6222 -731
rect 6508 -759 6538 -731
rect 6772 -759 6802 -731
rect 128 -1028 158 -1000
rect 392 -1028 422 -1000
rect 708 -1028 738 -1000
rect 972 -1028 1002 -1000
rect 1288 -1028 1318 -1000
rect 1552 -1028 1582 -1000
rect 1868 -1028 1898 -1000
rect 2132 -1028 2162 -1000
rect 2448 -1028 2478 -1000
rect 2712 -1028 2742 -1000
rect 3028 -1028 3058 -1000
rect 3292 -1028 3322 -1000
rect 3608 -1028 3638 -1000
rect 3872 -1028 3902 -1000
rect 4188 -1028 4218 -1000
rect 4452 -1028 4482 -1000
rect 4768 -1029 4798 -1001
rect 5032 -1029 5062 -1001
rect 5348 -1029 5378 -1001
rect 5612 -1029 5642 -1001
rect 5928 -1029 5958 -1001
rect 6192 -1029 6222 -1001
rect 6508 -1029 6538 -1001
rect 6772 -1029 6802 -1001
rect 128 -1298 158 -1270
rect 392 -1298 422 -1270
rect 708 -1298 738 -1270
rect 972 -1298 1002 -1270
rect 1288 -1298 1318 -1270
rect 1552 -1298 1582 -1270
rect 1868 -1298 1898 -1270
rect 2132 -1298 2162 -1270
rect 2448 -1298 2478 -1270
rect 2712 -1298 2742 -1270
rect 3028 -1298 3058 -1270
rect 3292 -1298 3322 -1270
rect 3608 -1298 3638 -1270
rect 3872 -1298 3902 -1270
rect 4188 -1298 4218 -1270
rect 4452 -1298 4482 -1270
rect 4768 -1299 4798 -1271
rect 5032 -1299 5062 -1271
rect 5348 -1299 5378 -1271
rect 5612 -1299 5642 -1271
rect 5928 -1299 5958 -1271
rect 6192 -1299 6222 -1271
rect 6508 -1299 6538 -1271
rect 6772 -1299 6802 -1271
rect 128 -1568 158 -1540
rect 392 -1568 422 -1540
rect 708 -1568 738 -1540
rect 972 -1568 1002 -1540
rect 1288 -1568 1318 -1540
rect 1552 -1568 1582 -1540
rect 1868 -1568 1898 -1540
rect 2132 -1568 2162 -1540
rect 2448 -1568 2478 -1540
rect 2712 -1568 2742 -1540
rect 3028 -1568 3058 -1540
rect 3292 -1568 3322 -1540
rect 3608 -1568 3638 -1540
rect 3872 -1568 3902 -1540
rect 4188 -1568 4218 -1540
rect 4452 -1568 4482 -1540
rect 4768 -1569 4798 -1541
rect 5032 -1569 5062 -1541
rect 5348 -1569 5378 -1541
rect 5612 -1569 5642 -1541
rect 5928 -1569 5958 -1541
rect 6192 -1569 6222 -1541
rect 6508 -1569 6538 -1541
rect 6772 -1569 6802 -1541
rect 128 -1838 158 -1810
rect 392 -1838 422 -1810
rect 708 -1838 738 -1810
rect 972 -1838 1002 -1810
rect 1288 -1838 1318 -1810
rect 1552 -1838 1582 -1810
rect 1868 -1838 1898 -1810
rect 2132 -1838 2162 -1810
rect 2448 -1838 2478 -1810
rect 2712 -1838 2742 -1810
rect 3028 -1838 3058 -1810
rect 3292 -1838 3322 -1810
rect 3608 -1838 3638 -1810
rect 3872 -1838 3902 -1810
rect 4188 -1838 4218 -1810
rect 4452 -1838 4482 -1810
rect 4768 -1839 4798 -1811
rect 5032 -1839 5062 -1811
rect 5348 -1839 5378 -1811
rect 5612 -1839 5642 -1811
rect 5928 -1839 5958 -1811
rect 6192 -1839 6222 -1811
rect 6508 -1839 6538 -1811
rect 6772 -1839 6802 -1811
rect 128 -2108 158 -2080
rect 392 -2108 422 -2080
rect 708 -2108 738 -2080
rect 972 -2108 1002 -2080
rect 1288 -2108 1318 -2080
rect 1552 -2108 1582 -2080
rect 1868 -2108 1898 -2080
rect 2132 -2108 2162 -2080
rect 2448 -2108 2478 -2080
rect 2712 -2108 2742 -2080
rect 3028 -2108 3058 -2080
rect 3292 -2108 3322 -2080
rect 3608 -2108 3638 -2080
rect 3872 -2108 3902 -2080
rect 4188 -2108 4218 -2080
rect 4452 -2108 4482 -2080
rect 4768 -2109 4798 -2081
rect 5032 -2109 5062 -2081
rect 5348 -2109 5378 -2081
rect 5612 -2109 5642 -2081
rect 5928 -2109 5958 -2081
rect 6192 -2109 6222 -2081
rect 6508 -2109 6538 -2081
rect 6772 -2109 6802 -2081
<< ppu >>
rect 221 2078 251 2106
rect 299 2078 329 2106
rect 801 2078 831 2106
rect 879 2078 909 2106
rect 1381 2078 1411 2106
rect 1459 2078 1489 2106
rect 1961 2078 1991 2106
rect 2039 2078 2069 2106
rect 2541 2078 2571 2106
rect 2619 2078 2649 2106
rect 3121 2078 3151 2106
rect 3199 2078 3229 2106
rect 3701 2078 3731 2106
rect 3779 2078 3809 2106
rect 4281 2078 4311 2106
rect 4359 2078 4389 2106
rect 4861 2078 4891 2106
rect 4939 2078 4969 2106
rect 5441 2078 5471 2106
rect 5519 2078 5549 2106
rect 6021 2078 6051 2106
rect 6099 2078 6129 2106
rect 6601 2078 6631 2106
rect 6679 2078 6709 2106
rect 221 1808 251 1836
rect 299 1808 329 1836
rect 801 1808 831 1836
rect 879 1808 909 1836
rect 1381 1808 1411 1836
rect 1459 1808 1489 1836
rect 1961 1808 1991 1836
rect 2039 1808 2069 1836
rect 2541 1808 2571 1836
rect 2619 1808 2649 1836
rect 3121 1808 3151 1836
rect 3199 1808 3229 1836
rect 3701 1808 3731 1836
rect 3779 1808 3809 1836
rect 4281 1808 4311 1836
rect 4359 1808 4389 1836
rect 4861 1808 4891 1836
rect 4939 1808 4969 1836
rect 5441 1808 5471 1836
rect 5519 1808 5549 1836
rect 6021 1808 6051 1836
rect 6099 1808 6129 1836
rect 6601 1808 6631 1836
rect 6679 1808 6709 1836
rect 221 1538 251 1566
rect 299 1538 329 1566
rect 801 1538 831 1566
rect 879 1538 909 1566
rect 1381 1538 1411 1566
rect 1459 1538 1489 1566
rect 1961 1538 1991 1566
rect 2039 1538 2069 1566
rect 2541 1538 2571 1566
rect 2619 1538 2649 1566
rect 3121 1538 3151 1566
rect 3199 1538 3229 1566
rect 3701 1538 3731 1566
rect 3779 1538 3809 1566
rect 4281 1538 4311 1566
rect 4359 1538 4389 1566
rect 4861 1538 4891 1566
rect 4939 1538 4969 1566
rect 5441 1538 5471 1566
rect 5519 1538 5549 1566
rect 6021 1538 6051 1566
rect 6099 1538 6129 1566
rect 6601 1538 6631 1566
rect 6679 1538 6709 1566
rect 221 1268 251 1296
rect 299 1268 329 1296
rect 801 1268 831 1296
rect 879 1268 909 1296
rect 1381 1268 1411 1296
rect 1459 1268 1489 1296
rect 1961 1268 1991 1296
rect 2039 1268 2069 1296
rect 2541 1268 2571 1296
rect 2619 1268 2649 1296
rect 3121 1268 3151 1296
rect 3199 1268 3229 1296
rect 3701 1268 3731 1296
rect 3779 1268 3809 1296
rect 4281 1268 4311 1296
rect 4359 1268 4389 1296
rect 4861 1268 4891 1296
rect 4939 1268 4969 1296
rect 5441 1268 5471 1296
rect 5519 1268 5549 1296
rect 6021 1268 6051 1296
rect 6099 1268 6129 1296
rect 6601 1268 6631 1296
rect 6679 1268 6709 1296
rect 221 998 251 1026
rect 299 998 329 1026
rect 801 998 831 1026
rect 879 998 909 1026
rect 1381 998 1411 1026
rect 1459 998 1489 1026
rect 1961 998 1991 1026
rect 2039 998 2069 1026
rect 2541 998 2571 1026
rect 2619 998 2649 1026
rect 3121 998 3151 1026
rect 3199 998 3229 1026
rect 3701 998 3731 1026
rect 3779 998 3809 1026
rect 4281 998 4311 1026
rect 4359 998 4389 1026
rect 4861 997 4891 1025
rect 4939 997 4969 1025
rect 5441 997 5471 1025
rect 5519 997 5549 1025
rect 6021 997 6051 1025
rect 6099 997 6129 1025
rect 6601 997 6631 1025
rect 6679 997 6709 1025
rect 221 728 251 756
rect 299 728 329 756
rect 801 728 831 756
rect 879 728 909 756
rect 1381 728 1411 756
rect 1459 728 1489 756
rect 1961 728 1991 756
rect 2039 728 2069 756
rect 2541 728 2571 756
rect 2619 728 2649 756
rect 3121 728 3151 756
rect 3199 728 3229 756
rect 3701 728 3731 756
rect 3779 728 3809 756
rect 4281 728 4311 756
rect 4359 728 4389 756
rect 4861 727 4891 755
rect 4939 727 4969 755
rect 5441 727 5471 755
rect 5519 727 5549 755
rect 6021 727 6051 755
rect 6099 727 6129 755
rect 6601 727 6631 755
rect 6679 727 6709 755
rect 221 458 251 486
rect 299 458 329 486
rect 801 458 831 486
rect 879 458 909 486
rect 1381 458 1411 486
rect 1459 458 1489 486
rect 1961 458 1991 486
rect 2039 458 2069 486
rect 2541 458 2571 486
rect 2619 458 2649 486
rect 3121 458 3151 486
rect 3199 458 3229 486
rect 3701 458 3731 486
rect 3779 458 3809 486
rect 4281 458 4311 486
rect 4359 458 4389 486
rect 4861 457 4891 485
rect 4939 457 4969 485
rect 5441 457 5471 485
rect 5519 457 5549 485
rect 6021 457 6051 485
rect 6099 457 6129 485
rect 6601 457 6631 485
rect 6679 457 6709 485
rect 221 188 251 216
rect 299 188 329 216
rect 801 188 831 216
rect 879 188 909 216
rect 1381 188 1411 216
rect 1459 188 1489 216
rect 1961 188 1991 216
rect 2039 188 2069 216
rect 2541 188 2571 216
rect 2619 188 2649 216
rect 3121 188 3151 216
rect 3199 188 3229 216
rect 3701 188 3731 216
rect 3779 188 3809 216
rect 4281 188 4311 216
rect 4359 188 4389 216
rect 4861 187 4891 215
rect 4939 187 4969 215
rect 5441 187 5471 215
rect 5519 187 5549 215
rect 6021 187 6051 215
rect 6099 187 6129 215
rect 6601 187 6631 215
rect 6679 187 6709 215
rect 221 -82 251 -54
rect 299 -82 329 -54
rect 801 -82 831 -54
rect 879 -82 909 -54
rect 1381 -82 1411 -54
rect 1459 -82 1489 -54
rect 1961 -82 1991 -54
rect 2039 -82 2069 -54
rect 2541 -82 2571 -54
rect 2619 -82 2649 -54
rect 3121 -82 3151 -54
rect 3199 -82 3229 -54
rect 3701 -82 3731 -54
rect 3779 -82 3809 -54
rect 4281 -82 4311 -54
rect 4359 -82 4389 -54
rect 4861 -83 4891 -55
rect 4939 -83 4969 -55
rect 5441 -83 5471 -55
rect 5519 -83 5549 -55
rect 6021 -83 6051 -55
rect 6099 -83 6129 -55
rect 6601 -83 6631 -55
rect 6679 -83 6709 -55
rect 221 -352 251 -324
rect 299 -352 329 -324
rect 801 -352 831 -324
rect 879 -352 909 -324
rect 1381 -352 1411 -324
rect 1459 -352 1489 -324
rect 1961 -352 1991 -324
rect 2039 -352 2069 -324
rect 2541 -352 2571 -324
rect 2619 -352 2649 -324
rect 3121 -352 3151 -324
rect 3199 -352 3229 -324
rect 3701 -352 3731 -324
rect 3779 -352 3809 -324
rect 4281 -352 4311 -324
rect 4359 -352 4389 -324
rect 4861 -353 4891 -325
rect 4939 -353 4969 -325
rect 5441 -353 5471 -325
rect 5519 -353 5549 -325
rect 6021 -353 6051 -325
rect 6099 -353 6129 -325
rect 6601 -353 6631 -325
rect 6679 -353 6709 -325
rect 221 -622 251 -594
rect 299 -622 329 -594
rect 801 -622 831 -594
rect 879 -622 909 -594
rect 1381 -622 1411 -594
rect 1459 -622 1489 -594
rect 1961 -622 1991 -594
rect 2039 -622 2069 -594
rect 2541 -622 2571 -594
rect 2619 -622 2649 -594
rect 3121 -622 3151 -594
rect 3199 -622 3229 -594
rect 3701 -622 3731 -594
rect 3779 -622 3809 -594
rect 4281 -622 4311 -594
rect 4359 -622 4389 -594
rect 4861 -623 4891 -595
rect 4939 -623 4969 -595
rect 5441 -623 5471 -595
rect 5519 -623 5549 -595
rect 6021 -623 6051 -595
rect 6099 -623 6129 -595
rect 6601 -623 6631 -595
rect 6679 -623 6709 -595
rect 221 -892 251 -864
rect 299 -892 329 -864
rect 801 -892 831 -864
rect 879 -892 909 -864
rect 1381 -892 1411 -864
rect 1459 -892 1489 -864
rect 1961 -892 1991 -864
rect 2039 -892 2069 -864
rect 2541 -892 2571 -864
rect 2619 -892 2649 -864
rect 3121 -892 3151 -864
rect 3199 -892 3229 -864
rect 3701 -892 3731 -864
rect 3779 -892 3809 -864
rect 4281 -892 4311 -864
rect 4359 -892 4389 -864
rect 4861 -893 4891 -865
rect 4939 -893 4969 -865
rect 5441 -893 5471 -865
rect 5519 -893 5549 -865
rect 6021 -893 6051 -865
rect 6099 -893 6129 -865
rect 6601 -893 6631 -865
rect 6679 -893 6709 -865
rect 221 -1162 251 -1134
rect 299 -1162 329 -1134
rect 801 -1162 831 -1134
rect 879 -1162 909 -1134
rect 1381 -1162 1411 -1134
rect 1459 -1162 1489 -1134
rect 1961 -1162 1991 -1134
rect 2039 -1162 2069 -1134
rect 2541 -1162 2571 -1134
rect 2619 -1162 2649 -1134
rect 3121 -1162 3151 -1134
rect 3199 -1162 3229 -1134
rect 3701 -1162 3731 -1134
rect 3779 -1162 3809 -1134
rect 4281 -1162 4311 -1134
rect 4359 -1162 4389 -1134
rect 4861 -1163 4891 -1135
rect 4939 -1163 4969 -1135
rect 5441 -1163 5471 -1135
rect 5519 -1163 5549 -1135
rect 6021 -1163 6051 -1135
rect 6099 -1163 6129 -1135
rect 6601 -1163 6631 -1135
rect 6679 -1163 6709 -1135
rect 221 -1432 251 -1404
rect 299 -1432 329 -1404
rect 801 -1432 831 -1404
rect 879 -1432 909 -1404
rect 1381 -1432 1411 -1404
rect 1459 -1432 1489 -1404
rect 1961 -1432 1991 -1404
rect 2039 -1432 2069 -1404
rect 2541 -1432 2571 -1404
rect 2619 -1432 2649 -1404
rect 3121 -1432 3151 -1404
rect 3199 -1432 3229 -1404
rect 3701 -1432 3731 -1404
rect 3779 -1432 3809 -1404
rect 4281 -1432 4311 -1404
rect 4359 -1432 4389 -1404
rect 4861 -1433 4891 -1405
rect 4939 -1433 4969 -1405
rect 5441 -1433 5471 -1405
rect 5519 -1433 5549 -1405
rect 6021 -1433 6051 -1405
rect 6099 -1433 6129 -1405
rect 6601 -1433 6631 -1405
rect 6679 -1433 6709 -1405
rect 221 -1702 251 -1674
rect 299 -1702 329 -1674
rect 801 -1702 831 -1674
rect 879 -1702 909 -1674
rect 1381 -1702 1411 -1674
rect 1459 -1702 1489 -1674
rect 1961 -1702 1991 -1674
rect 2039 -1702 2069 -1674
rect 2541 -1702 2571 -1674
rect 2619 -1702 2649 -1674
rect 3121 -1702 3151 -1674
rect 3199 -1702 3229 -1674
rect 3701 -1702 3731 -1674
rect 3779 -1702 3809 -1674
rect 4281 -1702 4311 -1674
rect 4359 -1702 4389 -1674
rect 4861 -1703 4891 -1675
rect 4939 -1703 4969 -1675
rect 5441 -1703 5471 -1675
rect 5519 -1703 5549 -1675
rect 6021 -1703 6051 -1675
rect 6099 -1703 6129 -1675
rect 6601 -1703 6631 -1675
rect 6679 -1703 6709 -1675
rect 221 -1972 251 -1944
rect 299 -1972 329 -1944
rect 801 -1972 831 -1944
rect 879 -1972 909 -1944
rect 1381 -1972 1411 -1944
rect 1459 -1972 1489 -1944
rect 1961 -1972 1991 -1944
rect 2039 -1972 2069 -1944
rect 2541 -1972 2571 -1944
rect 2619 -1972 2649 -1944
rect 3121 -1972 3151 -1944
rect 3199 -1972 3229 -1944
rect 3701 -1972 3731 -1944
rect 3779 -1972 3809 -1944
rect 4281 -1972 4311 -1944
rect 4359 -1972 4389 -1944
rect 4861 -1973 4891 -1945
rect 4939 -1973 4969 -1945
rect 5441 -1973 5471 -1945
rect 5519 -1973 5549 -1945
rect 6021 -1973 6051 -1945
rect 6099 -1973 6129 -1945
rect 6601 -1973 6631 -1945
rect 6679 -1973 6709 -1945
<< ndiff >>
rect 88 2088 106 2116
rect 136 2088 154 2116
rect 396 2088 414 2116
rect 444 2088 463 2116
rect 668 2088 686 2116
rect 716 2088 734 2116
rect 976 2088 994 2116
rect 1024 2088 1043 2116
rect 1248 2088 1266 2116
rect 1296 2088 1314 2116
rect 1556 2088 1574 2116
rect 1604 2088 1623 2116
rect 1828 2088 1846 2116
rect 1876 2088 1894 2116
rect 2136 2088 2154 2116
rect 2184 2088 2203 2116
rect 2408 2088 2426 2116
rect 2456 2088 2474 2116
rect 2716 2088 2734 2116
rect 2764 2088 2783 2116
rect 2988 2088 3006 2116
rect 3036 2088 3054 2116
rect 3296 2088 3314 2116
rect 3344 2088 3363 2116
rect 3568 2088 3586 2116
rect 3616 2088 3634 2116
rect 3876 2088 3894 2116
rect 3924 2088 3943 2116
rect 4148 2088 4166 2116
rect 4196 2088 4214 2116
rect 4456 2088 4474 2116
rect 4504 2088 4523 2116
rect 4728 2088 4746 2116
rect 4776 2088 4794 2116
rect 5036 2088 5054 2116
rect 5084 2088 5103 2116
rect 5308 2088 5326 2116
rect 5356 2088 5374 2116
rect 5616 2088 5634 2116
rect 5664 2088 5683 2116
rect 5888 2088 5906 2116
rect 5936 2088 5954 2116
rect 6196 2088 6214 2116
rect 6244 2088 6263 2116
rect 6468 2088 6486 2116
rect 6516 2088 6534 2116
rect 6776 2088 6794 2116
rect 6824 2088 6843 2116
rect 14 1942 42 1984
rect 72 1970 97 1984
rect 196 1974 221 1984
rect 72 1942 128 1970
rect 158 1942 192 1970
tri 206 1967 213 1974 ne
rect 213 1942 221 1974
rect 251 1942 299 1984
rect 329 1974 354 1984
rect 329 1942 337 1974
rect 453 1970 478 1984
rect 358 1942 392 1970
rect 422 1942 478 1970
rect 508 1942 536 1984
rect 594 1942 622 1984
rect 652 1970 677 1984
rect 776 1974 801 1984
rect 652 1942 708 1970
rect 738 1942 772 1970
tri 786 1967 793 1974 ne
rect 793 1942 801 1974
rect 831 1942 879 1984
rect 909 1974 934 1984
rect 909 1942 917 1974
rect 1033 1970 1058 1984
rect 938 1942 972 1970
rect 1002 1942 1058 1970
rect 1088 1942 1116 1984
rect 1174 1942 1202 1984
rect 1232 1970 1257 1984
rect 1356 1974 1381 1984
rect 1232 1942 1288 1970
rect 1318 1942 1352 1970
tri 1366 1967 1373 1974 ne
rect 1373 1942 1381 1974
rect 1411 1942 1459 1984
rect 1489 1974 1514 1984
rect 1489 1942 1497 1974
rect 1613 1970 1638 1984
rect 1518 1942 1552 1970
rect 1582 1942 1638 1970
rect 1668 1942 1696 1984
rect 1754 1942 1782 1984
rect 1812 1970 1837 1984
rect 1936 1974 1961 1984
rect 1812 1942 1868 1970
rect 1898 1942 1932 1970
tri 1946 1967 1953 1974 ne
rect 1953 1942 1961 1974
rect 1991 1942 2039 1984
rect 2069 1974 2094 1984
rect 2069 1942 2077 1974
rect 2193 1970 2218 1984
rect 2098 1942 2132 1970
rect 2162 1942 2218 1970
rect 2248 1942 2276 1984
rect 2334 1942 2362 1984
rect 2392 1970 2417 1984
rect 2516 1974 2541 1984
rect 2392 1942 2448 1970
rect 2478 1942 2512 1970
tri 2526 1967 2533 1974 ne
rect 2533 1942 2541 1974
rect 2571 1942 2619 1984
rect 2649 1974 2674 1984
rect 2649 1942 2657 1974
rect 2773 1970 2798 1984
rect 2678 1942 2712 1970
rect 2742 1942 2798 1970
rect 2828 1942 2856 1984
rect 2914 1942 2942 1984
rect 2972 1970 2997 1984
rect 3096 1974 3121 1984
rect 2972 1942 3028 1970
rect 3058 1942 3092 1970
tri 3106 1967 3113 1974 ne
rect 3113 1942 3121 1974
rect 3151 1942 3199 1984
rect 3229 1974 3254 1984
rect 3229 1942 3237 1974
rect 3353 1970 3378 1984
rect 3258 1942 3292 1970
rect 3322 1942 3378 1970
rect 3408 1942 3436 1984
rect 3494 1942 3522 1984
rect 3552 1970 3577 1984
rect 3676 1974 3701 1984
rect 3552 1942 3608 1970
rect 3638 1942 3672 1970
tri 3686 1967 3693 1974 ne
rect 3693 1942 3701 1974
rect 3731 1942 3779 1984
rect 3809 1974 3834 1984
rect 3809 1942 3817 1974
rect 3933 1970 3958 1984
rect 3838 1942 3872 1970
rect 3902 1942 3958 1970
rect 3988 1942 4016 1984
rect 4074 1942 4102 1984
rect 4132 1970 4157 1984
rect 4256 1974 4281 1984
rect 4132 1942 4188 1970
rect 4218 1942 4252 1970
tri 4266 1967 4273 1974 ne
rect 4273 1942 4281 1974
rect 4311 1942 4359 1984
rect 4389 1974 4414 1984
rect 4389 1942 4397 1974
rect 4513 1970 4538 1984
rect 4418 1942 4452 1970
rect 4482 1942 4538 1970
rect 4568 1942 4596 1984
rect 4654 1942 4682 1984
rect 4712 1970 4737 1984
rect 4836 1974 4861 1984
rect 4712 1942 4768 1970
rect 4798 1942 4832 1970
tri 4846 1967 4853 1974 ne
rect 4853 1942 4861 1974
rect 4891 1942 4939 1984
rect 4969 1974 4994 1984
rect 4969 1942 4977 1974
rect 5093 1970 5118 1984
rect 4998 1942 5032 1970
rect 5062 1942 5118 1970
rect 5148 1942 5176 1984
rect 5234 1942 5262 1984
rect 5292 1970 5317 1984
rect 5416 1974 5441 1984
rect 5292 1942 5348 1970
rect 5378 1942 5412 1970
tri 5426 1967 5433 1974 ne
rect 5433 1942 5441 1974
rect 5471 1942 5519 1984
rect 5549 1974 5574 1984
rect 5549 1942 5557 1974
rect 5673 1970 5698 1984
rect 5578 1942 5612 1970
rect 5642 1942 5698 1970
rect 5728 1942 5756 1984
rect 5814 1942 5842 1984
rect 5872 1970 5897 1984
rect 5996 1974 6021 1984
rect 5872 1942 5928 1970
rect 5958 1942 5992 1970
tri 6006 1967 6013 1974 ne
rect 6013 1942 6021 1974
rect 6051 1942 6099 1984
rect 6129 1974 6154 1984
rect 6129 1942 6137 1974
rect 6253 1970 6278 1984
rect 6158 1942 6192 1970
rect 6222 1942 6278 1970
rect 6308 1942 6336 1984
rect 6394 1942 6422 1984
rect 6452 1970 6477 1984
rect 6576 1974 6601 1984
rect 6452 1942 6508 1970
rect 6538 1942 6572 1970
tri 6586 1967 6593 1974 ne
rect 6593 1942 6601 1974
rect 6631 1942 6679 1984
rect 6709 1974 6734 1984
rect 6709 1942 6717 1974
rect 6833 1970 6858 1984
rect 6738 1942 6772 1970
rect 6802 1942 6858 1970
rect 6888 1942 6916 1984
rect 165 1918 192 1942
rect 259 1920 291 1942
rect 259 1918 261 1920
rect 289 1918 291 1920
rect 358 1918 385 1942
rect 165 1904 259 1918
rect 291 1904 385 1918
rect 745 1918 772 1942
rect 839 1920 871 1942
rect 839 1918 841 1920
rect 869 1918 871 1920
rect 938 1918 965 1942
rect 745 1904 839 1918
rect 871 1904 965 1918
rect 1325 1918 1352 1942
rect 1419 1920 1451 1942
rect 1419 1918 1421 1920
rect 1449 1918 1451 1920
rect 1518 1918 1545 1942
rect 1325 1904 1419 1918
rect 1451 1904 1545 1918
rect 1905 1918 1932 1942
rect 1999 1920 2031 1942
rect 1999 1918 2001 1920
rect 2029 1918 2031 1920
rect 2098 1918 2125 1942
rect 1905 1904 1999 1918
rect 2031 1904 2125 1918
rect 2485 1918 2512 1942
rect 2579 1920 2611 1942
rect 2579 1918 2581 1920
rect 2609 1918 2611 1920
rect 2678 1918 2705 1942
rect 2485 1904 2579 1918
rect 2611 1904 2705 1918
rect 3065 1918 3092 1942
rect 3159 1920 3191 1942
rect 3159 1918 3161 1920
rect 3189 1918 3191 1920
rect 3258 1918 3285 1942
rect 3065 1904 3159 1918
rect 3191 1904 3285 1918
rect 3645 1918 3672 1942
rect 3739 1920 3771 1942
rect 3739 1918 3741 1920
rect 3769 1918 3771 1920
rect 3838 1918 3865 1942
rect 3645 1904 3739 1918
rect 3771 1904 3865 1918
rect 4225 1918 4252 1942
rect 4319 1920 4351 1942
rect 4319 1918 4321 1920
rect 4349 1918 4351 1920
rect 4418 1918 4445 1942
rect 4225 1904 4319 1918
rect 4351 1904 4445 1918
rect 4805 1918 4832 1942
rect 4899 1920 4931 1942
rect 4899 1918 4901 1920
rect 4929 1918 4931 1920
rect 4998 1918 5025 1942
rect 4805 1904 4899 1918
rect 4931 1904 5025 1918
rect 5385 1918 5412 1942
rect 5479 1920 5511 1942
rect 5479 1918 5481 1920
rect 5509 1918 5511 1920
rect 5578 1918 5605 1942
rect 5385 1904 5479 1918
rect 5511 1904 5605 1918
rect 5965 1918 5992 1942
rect 6059 1920 6091 1942
rect 6059 1918 6061 1920
rect 6089 1918 6091 1920
rect 6158 1918 6185 1942
rect 5965 1904 6059 1918
rect 6091 1904 6185 1918
rect 6545 1918 6572 1942
rect 6639 1920 6671 1942
rect 6639 1918 6641 1920
rect 6669 1918 6671 1920
rect 6738 1918 6765 1942
rect 6545 1904 6639 1918
rect 6671 1904 6765 1918
rect 88 1818 106 1846
rect 136 1818 154 1846
rect 396 1818 414 1846
rect 444 1818 463 1846
rect 668 1818 686 1846
rect 716 1818 734 1846
rect 976 1818 994 1846
rect 1024 1818 1043 1846
rect 1248 1818 1266 1846
rect 1296 1818 1314 1846
rect 1556 1818 1574 1846
rect 1604 1818 1623 1846
rect 1828 1818 1846 1846
rect 1876 1818 1894 1846
rect 2136 1818 2154 1846
rect 2184 1818 2203 1846
rect 2408 1818 2426 1846
rect 2456 1818 2474 1846
rect 2716 1818 2734 1846
rect 2764 1818 2783 1846
rect 2988 1818 3006 1846
rect 3036 1818 3054 1846
rect 3296 1818 3314 1846
rect 3344 1818 3363 1846
rect 3568 1818 3586 1846
rect 3616 1818 3634 1846
rect 3876 1818 3894 1846
rect 3924 1818 3943 1846
rect 4148 1818 4166 1846
rect 4196 1818 4214 1846
rect 4456 1818 4474 1846
rect 4504 1818 4523 1846
rect 4728 1818 4746 1846
rect 4776 1818 4794 1846
rect 5036 1818 5054 1846
rect 5084 1818 5103 1846
rect 5308 1818 5326 1846
rect 5356 1818 5374 1846
rect 5616 1818 5634 1846
rect 5664 1818 5683 1846
rect 5888 1818 5906 1846
rect 5936 1818 5954 1846
rect 6196 1818 6214 1846
rect 6244 1818 6263 1846
rect 6468 1818 6486 1846
rect 6516 1818 6534 1846
rect 6776 1818 6794 1846
rect 6824 1818 6843 1846
rect 14 1672 42 1714
rect 72 1700 97 1714
rect 196 1704 221 1714
rect 72 1672 128 1700
rect 158 1672 192 1700
tri 206 1697 213 1704 ne
rect 213 1672 221 1704
rect 251 1672 299 1714
rect 329 1704 354 1714
rect 329 1672 337 1704
rect 453 1700 478 1714
rect 358 1672 392 1700
rect 422 1672 478 1700
rect 508 1672 536 1714
rect 594 1672 622 1714
rect 652 1700 677 1714
rect 776 1704 801 1714
rect 652 1672 708 1700
rect 738 1672 772 1700
tri 786 1697 793 1704 ne
rect 793 1672 801 1704
rect 831 1672 879 1714
rect 909 1704 934 1714
rect 909 1672 917 1704
rect 1033 1700 1058 1714
rect 938 1672 972 1700
rect 1002 1672 1058 1700
rect 1088 1672 1116 1714
rect 1174 1672 1202 1714
rect 1232 1700 1257 1714
rect 1356 1704 1381 1714
rect 1232 1672 1288 1700
rect 1318 1672 1352 1700
tri 1366 1697 1373 1704 ne
rect 1373 1672 1381 1704
rect 1411 1672 1459 1714
rect 1489 1704 1514 1714
rect 1489 1672 1497 1704
rect 1613 1700 1638 1714
rect 1518 1672 1552 1700
rect 1582 1672 1638 1700
rect 1668 1672 1696 1714
rect 1754 1672 1782 1714
rect 1812 1700 1837 1714
rect 1936 1704 1961 1714
rect 1812 1672 1868 1700
rect 1898 1672 1932 1700
tri 1946 1697 1953 1704 ne
rect 1953 1672 1961 1704
rect 1991 1672 2039 1714
rect 2069 1704 2094 1714
rect 2069 1672 2077 1704
rect 2193 1700 2218 1714
rect 2098 1672 2132 1700
rect 2162 1672 2218 1700
rect 2248 1672 2276 1714
rect 2334 1672 2362 1714
rect 2392 1700 2417 1714
rect 2516 1704 2541 1714
rect 2392 1672 2448 1700
rect 2478 1672 2512 1700
tri 2526 1697 2533 1704 ne
rect 2533 1672 2541 1704
rect 2571 1672 2619 1714
rect 2649 1704 2674 1714
rect 2649 1672 2657 1704
rect 2773 1700 2798 1714
rect 2678 1672 2712 1700
rect 2742 1672 2798 1700
rect 2828 1672 2856 1714
rect 2914 1672 2942 1714
rect 2972 1700 2997 1714
rect 3096 1704 3121 1714
rect 2972 1672 3028 1700
rect 3058 1672 3092 1700
tri 3106 1697 3113 1704 ne
rect 3113 1672 3121 1704
rect 3151 1672 3199 1714
rect 3229 1704 3254 1714
rect 3229 1672 3237 1704
rect 3353 1700 3378 1714
rect 3258 1672 3292 1700
rect 3322 1672 3378 1700
rect 3408 1672 3436 1714
rect 3494 1672 3522 1714
rect 3552 1700 3577 1714
rect 3676 1704 3701 1714
rect 3552 1672 3608 1700
rect 3638 1672 3672 1700
tri 3686 1697 3693 1704 ne
rect 3693 1672 3701 1704
rect 3731 1672 3779 1714
rect 3809 1704 3834 1714
rect 3809 1672 3817 1704
rect 3933 1700 3958 1714
rect 3838 1672 3872 1700
rect 3902 1672 3958 1700
rect 3988 1672 4016 1714
rect 4074 1672 4102 1714
rect 4132 1700 4157 1714
rect 4256 1704 4281 1714
rect 4132 1672 4188 1700
rect 4218 1672 4252 1700
tri 4266 1697 4273 1704 ne
rect 4273 1672 4281 1704
rect 4311 1672 4359 1714
rect 4389 1704 4414 1714
rect 4389 1672 4397 1704
rect 4513 1700 4538 1714
rect 4418 1672 4452 1700
rect 4482 1672 4538 1700
rect 4568 1672 4596 1714
rect 4654 1672 4682 1714
rect 4712 1700 4737 1714
rect 4836 1704 4861 1714
rect 4712 1672 4768 1700
rect 4798 1672 4832 1700
tri 4846 1697 4853 1704 ne
rect 4853 1672 4861 1704
rect 4891 1672 4939 1714
rect 4969 1704 4994 1714
rect 4969 1672 4977 1704
rect 5093 1700 5118 1714
rect 4998 1672 5032 1700
rect 5062 1672 5118 1700
rect 5148 1672 5176 1714
rect 5234 1672 5262 1714
rect 5292 1700 5317 1714
rect 5416 1704 5441 1714
rect 5292 1672 5348 1700
rect 5378 1672 5412 1700
tri 5426 1697 5433 1704 ne
rect 5433 1672 5441 1704
rect 5471 1672 5519 1714
rect 5549 1704 5574 1714
rect 5549 1672 5557 1704
rect 5673 1700 5698 1714
rect 5578 1672 5612 1700
rect 5642 1672 5698 1700
rect 5728 1672 5756 1714
rect 5814 1672 5842 1714
rect 5872 1700 5897 1714
rect 5996 1704 6021 1714
rect 5872 1672 5928 1700
rect 5958 1672 5992 1700
tri 6006 1697 6013 1704 ne
rect 6013 1672 6021 1704
rect 6051 1672 6099 1714
rect 6129 1704 6154 1714
rect 6129 1672 6137 1704
rect 6253 1700 6278 1714
rect 6158 1672 6192 1700
rect 6222 1672 6278 1700
rect 6308 1672 6336 1714
rect 6394 1672 6422 1714
rect 6452 1700 6477 1714
rect 6576 1704 6601 1714
rect 6452 1672 6508 1700
rect 6538 1672 6572 1700
tri 6586 1697 6593 1704 ne
rect 6593 1672 6601 1704
rect 6631 1672 6679 1714
rect 6709 1704 6734 1714
rect 6709 1672 6717 1704
rect 6833 1700 6858 1714
rect 6738 1672 6772 1700
rect 6802 1672 6858 1700
rect 6888 1672 6916 1714
rect 165 1648 192 1672
rect 259 1650 291 1672
rect 259 1648 261 1650
rect 289 1648 291 1650
rect 358 1648 385 1672
rect 165 1634 259 1648
rect 291 1634 385 1648
rect 745 1648 772 1672
rect 839 1650 871 1672
rect 839 1648 841 1650
rect 869 1648 871 1650
rect 938 1648 965 1672
rect 745 1634 839 1648
rect 871 1634 965 1648
rect 1325 1648 1352 1672
rect 1419 1650 1451 1672
rect 1419 1648 1421 1650
rect 1449 1648 1451 1650
rect 1518 1648 1545 1672
rect 1325 1634 1419 1648
rect 1451 1634 1545 1648
rect 1905 1648 1932 1672
rect 1999 1650 2031 1672
rect 1999 1648 2001 1650
rect 2029 1648 2031 1650
rect 2098 1648 2125 1672
rect 1905 1634 1999 1648
rect 2031 1634 2125 1648
rect 2485 1648 2512 1672
rect 2579 1650 2611 1672
rect 2579 1648 2581 1650
rect 2609 1648 2611 1650
rect 2678 1648 2705 1672
rect 2485 1634 2579 1648
rect 2611 1634 2705 1648
rect 3065 1648 3092 1672
rect 3159 1650 3191 1672
rect 3159 1648 3161 1650
rect 3189 1648 3191 1650
rect 3258 1648 3285 1672
rect 3065 1634 3159 1648
rect 3191 1634 3285 1648
rect 3645 1648 3672 1672
rect 3739 1650 3771 1672
rect 3739 1648 3741 1650
rect 3769 1648 3771 1650
rect 3838 1648 3865 1672
rect 3645 1634 3739 1648
rect 3771 1634 3865 1648
rect 4225 1648 4252 1672
rect 4319 1650 4351 1672
rect 4319 1648 4321 1650
rect 4349 1648 4351 1650
rect 4418 1648 4445 1672
rect 4225 1634 4319 1648
rect 4351 1634 4445 1648
rect 4805 1648 4832 1672
rect 4899 1650 4931 1672
rect 4899 1648 4901 1650
rect 4929 1648 4931 1650
rect 4998 1648 5025 1672
rect 4805 1634 4899 1648
rect 4931 1634 5025 1648
rect 5385 1648 5412 1672
rect 5479 1650 5511 1672
rect 5479 1648 5481 1650
rect 5509 1648 5511 1650
rect 5578 1648 5605 1672
rect 5385 1634 5479 1648
rect 5511 1634 5605 1648
rect 5965 1648 5992 1672
rect 6059 1650 6091 1672
rect 6059 1648 6061 1650
rect 6089 1648 6091 1650
rect 6158 1648 6185 1672
rect 5965 1634 6059 1648
rect 6091 1634 6185 1648
rect 6545 1648 6572 1672
rect 6639 1650 6671 1672
rect 6639 1648 6641 1650
rect 6669 1648 6671 1650
rect 6738 1648 6765 1672
rect 6545 1634 6639 1648
rect 6671 1634 6765 1648
rect 88 1548 106 1576
rect 136 1548 154 1576
rect 396 1548 414 1576
rect 444 1548 463 1576
rect 668 1548 686 1576
rect 716 1548 734 1576
rect 976 1548 994 1576
rect 1024 1548 1043 1576
rect 1248 1548 1266 1576
rect 1296 1548 1314 1576
rect 1556 1548 1574 1576
rect 1604 1548 1623 1576
rect 1828 1548 1846 1576
rect 1876 1548 1894 1576
rect 2136 1548 2154 1576
rect 2184 1548 2203 1576
rect 2408 1548 2426 1576
rect 2456 1548 2474 1576
rect 2716 1548 2734 1576
rect 2764 1548 2783 1576
rect 2988 1548 3006 1576
rect 3036 1548 3054 1576
rect 3296 1548 3314 1576
rect 3344 1548 3363 1576
rect 3568 1548 3586 1576
rect 3616 1548 3634 1576
rect 3876 1548 3894 1576
rect 3924 1548 3943 1576
rect 4148 1548 4166 1576
rect 4196 1548 4214 1576
rect 4456 1548 4474 1576
rect 4504 1548 4523 1576
rect 4728 1548 4746 1576
rect 4776 1548 4794 1576
rect 5036 1548 5054 1576
rect 5084 1548 5103 1576
rect 5308 1548 5326 1576
rect 5356 1548 5374 1576
rect 5616 1548 5634 1576
rect 5664 1548 5683 1576
rect 5888 1548 5906 1576
rect 5936 1548 5954 1576
rect 6196 1548 6214 1576
rect 6244 1548 6263 1576
rect 6468 1548 6486 1576
rect 6516 1548 6534 1576
rect 6776 1548 6794 1576
rect 6824 1548 6843 1576
rect 14 1402 42 1444
rect 72 1430 97 1444
rect 196 1434 221 1444
rect 72 1402 128 1430
rect 158 1402 192 1430
tri 206 1427 213 1434 ne
rect 213 1402 221 1434
rect 251 1402 299 1444
rect 329 1434 354 1444
rect 329 1402 337 1434
rect 453 1430 478 1444
rect 358 1402 392 1430
rect 422 1402 478 1430
rect 508 1402 536 1444
rect 594 1402 622 1444
rect 652 1430 677 1444
rect 776 1434 801 1444
rect 652 1402 708 1430
rect 738 1402 772 1430
tri 786 1427 793 1434 ne
rect 793 1402 801 1434
rect 831 1402 879 1444
rect 909 1434 934 1444
rect 909 1402 917 1434
rect 1033 1430 1058 1444
rect 938 1402 972 1430
rect 1002 1402 1058 1430
rect 1088 1402 1116 1444
rect 1174 1402 1202 1444
rect 1232 1430 1257 1444
rect 1356 1434 1381 1444
rect 1232 1402 1288 1430
rect 1318 1402 1352 1430
tri 1366 1427 1373 1434 ne
rect 1373 1402 1381 1434
rect 1411 1402 1459 1444
rect 1489 1434 1514 1444
rect 1489 1402 1497 1434
rect 1613 1430 1638 1444
rect 1518 1402 1552 1430
rect 1582 1402 1638 1430
rect 1668 1402 1696 1444
rect 1754 1402 1782 1444
rect 1812 1430 1837 1444
rect 1936 1434 1961 1444
rect 1812 1402 1868 1430
rect 1898 1402 1932 1430
tri 1946 1427 1953 1434 ne
rect 1953 1402 1961 1434
rect 1991 1402 2039 1444
rect 2069 1434 2094 1444
rect 2069 1402 2077 1434
rect 2193 1430 2218 1444
rect 2098 1402 2132 1430
rect 2162 1402 2218 1430
rect 2248 1402 2276 1444
rect 2334 1402 2362 1444
rect 2392 1430 2417 1444
rect 2516 1434 2541 1444
rect 2392 1402 2448 1430
rect 2478 1402 2512 1430
tri 2526 1427 2533 1434 ne
rect 2533 1402 2541 1434
rect 2571 1402 2619 1444
rect 2649 1434 2674 1444
rect 2649 1402 2657 1434
rect 2773 1430 2798 1444
rect 2678 1402 2712 1430
rect 2742 1402 2798 1430
rect 2828 1402 2856 1444
rect 2914 1402 2942 1444
rect 2972 1430 2997 1444
rect 3096 1434 3121 1444
rect 2972 1402 3028 1430
rect 3058 1402 3092 1430
tri 3106 1427 3113 1434 ne
rect 3113 1402 3121 1434
rect 3151 1402 3199 1444
rect 3229 1434 3254 1444
rect 3229 1402 3237 1434
rect 3353 1430 3378 1444
rect 3258 1402 3292 1430
rect 3322 1402 3378 1430
rect 3408 1402 3436 1444
rect 3494 1402 3522 1444
rect 3552 1430 3577 1444
rect 3676 1434 3701 1444
rect 3552 1402 3608 1430
rect 3638 1402 3672 1430
tri 3686 1427 3693 1434 ne
rect 3693 1402 3701 1434
rect 3731 1402 3779 1444
rect 3809 1434 3834 1444
rect 3809 1402 3817 1434
rect 3933 1430 3958 1444
rect 3838 1402 3872 1430
rect 3902 1402 3958 1430
rect 3988 1402 4016 1444
rect 4074 1402 4102 1444
rect 4132 1430 4157 1444
rect 4256 1434 4281 1444
rect 4132 1402 4188 1430
rect 4218 1402 4252 1430
tri 4266 1427 4273 1434 ne
rect 4273 1402 4281 1434
rect 4311 1402 4359 1444
rect 4389 1434 4414 1444
rect 4389 1402 4397 1434
rect 4513 1430 4538 1444
rect 4418 1402 4452 1430
rect 4482 1402 4538 1430
rect 4568 1402 4596 1444
rect 4654 1402 4682 1444
rect 4712 1430 4737 1444
rect 4836 1434 4861 1444
rect 4712 1402 4768 1430
rect 4798 1402 4832 1430
tri 4846 1427 4853 1434 ne
rect 4853 1402 4861 1434
rect 4891 1402 4939 1444
rect 4969 1434 4994 1444
rect 4969 1402 4977 1434
rect 5093 1430 5118 1444
rect 4998 1402 5032 1430
rect 5062 1402 5118 1430
rect 5148 1402 5176 1444
rect 5234 1402 5262 1444
rect 5292 1430 5317 1444
rect 5416 1434 5441 1444
rect 5292 1402 5348 1430
rect 5378 1402 5412 1430
tri 5426 1427 5433 1434 ne
rect 5433 1402 5441 1434
rect 5471 1402 5519 1444
rect 5549 1434 5574 1444
rect 5549 1402 5557 1434
rect 5673 1430 5698 1444
rect 5578 1402 5612 1430
rect 5642 1402 5698 1430
rect 5728 1402 5756 1444
rect 5814 1402 5842 1444
rect 5872 1430 5897 1444
rect 5996 1434 6021 1444
rect 5872 1402 5928 1430
rect 5958 1402 5992 1430
tri 6006 1427 6013 1434 ne
rect 6013 1402 6021 1434
rect 6051 1402 6099 1444
rect 6129 1434 6154 1444
rect 6129 1402 6137 1434
rect 6253 1430 6278 1444
rect 6158 1402 6192 1430
rect 6222 1402 6278 1430
rect 6308 1402 6336 1444
rect 6394 1402 6422 1444
rect 6452 1430 6477 1444
rect 6576 1434 6601 1444
rect 6452 1402 6508 1430
rect 6538 1402 6572 1430
tri 6586 1427 6593 1434 ne
rect 6593 1402 6601 1434
rect 6631 1402 6679 1444
rect 6709 1434 6734 1444
rect 6709 1402 6717 1434
rect 6833 1430 6858 1444
rect 6738 1402 6772 1430
rect 6802 1402 6858 1430
rect 6888 1402 6916 1444
rect 165 1378 192 1402
rect 259 1380 291 1402
rect 259 1378 261 1380
rect 289 1378 291 1380
rect 358 1378 385 1402
rect 165 1364 259 1378
rect 291 1364 385 1378
rect 745 1378 772 1402
rect 839 1380 871 1402
rect 839 1378 841 1380
rect 869 1378 871 1380
rect 938 1378 965 1402
rect 745 1364 839 1378
rect 871 1364 965 1378
rect 1325 1378 1352 1402
rect 1419 1380 1451 1402
rect 1419 1378 1421 1380
rect 1449 1378 1451 1380
rect 1518 1378 1545 1402
rect 1325 1364 1419 1378
rect 1451 1364 1545 1378
rect 1905 1378 1932 1402
rect 1999 1380 2031 1402
rect 1999 1378 2001 1380
rect 2029 1378 2031 1380
rect 2098 1378 2125 1402
rect 1905 1364 1999 1378
rect 2031 1364 2125 1378
rect 2485 1378 2512 1402
rect 2579 1380 2611 1402
rect 2579 1378 2581 1380
rect 2609 1378 2611 1380
rect 2678 1378 2705 1402
rect 2485 1364 2579 1378
rect 2611 1364 2705 1378
rect 3065 1378 3092 1402
rect 3159 1380 3191 1402
rect 3159 1378 3161 1380
rect 3189 1378 3191 1380
rect 3258 1378 3285 1402
rect 3065 1364 3159 1378
rect 3191 1364 3285 1378
rect 3645 1378 3672 1402
rect 3739 1380 3771 1402
rect 3739 1378 3741 1380
rect 3769 1378 3771 1380
rect 3838 1378 3865 1402
rect 3645 1364 3739 1378
rect 3771 1364 3865 1378
rect 4225 1378 4252 1402
rect 4319 1380 4351 1402
rect 4319 1378 4321 1380
rect 4349 1378 4351 1380
rect 4418 1378 4445 1402
rect 4225 1364 4319 1378
rect 4351 1364 4445 1378
rect 4805 1378 4832 1402
rect 4899 1380 4931 1402
rect 4899 1378 4901 1380
rect 4929 1378 4931 1380
rect 4998 1378 5025 1402
rect 4805 1364 4899 1378
rect 4931 1364 5025 1378
rect 5385 1378 5412 1402
rect 5479 1380 5511 1402
rect 5479 1378 5481 1380
rect 5509 1378 5511 1380
rect 5578 1378 5605 1402
rect 5385 1364 5479 1378
rect 5511 1364 5605 1378
rect 5965 1378 5992 1402
rect 6059 1380 6091 1402
rect 6059 1378 6061 1380
rect 6089 1378 6091 1380
rect 6158 1378 6185 1402
rect 5965 1364 6059 1378
rect 6091 1364 6185 1378
rect 6545 1378 6572 1402
rect 6639 1380 6671 1402
rect 6639 1378 6641 1380
rect 6669 1378 6671 1380
rect 6738 1378 6765 1402
rect 6545 1364 6639 1378
rect 6671 1364 6765 1378
rect 88 1278 106 1306
rect 136 1278 154 1306
rect 396 1278 414 1306
rect 444 1278 463 1306
rect 668 1278 686 1306
rect 716 1278 734 1306
rect 976 1278 994 1306
rect 1024 1278 1043 1306
rect 1248 1278 1266 1306
rect 1296 1278 1314 1306
rect 1556 1278 1574 1306
rect 1604 1278 1623 1306
rect 1828 1278 1846 1306
rect 1876 1278 1894 1306
rect 2136 1278 2154 1306
rect 2184 1278 2203 1306
rect 2408 1278 2426 1306
rect 2456 1278 2474 1306
rect 2716 1278 2734 1306
rect 2764 1278 2783 1306
rect 2988 1278 3006 1306
rect 3036 1278 3054 1306
rect 3296 1278 3314 1306
rect 3344 1278 3363 1306
rect 3568 1278 3586 1306
rect 3616 1278 3634 1306
rect 3876 1278 3894 1306
rect 3924 1278 3943 1306
rect 4148 1278 4166 1306
rect 4196 1278 4214 1306
rect 4456 1278 4474 1306
rect 4504 1278 4523 1306
rect 4728 1278 4746 1306
rect 4776 1278 4794 1306
rect 5036 1278 5054 1306
rect 5084 1278 5103 1306
rect 5308 1278 5326 1306
rect 5356 1278 5374 1306
rect 5616 1278 5634 1306
rect 5664 1278 5683 1306
rect 5888 1278 5906 1306
rect 5936 1278 5954 1306
rect 6196 1278 6214 1306
rect 6244 1278 6263 1306
rect 6468 1278 6486 1306
rect 6516 1278 6534 1306
rect 6776 1278 6794 1306
rect 6824 1278 6843 1306
rect 14 1132 42 1174
rect 72 1160 97 1174
rect 196 1164 221 1174
rect 72 1132 128 1160
rect 158 1132 192 1160
tri 206 1157 213 1164 ne
rect 213 1132 221 1164
rect 251 1132 299 1174
rect 329 1164 354 1174
rect 329 1132 337 1164
rect 453 1160 478 1174
rect 358 1132 392 1160
rect 422 1132 478 1160
rect 508 1132 536 1174
rect 594 1132 622 1174
rect 652 1160 677 1174
rect 776 1164 801 1174
rect 652 1132 708 1160
rect 738 1132 772 1160
tri 786 1157 793 1164 ne
rect 793 1132 801 1164
rect 831 1132 879 1174
rect 909 1164 934 1174
rect 909 1132 917 1164
rect 1033 1160 1058 1174
rect 938 1132 972 1160
rect 1002 1132 1058 1160
rect 1088 1132 1116 1174
rect 1174 1132 1202 1174
rect 1232 1160 1257 1174
rect 1356 1164 1381 1174
rect 1232 1132 1288 1160
rect 1318 1132 1352 1160
tri 1366 1157 1373 1164 ne
rect 1373 1132 1381 1164
rect 1411 1132 1459 1174
rect 1489 1164 1514 1174
rect 1489 1132 1497 1164
rect 1613 1160 1638 1174
rect 1518 1132 1552 1160
rect 1582 1132 1638 1160
rect 1668 1132 1696 1174
rect 1754 1132 1782 1174
rect 1812 1160 1837 1174
rect 1936 1164 1961 1174
rect 1812 1132 1868 1160
rect 1898 1132 1932 1160
tri 1946 1157 1953 1164 ne
rect 1953 1132 1961 1164
rect 1991 1132 2039 1174
rect 2069 1164 2094 1174
rect 2069 1132 2077 1164
rect 2193 1160 2218 1174
rect 2098 1132 2132 1160
rect 2162 1132 2218 1160
rect 2248 1132 2276 1174
rect 2334 1132 2362 1174
rect 2392 1160 2417 1174
rect 2516 1164 2541 1174
rect 2392 1132 2448 1160
rect 2478 1132 2512 1160
tri 2526 1157 2533 1164 ne
rect 2533 1132 2541 1164
rect 2571 1132 2619 1174
rect 2649 1164 2674 1174
rect 2649 1132 2657 1164
rect 2773 1160 2798 1174
rect 2678 1132 2712 1160
rect 2742 1132 2798 1160
rect 2828 1132 2856 1174
rect 2914 1132 2942 1174
rect 2972 1160 2997 1174
rect 3096 1164 3121 1174
rect 2972 1132 3028 1160
rect 3058 1132 3092 1160
tri 3106 1157 3113 1164 ne
rect 3113 1132 3121 1164
rect 3151 1132 3199 1174
rect 3229 1164 3254 1174
rect 3229 1132 3237 1164
rect 3353 1160 3378 1174
rect 3258 1132 3292 1160
rect 3322 1132 3378 1160
rect 3408 1132 3436 1174
rect 3494 1132 3522 1174
rect 3552 1160 3577 1174
rect 3676 1164 3701 1174
rect 3552 1132 3608 1160
rect 3638 1132 3672 1160
tri 3686 1157 3693 1164 ne
rect 3693 1132 3701 1164
rect 3731 1132 3779 1174
rect 3809 1164 3834 1174
rect 3809 1132 3817 1164
rect 3933 1160 3958 1174
rect 3838 1132 3872 1160
rect 3902 1132 3958 1160
rect 3988 1132 4016 1174
rect 4074 1132 4102 1174
rect 4132 1160 4157 1174
rect 4256 1164 4281 1174
rect 4132 1132 4188 1160
rect 4218 1132 4252 1160
tri 4266 1157 4273 1164 ne
rect 4273 1132 4281 1164
rect 4311 1132 4359 1174
rect 4389 1164 4414 1174
rect 4389 1132 4397 1164
rect 4513 1160 4538 1174
rect 4418 1132 4452 1160
rect 4482 1132 4538 1160
rect 4568 1132 4596 1174
rect 4654 1132 4682 1174
rect 4712 1160 4737 1174
rect 4836 1164 4861 1174
rect 4712 1132 4768 1160
rect 4798 1132 4832 1160
tri 4846 1157 4853 1164 ne
rect 4853 1132 4861 1164
rect 4891 1132 4939 1174
rect 4969 1164 4994 1174
rect 4969 1132 4977 1164
rect 5093 1160 5118 1174
rect 4998 1132 5032 1160
rect 5062 1132 5118 1160
rect 5148 1132 5176 1174
rect 5234 1132 5262 1174
rect 5292 1160 5317 1174
rect 5416 1164 5441 1174
rect 5292 1132 5348 1160
rect 5378 1132 5412 1160
tri 5426 1157 5433 1164 ne
rect 5433 1132 5441 1164
rect 5471 1132 5519 1174
rect 5549 1164 5574 1174
rect 5549 1132 5557 1164
rect 5673 1160 5698 1174
rect 5578 1132 5612 1160
rect 5642 1132 5698 1160
rect 5728 1132 5756 1174
rect 5814 1132 5842 1174
rect 5872 1160 5897 1174
rect 5996 1164 6021 1174
rect 5872 1132 5928 1160
rect 5958 1132 5992 1160
tri 6006 1157 6013 1164 ne
rect 6013 1132 6021 1164
rect 6051 1132 6099 1174
rect 6129 1164 6154 1174
rect 6129 1132 6137 1164
rect 6253 1160 6278 1174
rect 6158 1132 6192 1160
rect 6222 1132 6278 1160
rect 6308 1132 6336 1174
rect 6394 1132 6422 1174
rect 6452 1160 6477 1174
rect 6576 1164 6601 1174
rect 6452 1132 6508 1160
rect 6538 1132 6572 1160
tri 6586 1157 6593 1164 ne
rect 6593 1132 6601 1164
rect 6631 1132 6679 1174
rect 6709 1164 6734 1174
rect 6709 1132 6717 1164
rect 6833 1160 6858 1174
rect 6738 1132 6772 1160
rect 6802 1132 6858 1160
rect 6888 1132 6916 1174
rect 165 1108 192 1132
rect 259 1110 291 1132
rect 259 1108 261 1110
rect 289 1108 291 1110
rect 358 1108 385 1132
rect 165 1094 259 1108
rect 291 1094 385 1108
rect 745 1108 772 1132
rect 839 1110 871 1132
rect 839 1108 841 1110
rect 869 1108 871 1110
rect 938 1108 965 1132
rect 745 1094 839 1108
rect 871 1094 965 1108
rect 1325 1108 1352 1132
rect 1419 1110 1451 1132
rect 1419 1108 1421 1110
rect 1449 1108 1451 1110
rect 1518 1108 1545 1132
rect 1325 1094 1419 1108
rect 1451 1094 1545 1108
rect 1905 1108 1932 1132
rect 1999 1110 2031 1132
rect 1999 1108 2001 1110
rect 2029 1108 2031 1110
rect 2098 1108 2125 1132
rect 1905 1094 1999 1108
rect 2031 1094 2125 1108
rect 2485 1108 2512 1132
rect 2579 1110 2611 1132
rect 2579 1108 2581 1110
rect 2609 1108 2611 1110
rect 2678 1108 2705 1132
rect 2485 1094 2579 1108
rect 2611 1094 2705 1108
rect 3065 1108 3092 1132
rect 3159 1110 3191 1132
rect 3159 1108 3161 1110
rect 3189 1108 3191 1110
rect 3258 1108 3285 1132
rect 3065 1094 3159 1108
rect 3191 1094 3285 1108
rect 3645 1108 3672 1132
rect 3739 1110 3771 1132
rect 3739 1108 3741 1110
rect 3769 1108 3771 1110
rect 3838 1108 3865 1132
rect 3645 1094 3739 1108
rect 3771 1094 3865 1108
rect 4225 1108 4252 1132
rect 4319 1110 4351 1132
rect 4319 1108 4321 1110
rect 4349 1108 4351 1110
rect 4418 1108 4445 1132
rect 4225 1094 4319 1108
rect 4351 1094 4445 1108
rect 4805 1108 4832 1132
rect 4899 1110 4931 1132
rect 4899 1108 4901 1110
rect 4929 1108 4931 1110
rect 4998 1108 5025 1132
rect 4805 1094 4899 1108
rect 4931 1094 5025 1108
rect 5385 1108 5412 1132
rect 5479 1110 5511 1132
rect 5479 1108 5481 1110
rect 5509 1108 5511 1110
rect 5578 1108 5605 1132
rect 5385 1094 5479 1108
rect 5511 1094 5605 1108
rect 5965 1108 5992 1132
rect 6059 1110 6091 1132
rect 6059 1108 6061 1110
rect 6089 1108 6091 1110
rect 6158 1108 6185 1132
rect 5965 1094 6059 1108
rect 6091 1094 6185 1108
rect 6545 1108 6572 1132
rect 6639 1110 6671 1132
rect 6639 1108 6641 1110
rect 6669 1108 6671 1110
rect 6738 1108 6765 1132
rect 6545 1094 6639 1108
rect 6671 1094 6765 1108
rect 88 1008 106 1036
rect 136 1008 154 1036
rect 396 1008 414 1036
rect 444 1008 463 1036
rect 668 1008 686 1036
rect 716 1008 734 1036
rect 976 1008 994 1036
rect 1024 1008 1043 1036
rect 1248 1008 1266 1036
rect 1296 1008 1314 1036
rect 1556 1008 1574 1036
rect 1604 1008 1623 1036
rect 1828 1008 1846 1036
rect 1876 1008 1894 1036
rect 2136 1008 2154 1036
rect 2184 1008 2203 1036
rect 2408 1008 2426 1036
rect 2456 1008 2474 1036
rect 2716 1008 2734 1036
rect 2764 1008 2783 1036
rect 2988 1008 3006 1036
rect 3036 1008 3054 1036
rect 3296 1008 3314 1036
rect 3344 1008 3363 1036
rect 3568 1008 3586 1036
rect 3616 1008 3634 1036
rect 3876 1008 3894 1036
rect 3924 1008 3943 1036
rect 4148 1008 4166 1036
rect 4196 1008 4214 1036
rect 4456 1008 4474 1036
rect 4504 1008 4523 1036
rect 4728 1007 4746 1035
rect 4776 1007 4794 1035
rect 5036 1007 5054 1035
rect 5084 1007 5103 1035
rect 5308 1007 5326 1035
rect 5356 1007 5374 1035
rect 14 862 42 904
rect 72 890 97 904
rect 196 894 221 904
rect 72 862 128 890
rect 158 862 192 890
tri 206 887 213 894 ne
rect 213 862 221 894
rect 251 862 299 904
rect 329 894 354 904
rect 329 862 337 894
rect 453 890 478 904
rect 358 862 392 890
rect 422 862 478 890
rect 508 862 536 904
rect 594 862 622 904
rect 652 890 677 904
rect 776 894 801 904
rect 652 862 708 890
rect 738 862 772 890
tri 786 887 793 894 ne
rect 793 862 801 894
rect 831 862 879 904
rect 909 894 934 904
rect 909 862 917 894
rect 1033 890 1058 904
rect 938 862 972 890
rect 1002 862 1058 890
rect 1088 862 1116 904
rect 1174 862 1202 904
rect 1232 890 1257 904
rect 1356 894 1381 904
rect 1232 862 1288 890
rect 1318 862 1352 890
tri 1366 887 1373 894 ne
rect 1373 862 1381 894
rect 1411 862 1459 904
rect 1489 894 1514 904
rect 1489 862 1497 894
rect 1613 890 1638 904
rect 1518 862 1552 890
rect 1582 862 1638 890
rect 1668 862 1696 904
rect 1754 862 1782 904
rect 1812 890 1837 904
rect 1936 894 1961 904
rect 1812 862 1868 890
rect 1898 862 1932 890
tri 1946 887 1953 894 ne
rect 1953 862 1961 894
rect 1991 862 2039 904
rect 2069 894 2094 904
rect 2069 862 2077 894
rect 2193 890 2218 904
rect 2098 862 2132 890
rect 2162 862 2218 890
rect 2248 862 2276 904
rect 2334 862 2362 904
rect 2392 890 2417 904
rect 2516 894 2541 904
rect 2392 862 2448 890
rect 2478 862 2512 890
tri 2526 887 2533 894 ne
rect 2533 862 2541 894
rect 2571 862 2619 904
rect 2649 894 2674 904
rect 2649 862 2657 894
rect 2773 890 2798 904
rect 2678 862 2712 890
rect 2742 862 2798 890
rect 2828 862 2856 904
rect 2914 862 2942 904
rect 2972 890 2997 904
rect 3096 894 3121 904
rect 2972 862 3028 890
rect 3058 862 3092 890
tri 3106 887 3113 894 ne
rect 3113 862 3121 894
rect 3151 862 3199 904
rect 3229 894 3254 904
rect 3229 862 3237 894
rect 3353 890 3378 904
rect 3258 862 3292 890
rect 3322 862 3378 890
rect 3408 862 3436 904
rect 3494 862 3522 904
rect 3552 890 3577 904
rect 3676 894 3701 904
rect 3552 862 3608 890
rect 3638 862 3672 890
tri 3686 887 3693 894 ne
rect 3693 862 3701 894
rect 3731 862 3779 904
rect 3809 894 3834 904
rect 3809 862 3817 894
rect 3933 890 3958 904
rect 3838 862 3872 890
rect 3902 862 3958 890
rect 3988 862 4016 904
rect 4074 862 4102 904
rect 4132 890 4157 904
rect 4256 894 4281 904
rect 4132 862 4188 890
rect 4218 862 4252 890
tri 4266 887 4273 894 ne
rect 4273 862 4281 894
rect 4311 862 4359 904
rect 4389 894 4414 904
rect 4389 862 4397 894
rect 4513 890 4538 904
rect 4418 862 4452 890
rect 4482 862 4538 890
rect 4568 862 4596 904
rect 5616 1007 5634 1035
rect 5664 1007 5683 1035
rect 5888 1007 5906 1035
rect 5936 1007 5954 1035
rect 6196 1007 6214 1035
rect 6244 1007 6263 1035
rect 6468 1007 6486 1035
rect 6516 1007 6534 1035
rect 6776 1007 6794 1035
rect 6824 1007 6843 1035
rect 165 838 192 862
rect 259 840 291 862
rect 259 838 261 840
rect 289 838 291 840
rect 358 838 385 862
rect 165 824 259 838
rect 291 824 385 838
rect 745 838 772 862
rect 839 840 871 862
rect 839 838 841 840
rect 869 838 871 840
rect 938 838 965 862
rect 745 824 839 838
rect 871 824 965 838
rect 1325 838 1352 862
rect 1419 840 1451 862
rect 1419 838 1421 840
rect 1449 838 1451 840
rect 1518 838 1545 862
rect 1325 824 1419 838
rect 1451 824 1545 838
rect 1905 838 1932 862
rect 1999 840 2031 862
rect 1999 838 2001 840
rect 2029 838 2031 840
rect 2098 838 2125 862
rect 1905 824 1999 838
rect 2031 824 2125 838
rect 2485 838 2512 862
rect 2579 840 2611 862
rect 2579 838 2581 840
rect 2609 838 2611 840
rect 2678 838 2705 862
rect 2485 824 2579 838
rect 2611 824 2705 838
rect 3065 838 3092 862
rect 3159 840 3191 862
rect 3159 838 3161 840
rect 3189 838 3191 840
rect 3258 838 3285 862
rect 3065 824 3159 838
rect 3191 824 3285 838
rect 3645 838 3672 862
rect 3739 840 3771 862
rect 3739 838 3741 840
rect 3769 838 3771 840
rect 3838 838 3865 862
rect 3645 824 3739 838
rect 3771 824 3865 838
rect 4225 838 4252 862
rect 4319 840 4351 862
rect 4319 838 4321 840
rect 4349 838 4351 840
rect 4418 838 4445 862
rect 4654 861 4682 903
rect 4712 889 4737 903
rect 4836 893 4861 903
rect 4712 861 4768 889
rect 4798 861 4832 889
tri 4846 886 4853 893 ne
rect 4853 861 4861 893
rect 4891 861 4939 903
rect 4969 893 4994 903
rect 4969 861 4977 893
rect 5093 889 5118 903
rect 4998 861 5032 889
rect 5062 861 5118 889
rect 5148 861 5176 903
rect 5234 861 5262 903
rect 5292 889 5317 903
rect 5416 893 5441 903
rect 5292 861 5348 889
rect 5378 861 5412 889
tri 5426 886 5433 893 ne
rect 5433 861 5441 893
rect 5471 861 5519 903
rect 5549 893 5574 903
rect 5549 861 5557 893
rect 5673 889 5698 903
rect 5578 861 5612 889
rect 5642 861 5698 889
rect 5728 861 5756 903
rect 5814 861 5842 903
rect 5872 889 5897 903
rect 5996 893 6021 903
rect 5872 861 5928 889
rect 5958 861 5992 889
tri 6006 886 6013 893 ne
rect 6013 861 6021 893
rect 6051 861 6099 903
rect 6129 893 6154 903
rect 6129 861 6137 893
rect 6253 889 6278 903
rect 6158 861 6192 889
rect 6222 861 6278 889
rect 6308 861 6336 903
rect 6394 861 6422 903
rect 6452 889 6477 903
rect 6576 893 6601 903
rect 6452 861 6508 889
rect 6538 861 6572 889
tri 6586 886 6593 893 ne
rect 6593 861 6601 893
rect 6631 861 6679 903
rect 6709 893 6734 903
rect 6709 861 6717 893
rect 6833 889 6858 903
rect 6738 861 6772 889
rect 6802 861 6858 889
rect 6888 861 6916 903
rect 4225 824 4319 838
rect 4351 824 4445 838
rect 4805 837 4832 861
rect 4899 839 4931 861
rect 4899 837 4901 839
rect 4929 837 4931 839
rect 4998 837 5025 861
rect 4805 823 4899 837
rect 4931 823 5025 837
rect 5385 837 5412 861
rect 5479 839 5511 861
rect 5479 837 5481 839
rect 5509 837 5511 839
rect 5578 837 5605 861
rect 5385 823 5479 837
rect 5511 823 5605 837
rect 5965 837 5992 861
rect 6059 839 6091 861
rect 6059 837 6061 839
rect 6089 837 6091 839
rect 6158 837 6185 861
rect 5965 823 6059 837
rect 6091 823 6185 837
rect 6545 837 6572 861
rect 6639 839 6671 861
rect 6639 837 6641 839
rect 6669 837 6671 839
rect 6738 837 6765 861
rect 6545 823 6639 837
rect 6671 823 6765 837
rect 88 738 106 766
rect 136 738 154 766
rect 396 738 414 766
rect 444 738 463 766
rect 668 738 686 766
rect 716 738 734 766
rect 976 738 994 766
rect 1024 738 1043 766
rect 1248 738 1266 766
rect 1296 738 1314 766
rect 1556 738 1574 766
rect 1604 738 1623 766
rect 1828 738 1846 766
rect 1876 738 1894 766
rect 2136 738 2154 766
rect 2184 738 2203 766
rect 2408 738 2426 766
rect 2456 738 2474 766
rect 2716 738 2734 766
rect 2764 738 2783 766
rect 2988 738 3006 766
rect 3036 738 3054 766
rect 3296 738 3314 766
rect 3344 738 3363 766
rect 3568 738 3586 766
rect 3616 738 3634 766
rect 3876 738 3894 766
rect 3924 738 3943 766
rect 4148 738 4166 766
rect 4196 738 4214 766
rect 4456 738 4474 766
rect 4504 738 4523 766
rect 4728 737 4746 765
rect 4776 737 4794 765
rect 5036 737 5054 765
rect 5084 737 5103 765
rect 5308 737 5326 765
rect 5356 737 5374 765
rect 14 592 42 634
rect 72 620 97 634
rect 196 624 221 634
rect 72 592 128 620
rect 158 592 192 620
tri 206 617 213 624 ne
rect 213 592 221 624
rect 251 592 299 634
rect 329 624 354 634
rect 329 592 337 624
rect 453 620 478 634
rect 358 592 392 620
rect 422 592 478 620
rect 508 592 536 634
rect 594 592 622 634
rect 652 620 677 634
rect 776 624 801 634
rect 652 592 708 620
rect 738 592 772 620
tri 786 617 793 624 ne
rect 793 592 801 624
rect 831 592 879 634
rect 909 624 934 634
rect 909 592 917 624
rect 1033 620 1058 634
rect 938 592 972 620
rect 1002 592 1058 620
rect 1088 592 1116 634
rect 1174 592 1202 634
rect 1232 620 1257 634
rect 1356 624 1381 634
rect 1232 592 1288 620
rect 1318 592 1352 620
tri 1366 617 1373 624 ne
rect 1373 592 1381 624
rect 1411 592 1459 634
rect 1489 624 1514 634
rect 1489 592 1497 624
rect 1613 620 1638 634
rect 1518 592 1552 620
rect 1582 592 1638 620
rect 1668 592 1696 634
rect 1754 592 1782 634
rect 1812 620 1837 634
rect 1936 624 1961 634
rect 1812 592 1868 620
rect 1898 592 1932 620
tri 1946 617 1953 624 ne
rect 1953 592 1961 624
rect 1991 592 2039 634
rect 2069 624 2094 634
rect 2069 592 2077 624
rect 2193 620 2218 634
rect 2098 592 2132 620
rect 2162 592 2218 620
rect 2248 592 2276 634
rect 2334 592 2362 634
rect 2392 620 2417 634
rect 2516 624 2541 634
rect 2392 592 2448 620
rect 2478 592 2512 620
tri 2526 617 2533 624 ne
rect 2533 592 2541 624
rect 2571 592 2619 634
rect 2649 624 2674 634
rect 2649 592 2657 624
rect 2773 620 2798 634
rect 2678 592 2712 620
rect 2742 592 2798 620
rect 2828 592 2856 634
rect 2914 592 2942 634
rect 2972 620 2997 634
rect 3096 624 3121 634
rect 2972 592 3028 620
rect 3058 592 3092 620
tri 3106 617 3113 624 ne
rect 3113 592 3121 624
rect 3151 592 3199 634
rect 3229 624 3254 634
rect 3229 592 3237 624
rect 3353 620 3378 634
rect 3258 592 3292 620
rect 3322 592 3378 620
rect 3408 592 3436 634
rect 3494 592 3522 634
rect 3552 620 3577 634
rect 3676 624 3701 634
rect 3552 592 3608 620
rect 3638 592 3672 620
tri 3686 617 3693 624 ne
rect 3693 592 3701 624
rect 3731 592 3779 634
rect 3809 624 3834 634
rect 3809 592 3817 624
rect 3933 620 3958 634
rect 3838 592 3872 620
rect 3902 592 3958 620
rect 3988 592 4016 634
rect 4074 592 4102 634
rect 4132 620 4157 634
rect 4256 624 4281 634
rect 4132 592 4188 620
rect 4218 592 4252 620
tri 4266 617 4273 624 ne
rect 4273 592 4281 624
rect 4311 592 4359 634
rect 4389 624 4414 634
rect 4389 592 4397 624
rect 4513 620 4538 634
rect 4418 592 4452 620
rect 4482 592 4538 620
rect 4568 592 4596 634
rect 5616 737 5634 765
rect 5664 737 5683 765
rect 5888 737 5906 765
rect 5936 737 5954 765
rect 6196 737 6214 765
rect 6244 737 6263 765
rect 6468 737 6486 765
rect 6516 737 6534 765
rect 6776 737 6794 765
rect 6824 737 6843 765
rect 165 568 192 592
rect 259 570 291 592
rect 259 568 261 570
rect 289 568 291 570
rect 358 568 385 592
rect 165 554 259 568
rect 291 554 385 568
rect 745 568 772 592
rect 839 570 871 592
rect 839 568 841 570
rect 869 568 871 570
rect 938 568 965 592
rect 745 554 839 568
rect 871 554 965 568
rect 1325 568 1352 592
rect 1419 570 1451 592
rect 1419 568 1421 570
rect 1449 568 1451 570
rect 1518 568 1545 592
rect 1325 554 1419 568
rect 1451 554 1545 568
rect 1905 568 1932 592
rect 1999 570 2031 592
rect 1999 568 2001 570
rect 2029 568 2031 570
rect 2098 568 2125 592
rect 1905 554 1999 568
rect 2031 554 2125 568
rect 2485 568 2512 592
rect 2579 570 2611 592
rect 2579 568 2581 570
rect 2609 568 2611 570
rect 2678 568 2705 592
rect 2485 554 2579 568
rect 2611 554 2705 568
rect 3065 568 3092 592
rect 3159 570 3191 592
rect 3159 568 3161 570
rect 3189 568 3191 570
rect 3258 568 3285 592
rect 3065 554 3159 568
rect 3191 554 3285 568
rect 3645 568 3672 592
rect 3739 570 3771 592
rect 3739 568 3741 570
rect 3769 568 3771 570
rect 3838 568 3865 592
rect 3645 554 3739 568
rect 3771 554 3865 568
rect 4225 568 4252 592
rect 4319 570 4351 592
rect 4319 568 4321 570
rect 4349 568 4351 570
rect 4418 568 4445 592
rect 4654 591 4682 633
rect 4712 619 4737 633
rect 4836 623 4861 633
rect 4712 591 4768 619
rect 4798 591 4832 619
tri 4846 616 4853 623 ne
rect 4853 591 4861 623
rect 4891 591 4939 633
rect 4969 623 4994 633
rect 4969 591 4977 623
rect 5093 619 5118 633
rect 4998 591 5032 619
rect 5062 591 5118 619
rect 5148 591 5176 633
rect 5234 591 5262 633
rect 5292 619 5317 633
rect 5416 623 5441 633
rect 5292 591 5348 619
rect 5378 591 5412 619
tri 5426 616 5433 623 ne
rect 5433 591 5441 623
rect 5471 591 5519 633
rect 5549 623 5574 633
rect 5549 591 5557 623
rect 5673 619 5698 633
rect 5578 591 5612 619
rect 5642 591 5698 619
rect 5728 591 5756 633
rect 5814 591 5842 633
rect 5872 619 5897 633
rect 5996 623 6021 633
rect 5872 591 5928 619
rect 5958 591 5992 619
tri 6006 616 6013 623 ne
rect 6013 591 6021 623
rect 6051 591 6099 633
rect 6129 623 6154 633
rect 6129 591 6137 623
rect 6253 619 6278 633
rect 6158 591 6192 619
rect 6222 591 6278 619
rect 6308 591 6336 633
rect 6394 591 6422 633
rect 6452 619 6477 633
rect 6576 623 6601 633
rect 6452 591 6508 619
rect 6538 591 6572 619
tri 6586 616 6593 623 ne
rect 6593 591 6601 623
rect 6631 591 6679 633
rect 6709 623 6734 633
rect 6709 591 6717 623
rect 6833 619 6858 633
rect 6738 591 6772 619
rect 6802 591 6858 619
rect 6888 591 6916 633
rect 4225 554 4319 568
rect 4351 554 4445 568
rect 4805 567 4832 591
rect 4899 569 4931 591
rect 4899 567 4901 569
rect 4929 567 4931 569
rect 4998 567 5025 591
rect 4805 553 4899 567
rect 4931 553 5025 567
rect 5385 567 5412 591
rect 5479 569 5511 591
rect 5479 567 5481 569
rect 5509 567 5511 569
rect 5578 567 5605 591
rect 5385 553 5479 567
rect 5511 553 5605 567
rect 5965 567 5992 591
rect 6059 569 6091 591
rect 6059 567 6061 569
rect 6089 567 6091 569
rect 6158 567 6185 591
rect 5965 553 6059 567
rect 6091 553 6185 567
rect 6545 567 6572 591
rect 6639 569 6671 591
rect 6639 567 6641 569
rect 6669 567 6671 569
rect 6738 567 6765 591
rect 6545 553 6639 567
rect 6671 553 6765 567
rect 88 468 106 496
rect 136 468 154 496
rect 396 468 414 496
rect 444 468 463 496
rect 668 468 686 496
rect 716 468 734 496
rect 976 468 994 496
rect 1024 468 1043 496
rect 1248 468 1266 496
rect 1296 468 1314 496
rect 1556 468 1574 496
rect 1604 468 1623 496
rect 1828 468 1846 496
rect 1876 468 1894 496
rect 2136 468 2154 496
rect 2184 468 2203 496
rect 2408 468 2426 496
rect 2456 468 2474 496
rect 2716 468 2734 496
rect 2764 468 2783 496
rect 2988 468 3006 496
rect 3036 468 3054 496
rect 3296 468 3314 496
rect 3344 468 3363 496
rect 3568 468 3586 496
rect 3616 468 3634 496
rect 3876 468 3894 496
rect 3924 468 3943 496
rect 4148 468 4166 496
rect 4196 468 4214 496
rect 4456 468 4474 496
rect 4504 468 4523 496
rect 4728 467 4746 495
rect 4776 467 4794 495
rect 5036 467 5054 495
rect 5084 467 5103 495
rect 5308 467 5326 495
rect 5356 467 5374 495
rect 14 322 42 364
rect 72 350 97 364
rect 196 354 221 364
rect 72 322 128 350
rect 158 322 192 350
tri 206 347 213 354 ne
rect 213 322 221 354
rect 251 322 299 364
rect 329 354 354 364
rect 329 322 337 354
rect 453 350 478 364
rect 358 322 392 350
rect 422 322 478 350
rect 508 322 536 364
rect 594 322 622 364
rect 652 350 677 364
rect 776 354 801 364
rect 652 322 708 350
rect 738 322 772 350
tri 786 347 793 354 ne
rect 793 322 801 354
rect 831 322 879 364
rect 909 354 934 364
rect 909 322 917 354
rect 1033 350 1058 364
rect 938 322 972 350
rect 1002 322 1058 350
rect 1088 322 1116 364
rect 1174 322 1202 364
rect 1232 350 1257 364
rect 1356 354 1381 364
rect 1232 322 1288 350
rect 1318 322 1352 350
tri 1366 347 1373 354 ne
rect 1373 322 1381 354
rect 1411 322 1459 364
rect 1489 354 1514 364
rect 1489 322 1497 354
rect 1613 350 1638 364
rect 1518 322 1552 350
rect 1582 322 1638 350
rect 1668 322 1696 364
rect 1754 322 1782 364
rect 1812 350 1837 364
rect 1936 354 1961 364
rect 1812 322 1868 350
rect 1898 322 1932 350
tri 1946 347 1953 354 ne
rect 1953 322 1961 354
rect 1991 322 2039 364
rect 2069 354 2094 364
rect 2069 322 2077 354
rect 2193 350 2218 364
rect 2098 322 2132 350
rect 2162 322 2218 350
rect 2248 322 2276 364
rect 2334 322 2362 364
rect 2392 350 2417 364
rect 2516 354 2541 364
rect 2392 322 2448 350
rect 2478 322 2512 350
tri 2526 347 2533 354 ne
rect 2533 322 2541 354
rect 2571 322 2619 364
rect 2649 354 2674 364
rect 2649 322 2657 354
rect 2773 350 2798 364
rect 2678 322 2712 350
rect 2742 322 2798 350
rect 2828 322 2856 364
rect 2914 322 2942 364
rect 2972 350 2997 364
rect 3096 354 3121 364
rect 2972 322 3028 350
rect 3058 322 3092 350
tri 3106 347 3113 354 ne
rect 3113 322 3121 354
rect 3151 322 3199 364
rect 3229 354 3254 364
rect 3229 322 3237 354
rect 3353 350 3378 364
rect 3258 322 3292 350
rect 3322 322 3378 350
rect 3408 322 3436 364
rect 3494 322 3522 364
rect 3552 350 3577 364
rect 3676 354 3701 364
rect 3552 322 3608 350
rect 3638 322 3672 350
tri 3686 347 3693 354 ne
rect 3693 322 3701 354
rect 3731 322 3779 364
rect 3809 354 3834 364
rect 3809 322 3817 354
rect 3933 350 3958 364
rect 3838 322 3872 350
rect 3902 322 3958 350
rect 3988 322 4016 364
rect 4074 322 4102 364
rect 4132 350 4157 364
rect 4256 354 4281 364
rect 4132 322 4188 350
rect 4218 322 4252 350
tri 4266 347 4273 354 ne
rect 4273 322 4281 354
rect 4311 322 4359 364
rect 4389 354 4414 364
rect 4389 322 4397 354
rect 4513 350 4538 364
rect 4418 322 4452 350
rect 4482 322 4538 350
rect 4568 322 4596 364
rect 5616 467 5634 495
rect 5664 467 5683 495
rect 5888 467 5906 495
rect 5936 467 5954 495
rect 6196 467 6214 495
rect 6244 467 6263 495
rect 6468 467 6486 495
rect 6516 467 6534 495
rect 6776 467 6794 495
rect 6824 467 6843 495
rect 165 298 192 322
rect 259 300 291 322
rect 259 298 261 300
rect 289 298 291 300
rect 358 298 385 322
rect 165 284 259 298
rect 291 284 385 298
rect 745 298 772 322
rect 839 300 871 322
rect 839 298 841 300
rect 869 298 871 300
rect 938 298 965 322
rect 745 284 839 298
rect 871 284 965 298
rect 1325 298 1352 322
rect 1419 300 1451 322
rect 1419 298 1421 300
rect 1449 298 1451 300
rect 1518 298 1545 322
rect 1325 284 1419 298
rect 1451 284 1545 298
rect 1905 298 1932 322
rect 1999 300 2031 322
rect 1999 298 2001 300
rect 2029 298 2031 300
rect 2098 298 2125 322
rect 1905 284 1999 298
rect 2031 284 2125 298
rect 2485 298 2512 322
rect 2579 300 2611 322
rect 2579 298 2581 300
rect 2609 298 2611 300
rect 2678 298 2705 322
rect 2485 284 2579 298
rect 2611 284 2705 298
rect 3065 298 3092 322
rect 3159 300 3191 322
rect 3159 298 3161 300
rect 3189 298 3191 300
rect 3258 298 3285 322
rect 3065 284 3159 298
rect 3191 284 3285 298
rect 3645 298 3672 322
rect 3739 300 3771 322
rect 3739 298 3741 300
rect 3769 298 3771 300
rect 3838 298 3865 322
rect 3645 284 3739 298
rect 3771 284 3865 298
rect 4225 298 4252 322
rect 4319 300 4351 322
rect 4319 298 4321 300
rect 4349 298 4351 300
rect 4418 298 4445 322
rect 4654 321 4682 363
rect 4712 349 4737 363
rect 4836 353 4861 363
rect 4712 321 4768 349
rect 4798 321 4832 349
tri 4846 346 4853 353 ne
rect 4853 321 4861 353
rect 4891 321 4939 363
rect 4969 353 4994 363
rect 4969 321 4977 353
rect 5093 349 5118 363
rect 4998 321 5032 349
rect 5062 321 5118 349
rect 5148 321 5176 363
rect 5234 321 5262 363
rect 5292 349 5317 363
rect 5416 353 5441 363
rect 5292 321 5348 349
rect 5378 321 5412 349
tri 5426 346 5433 353 ne
rect 5433 321 5441 353
rect 5471 321 5519 363
rect 5549 353 5574 363
rect 5549 321 5557 353
rect 5673 349 5698 363
rect 5578 321 5612 349
rect 5642 321 5698 349
rect 5728 321 5756 363
rect 5814 321 5842 363
rect 5872 349 5897 363
rect 5996 353 6021 363
rect 5872 321 5928 349
rect 5958 321 5992 349
tri 6006 346 6013 353 ne
rect 6013 321 6021 353
rect 6051 321 6099 363
rect 6129 353 6154 363
rect 6129 321 6137 353
rect 6253 349 6278 363
rect 6158 321 6192 349
rect 6222 321 6278 349
rect 6308 321 6336 363
rect 6394 321 6422 363
rect 6452 349 6477 363
rect 6576 353 6601 363
rect 6452 321 6508 349
rect 6538 321 6572 349
tri 6586 346 6593 353 ne
rect 6593 321 6601 353
rect 6631 321 6679 363
rect 6709 353 6734 363
rect 6709 321 6717 353
rect 6833 349 6858 363
rect 6738 321 6772 349
rect 6802 321 6858 349
rect 6888 321 6916 363
rect 4225 284 4319 298
rect 4351 284 4445 298
rect 4805 297 4832 321
rect 4899 299 4931 321
rect 4899 297 4901 299
rect 4929 297 4931 299
rect 4998 297 5025 321
rect 4805 283 4899 297
rect 4931 283 5025 297
rect 5385 297 5412 321
rect 5479 299 5511 321
rect 5479 297 5481 299
rect 5509 297 5511 299
rect 5578 297 5605 321
rect 5385 283 5479 297
rect 5511 283 5605 297
rect 5965 297 5992 321
rect 6059 299 6091 321
rect 6059 297 6061 299
rect 6089 297 6091 299
rect 6158 297 6185 321
rect 5965 283 6059 297
rect 6091 283 6185 297
rect 6545 297 6572 321
rect 6639 299 6671 321
rect 6639 297 6641 299
rect 6669 297 6671 299
rect 6738 297 6765 321
rect 6545 283 6639 297
rect 6671 283 6765 297
rect 88 198 106 226
rect 136 198 154 226
rect 396 198 414 226
rect 444 198 463 226
rect 668 198 686 226
rect 716 198 734 226
rect 976 198 994 226
rect 1024 198 1043 226
rect 1248 198 1266 226
rect 1296 198 1314 226
rect 1556 198 1574 226
rect 1604 198 1623 226
rect 1828 198 1846 226
rect 1876 198 1894 226
rect 2136 198 2154 226
rect 2184 198 2203 226
rect 2408 198 2426 226
rect 2456 198 2474 226
rect 2716 198 2734 226
rect 2764 198 2783 226
rect 2988 198 3006 226
rect 3036 198 3054 226
rect 3296 198 3314 226
rect 3344 198 3363 226
rect 3568 198 3586 226
rect 3616 198 3634 226
rect 3876 198 3894 226
rect 3924 198 3943 226
rect 4148 198 4166 226
rect 4196 198 4214 226
rect 4456 198 4474 226
rect 4504 198 4523 226
rect 4728 197 4746 225
rect 4776 197 4794 225
rect 5036 197 5054 225
rect 5084 197 5103 225
rect 5308 197 5326 225
rect 5356 197 5374 225
rect 14 52 42 94
rect 72 80 97 94
rect 196 84 221 94
rect 72 52 128 80
rect 158 52 192 80
tri 206 77 213 84 ne
rect 213 52 221 84
rect 251 52 299 94
rect 329 84 354 94
rect 329 52 337 84
rect 453 80 478 94
rect 358 52 392 80
rect 422 52 478 80
rect 508 52 536 94
rect 594 52 622 94
rect 652 80 677 94
rect 776 84 801 94
rect 652 52 708 80
rect 738 52 772 80
tri 786 77 793 84 ne
rect 793 52 801 84
rect 831 52 879 94
rect 909 84 934 94
rect 909 52 917 84
rect 1033 80 1058 94
rect 938 52 972 80
rect 1002 52 1058 80
rect 1088 52 1116 94
rect 1174 52 1202 94
rect 1232 80 1257 94
rect 1356 84 1381 94
rect 1232 52 1288 80
rect 1318 52 1352 80
tri 1366 77 1373 84 ne
rect 1373 52 1381 84
rect 1411 52 1459 94
rect 1489 84 1514 94
rect 1489 52 1497 84
rect 1613 80 1638 94
rect 1518 52 1552 80
rect 1582 52 1638 80
rect 1668 52 1696 94
rect 1754 52 1782 94
rect 1812 80 1837 94
rect 1936 84 1961 94
rect 1812 52 1868 80
rect 1898 52 1932 80
tri 1946 77 1953 84 ne
rect 1953 52 1961 84
rect 1991 52 2039 94
rect 2069 84 2094 94
rect 2069 52 2077 84
rect 2193 80 2218 94
rect 2098 52 2132 80
rect 2162 52 2218 80
rect 2248 52 2276 94
rect 2334 52 2362 94
rect 2392 80 2417 94
rect 2516 84 2541 94
rect 2392 52 2448 80
rect 2478 52 2512 80
tri 2526 77 2533 84 ne
rect 2533 52 2541 84
rect 2571 52 2619 94
rect 2649 84 2674 94
rect 2649 52 2657 84
rect 2773 80 2798 94
rect 2678 52 2712 80
rect 2742 52 2798 80
rect 2828 52 2856 94
rect 2914 52 2942 94
rect 2972 80 2997 94
rect 3096 84 3121 94
rect 2972 52 3028 80
rect 3058 52 3092 80
tri 3106 77 3113 84 ne
rect 3113 52 3121 84
rect 3151 52 3199 94
rect 3229 84 3254 94
rect 3229 52 3237 84
rect 3353 80 3378 94
rect 3258 52 3292 80
rect 3322 52 3378 80
rect 3408 52 3436 94
rect 3494 52 3522 94
rect 3552 80 3577 94
rect 3676 84 3701 94
rect 3552 52 3608 80
rect 3638 52 3672 80
tri 3686 77 3693 84 ne
rect 3693 52 3701 84
rect 3731 52 3779 94
rect 3809 84 3834 94
rect 3809 52 3817 84
rect 3933 80 3958 94
rect 3838 52 3872 80
rect 3902 52 3958 80
rect 3988 52 4016 94
rect 4074 52 4102 94
rect 4132 80 4157 94
rect 4256 84 4281 94
rect 4132 52 4188 80
rect 4218 52 4252 80
tri 4266 77 4273 84 ne
rect 4273 52 4281 84
rect 4311 52 4359 94
rect 4389 84 4414 94
rect 4389 52 4397 84
rect 4513 80 4538 94
rect 4418 52 4452 80
rect 4482 52 4538 80
rect 4568 52 4596 94
rect 5616 197 5634 225
rect 5664 197 5683 225
rect 5888 197 5906 225
rect 5936 197 5954 225
rect 6196 197 6214 225
rect 6244 197 6263 225
rect 6468 197 6486 225
rect 6516 197 6534 225
rect 6776 197 6794 225
rect 6824 197 6843 225
rect 165 28 192 52
rect 259 30 291 52
rect 259 28 261 30
rect 289 28 291 30
rect 358 28 385 52
rect 165 14 259 28
rect 291 14 385 28
rect 745 28 772 52
rect 839 30 871 52
rect 839 28 841 30
rect 869 28 871 30
rect 938 28 965 52
rect 745 14 839 28
rect 871 14 965 28
rect 1325 28 1352 52
rect 1419 30 1451 52
rect 1419 28 1421 30
rect 1449 28 1451 30
rect 1518 28 1545 52
rect 1325 14 1419 28
rect 1451 14 1545 28
rect 1905 28 1932 52
rect 1999 30 2031 52
rect 1999 28 2001 30
rect 2029 28 2031 30
rect 2098 28 2125 52
rect 1905 14 1999 28
rect 2031 14 2125 28
rect 2485 28 2512 52
rect 2579 30 2611 52
rect 2579 28 2581 30
rect 2609 28 2611 30
rect 2678 28 2705 52
rect 2485 14 2579 28
rect 2611 14 2705 28
rect 3065 28 3092 52
rect 3159 30 3191 52
rect 3159 28 3161 30
rect 3189 28 3191 30
rect 3258 28 3285 52
rect 3065 14 3159 28
rect 3191 14 3285 28
rect 3645 28 3672 52
rect 3739 30 3771 52
rect 3739 28 3741 30
rect 3769 28 3771 30
rect 3838 28 3865 52
rect 3645 14 3739 28
rect 3771 14 3865 28
rect 4225 28 4252 52
rect 4319 30 4351 52
rect 4319 28 4321 30
rect 4349 28 4351 30
rect 4418 28 4445 52
rect 4654 51 4682 93
rect 4712 79 4737 93
rect 4836 83 4861 93
rect 4712 51 4768 79
rect 4798 51 4832 79
tri 4846 76 4853 83 ne
rect 4853 51 4861 83
rect 4891 51 4939 93
rect 4969 83 4994 93
rect 4969 51 4977 83
rect 5093 79 5118 93
rect 4998 51 5032 79
rect 5062 51 5118 79
rect 5148 51 5176 93
rect 5234 51 5262 93
rect 5292 79 5317 93
rect 5416 83 5441 93
rect 5292 51 5348 79
rect 5378 51 5412 79
tri 5426 76 5433 83 ne
rect 5433 51 5441 83
rect 5471 51 5519 93
rect 5549 83 5574 93
rect 5549 51 5557 83
rect 5673 79 5698 93
rect 5578 51 5612 79
rect 5642 51 5698 79
rect 5728 51 5756 93
rect 5814 51 5842 93
rect 5872 79 5897 93
rect 5996 83 6021 93
rect 5872 51 5928 79
rect 5958 51 5992 79
tri 6006 76 6013 83 ne
rect 6013 51 6021 83
rect 6051 51 6099 93
rect 6129 83 6154 93
rect 6129 51 6137 83
rect 6253 79 6278 93
rect 6158 51 6192 79
rect 6222 51 6278 79
rect 6308 51 6336 93
rect 6394 51 6422 93
rect 6452 79 6477 93
rect 6576 83 6601 93
rect 6452 51 6508 79
rect 6538 51 6572 79
tri 6586 76 6593 83 ne
rect 6593 51 6601 83
rect 6631 51 6679 93
rect 6709 83 6734 93
rect 6709 51 6717 83
rect 6833 79 6858 93
rect 6738 51 6772 79
rect 6802 51 6858 79
rect 6888 51 6916 93
rect 4225 14 4319 28
rect 4351 14 4445 28
rect 4805 27 4832 51
rect 4899 29 4931 51
rect 4899 27 4901 29
rect 4929 27 4931 29
rect 4998 27 5025 51
rect 4805 13 4899 27
rect 4931 13 5025 27
rect 5385 27 5412 51
rect 5479 29 5511 51
rect 5479 27 5481 29
rect 5509 27 5511 29
rect 5578 27 5605 51
rect 5385 13 5479 27
rect 5511 13 5605 27
rect 5965 27 5992 51
rect 6059 29 6091 51
rect 6059 27 6061 29
rect 6089 27 6091 29
rect 6158 27 6185 51
rect 5965 13 6059 27
rect 6091 13 6185 27
rect 6545 27 6572 51
rect 6639 29 6671 51
rect 6639 27 6641 29
rect 6669 27 6671 29
rect 6738 27 6765 51
rect 6545 13 6639 27
rect 6671 13 6765 27
rect 88 -72 106 -44
rect 136 -72 154 -44
rect 396 -72 414 -44
rect 444 -72 463 -44
rect 668 -72 686 -44
rect 716 -72 734 -44
rect 976 -72 994 -44
rect 1024 -72 1043 -44
rect 1248 -72 1266 -44
rect 1296 -72 1314 -44
rect 1556 -72 1574 -44
rect 1604 -72 1623 -44
rect 1828 -72 1846 -44
rect 1876 -72 1894 -44
rect 2136 -72 2154 -44
rect 2184 -72 2203 -44
rect 2408 -72 2426 -44
rect 2456 -72 2474 -44
rect 2716 -72 2734 -44
rect 2764 -72 2783 -44
rect 2988 -72 3006 -44
rect 3036 -72 3054 -44
rect 3296 -72 3314 -44
rect 3344 -72 3363 -44
rect 3568 -72 3586 -44
rect 3616 -72 3634 -44
rect 3876 -72 3894 -44
rect 3924 -72 3943 -44
rect 4148 -72 4166 -44
rect 4196 -72 4214 -44
rect 4456 -72 4474 -44
rect 4504 -72 4523 -44
rect 4728 -73 4746 -45
rect 4776 -73 4794 -45
rect 5036 -73 5054 -45
rect 5084 -73 5103 -45
rect 5308 -73 5326 -45
rect 5356 -73 5374 -45
rect 14 -218 42 -176
rect 72 -190 97 -176
rect 196 -186 221 -176
rect 72 -218 128 -190
rect 158 -218 192 -190
tri 206 -193 213 -186 ne
rect 213 -218 221 -186
rect 251 -218 299 -176
rect 329 -186 354 -176
rect 329 -218 337 -186
rect 453 -190 478 -176
rect 358 -218 392 -190
rect 422 -218 478 -190
rect 508 -218 536 -176
rect 594 -218 622 -176
rect 652 -190 677 -176
rect 776 -186 801 -176
rect 652 -218 708 -190
rect 738 -218 772 -190
tri 786 -193 793 -186 ne
rect 793 -218 801 -186
rect 831 -218 879 -176
rect 909 -186 934 -176
rect 909 -218 917 -186
rect 1033 -190 1058 -176
rect 938 -218 972 -190
rect 1002 -218 1058 -190
rect 1088 -218 1116 -176
rect 1174 -218 1202 -176
rect 1232 -190 1257 -176
rect 1356 -186 1381 -176
rect 1232 -218 1288 -190
rect 1318 -218 1352 -190
tri 1366 -193 1373 -186 ne
rect 1373 -218 1381 -186
rect 1411 -218 1459 -176
rect 1489 -186 1514 -176
rect 1489 -218 1497 -186
rect 1613 -190 1638 -176
rect 1518 -218 1552 -190
rect 1582 -218 1638 -190
rect 1668 -218 1696 -176
rect 1754 -218 1782 -176
rect 1812 -190 1837 -176
rect 1936 -186 1961 -176
rect 1812 -218 1868 -190
rect 1898 -218 1932 -190
tri 1946 -193 1953 -186 ne
rect 1953 -218 1961 -186
rect 1991 -218 2039 -176
rect 2069 -186 2094 -176
rect 2069 -218 2077 -186
rect 2193 -190 2218 -176
rect 2098 -218 2132 -190
rect 2162 -218 2218 -190
rect 2248 -218 2276 -176
rect 2334 -218 2362 -176
rect 2392 -190 2417 -176
rect 2516 -186 2541 -176
rect 2392 -218 2448 -190
rect 2478 -218 2512 -190
tri 2526 -193 2533 -186 ne
rect 2533 -218 2541 -186
rect 2571 -218 2619 -176
rect 2649 -186 2674 -176
rect 2649 -218 2657 -186
rect 2773 -190 2798 -176
rect 2678 -218 2712 -190
rect 2742 -218 2798 -190
rect 2828 -218 2856 -176
rect 2914 -218 2942 -176
rect 2972 -190 2997 -176
rect 3096 -186 3121 -176
rect 2972 -218 3028 -190
rect 3058 -218 3092 -190
tri 3106 -193 3113 -186 ne
rect 3113 -218 3121 -186
rect 3151 -218 3199 -176
rect 3229 -186 3254 -176
rect 3229 -218 3237 -186
rect 3353 -190 3378 -176
rect 3258 -218 3292 -190
rect 3322 -218 3378 -190
rect 3408 -218 3436 -176
rect 3494 -218 3522 -176
rect 3552 -190 3577 -176
rect 3676 -186 3701 -176
rect 3552 -218 3608 -190
rect 3638 -218 3672 -190
tri 3686 -193 3693 -186 ne
rect 3693 -218 3701 -186
rect 3731 -218 3779 -176
rect 3809 -186 3834 -176
rect 3809 -218 3817 -186
rect 3933 -190 3958 -176
rect 3838 -218 3872 -190
rect 3902 -218 3958 -190
rect 3988 -218 4016 -176
rect 4074 -218 4102 -176
rect 4132 -190 4157 -176
rect 4256 -186 4281 -176
rect 4132 -218 4188 -190
rect 4218 -218 4252 -190
tri 4266 -193 4273 -186 ne
rect 4273 -218 4281 -186
rect 4311 -218 4359 -176
rect 4389 -186 4414 -176
rect 4389 -218 4397 -186
rect 4513 -190 4538 -176
rect 4418 -218 4452 -190
rect 4482 -218 4538 -190
rect 4568 -218 4596 -176
rect 5616 -73 5634 -45
rect 5664 -73 5683 -45
rect 5888 -73 5906 -45
rect 5936 -73 5954 -45
rect 6196 -73 6214 -45
rect 6244 -73 6263 -45
rect 6468 -73 6486 -45
rect 6516 -73 6534 -45
rect 6776 -73 6794 -45
rect 6824 -73 6843 -45
rect 165 -242 192 -218
rect 259 -240 291 -218
rect 259 -242 261 -240
rect 289 -242 291 -240
rect 358 -242 385 -218
rect 165 -256 259 -242
rect 291 -256 385 -242
rect 745 -242 772 -218
rect 839 -240 871 -218
rect 839 -242 841 -240
rect 869 -242 871 -240
rect 938 -242 965 -218
rect 745 -256 839 -242
rect 871 -256 965 -242
rect 1325 -242 1352 -218
rect 1419 -240 1451 -218
rect 1419 -242 1421 -240
rect 1449 -242 1451 -240
rect 1518 -242 1545 -218
rect 1325 -256 1419 -242
rect 1451 -256 1545 -242
rect 1905 -242 1932 -218
rect 1999 -240 2031 -218
rect 1999 -242 2001 -240
rect 2029 -242 2031 -240
rect 2098 -242 2125 -218
rect 1905 -256 1999 -242
rect 2031 -256 2125 -242
rect 2485 -242 2512 -218
rect 2579 -240 2611 -218
rect 2579 -242 2581 -240
rect 2609 -242 2611 -240
rect 2678 -242 2705 -218
rect 2485 -256 2579 -242
rect 2611 -256 2705 -242
rect 3065 -242 3092 -218
rect 3159 -240 3191 -218
rect 3159 -242 3161 -240
rect 3189 -242 3191 -240
rect 3258 -242 3285 -218
rect 3065 -256 3159 -242
rect 3191 -256 3285 -242
rect 3645 -242 3672 -218
rect 3739 -240 3771 -218
rect 3739 -242 3741 -240
rect 3769 -242 3771 -240
rect 3838 -242 3865 -218
rect 3645 -256 3739 -242
rect 3771 -256 3865 -242
rect 4225 -242 4252 -218
rect 4319 -240 4351 -218
rect 4319 -242 4321 -240
rect 4349 -242 4351 -240
rect 4418 -242 4445 -218
rect 4654 -219 4682 -177
rect 4712 -191 4737 -177
rect 4836 -187 4861 -177
rect 4712 -219 4768 -191
rect 4798 -219 4832 -191
tri 4846 -194 4853 -187 ne
rect 4853 -219 4861 -187
rect 4891 -219 4939 -177
rect 4969 -187 4994 -177
rect 4969 -219 4977 -187
rect 5093 -191 5118 -177
rect 4998 -219 5032 -191
rect 5062 -219 5118 -191
rect 5148 -219 5176 -177
rect 5234 -219 5262 -177
rect 5292 -191 5317 -177
rect 5416 -187 5441 -177
rect 5292 -219 5348 -191
rect 5378 -219 5412 -191
tri 5426 -194 5433 -187 ne
rect 5433 -219 5441 -187
rect 5471 -219 5519 -177
rect 5549 -187 5574 -177
rect 5549 -219 5557 -187
rect 5673 -191 5698 -177
rect 5578 -219 5612 -191
rect 5642 -219 5698 -191
rect 5728 -219 5756 -177
rect 5814 -219 5842 -177
rect 5872 -191 5897 -177
rect 5996 -187 6021 -177
rect 5872 -219 5928 -191
rect 5958 -219 5992 -191
tri 6006 -194 6013 -187 ne
rect 6013 -219 6021 -187
rect 6051 -219 6099 -177
rect 6129 -187 6154 -177
rect 6129 -219 6137 -187
rect 6253 -191 6278 -177
rect 6158 -219 6192 -191
rect 6222 -219 6278 -191
rect 6308 -219 6336 -177
rect 6394 -219 6422 -177
rect 6452 -191 6477 -177
rect 6576 -187 6601 -177
rect 6452 -219 6508 -191
rect 6538 -219 6572 -191
tri 6586 -194 6593 -187 ne
rect 6593 -219 6601 -187
rect 6631 -219 6679 -177
rect 6709 -187 6734 -177
rect 6709 -219 6717 -187
rect 6833 -191 6858 -177
rect 6738 -219 6772 -191
rect 6802 -219 6858 -191
rect 6888 -219 6916 -177
rect 4225 -256 4319 -242
rect 4351 -256 4445 -242
rect 4805 -243 4832 -219
rect 4899 -241 4931 -219
rect 4899 -243 4901 -241
rect 4929 -243 4931 -241
rect 4998 -243 5025 -219
rect 4805 -257 4899 -243
rect 4931 -257 5025 -243
rect 5385 -243 5412 -219
rect 5479 -241 5511 -219
rect 5479 -243 5481 -241
rect 5509 -243 5511 -241
rect 5578 -243 5605 -219
rect 5385 -257 5479 -243
rect 5511 -257 5605 -243
rect 5965 -243 5992 -219
rect 6059 -241 6091 -219
rect 6059 -243 6061 -241
rect 6089 -243 6091 -241
rect 6158 -243 6185 -219
rect 5965 -257 6059 -243
rect 6091 -257 6185 -243
rect 6545 -243 6572 -219
rect 6639 -241 6671 -219
rect 6639 -243 6641 -241
rect 6669 -243 6671 -241
rect 6738 -243 6765 -219
rect 6545 -257 6639 -243
rect 6671 -257 6765 -243
rect 88 -342 106 -314
rect 136 -342 154 -314
rect 396 -342 414 -314
rect 444 -342 463 -314
rect 668 -342 686 -314
rect 716 -342 734 -314
rect 976 -342 994 -314
rect 1024 -342 1043 -314
rect 1248 -342 1266 -314
rect 1296 -342 1314 -314
rect 1556 -342 1574 -314
rect 1604 -342 1623 -314
rect 1828 -342 1846 -314
rect 1876 -342 1894 -314
rect 2136 -342 2154 -314
rect 2184 -342 2203 -314
rect 2408 -342 2426 -314
rect 2456 -342 2474 -314
rect 2716 -342 2734 -314
rect 2764 -342 2783 -314
rect 2988 -342 3006 -314
rect 3036 -342 3054 -314
rect 3296 -342 3314 -314
rect 3344 -342 3363 -314
rect 3568 -342 3586 -314
rect 3616 -342 3634 -314
rect 3876 -342 3894 -314
rect 3924 -342 3943 -314
rect 4148 -342 4166 -314
rect 4196 -342 4214 -314
rect 4456 -342 4474 -314
rect 4504 -342 4523 -314
rect 4728 -343 4746 -315
rect 4776 -343 4794 -315
rect 5036 -343 5054 -315
rect 5084 -343 5103 -315
rect 5308 -343 5326 -315
rect 5356 -343 5374 -315
rect 14 -488 42 -446
rect 72 -460 97 -446
rect 196 -456 221 -446
rect 72 -488 128 -460
rect 158 -488 192 -460
tri 206 -463 213 -456 ne
rect 213 -488 221 -456
rect 251 -488 299 -446
rect 329 -456 354 -446
rect 329 -488 337 -456
rect 453 -460 478 -446
rect 358 -488 392 -460
rect 422 -488 478 -460
rect 508 -488 536 -446
rect 594 -488 622 -446
rect 652 -460 677 -446
rect 776 -456 801 -446
rect 652 -488 708 -460
rect 738 -488 772 -460
tri 786 -463 793 -456 ne
rect 793 -488 801 -456
rect 831 -488 879 -446
rect 909 -456 934 -446
rect 909 -488 917 -456
rect 1033 -460 1058 -446
rect 938 -488 972 -460
rect 1002 -488 1058 -460
rect 1088 -488 1116 -446
rect 1174 -488 1202 -446
rect 1232 -460 1257 -446
rect 1356 -456 1381 -446
rect 1232 -488 1288 -460
rect 1318 -488 1352 -460
tri 1366 -463 1373 -456 ne
rect 1373 -488 1381 -456
rect 1411 -488 1459 -446
rect 1489 -456 1514 -446
rect 1489 -488 1497 -456
rect 1613 -460 1638 -446
rect 1518 -488 1552 -460
rect 1582 -488 1638 -460
rect 1668 -488 1696 -446
rect 1754 -488 1782 -446
rect 1812 -460 1837 -446
rect 1936 -456 1961 -446
rect 1812 -488 1868 -460
rect 1898 -488 1932 -460
tri 1946 -463 1953 -456 ne
rect 1953 -488 1961 -456
rect 1991 -488 2039 -446
rect 2069 -456 2094 -446
rect 2069 -488 2077 -456
rect 2193 -460 2218 -446
rect 2098 -488 2132 -460
rect 2162 -488 2218 -460
rect 2248 -488 2276 -446
rect 2334 -488 2362 -446
rect 2392 -460 2417 -446
rect 2516 -456 2541 -446
rect 2392 -488 2448 -460
rect 2478 -488 2512 -460
tri 2526 -463 2533 -456 ne
rect 2533 -488 2541 -456
rect 2571 -488 2619 -446
rect 2649 -456 2674 -446
rect 2649 -488 2657 -456
rect 2773 -460 2798 -446
rect 2678 -488 2712 -460
rect 2742 -488 2798 -460
rect 2828 -488 2856 -446
rect 2914 -488 2942 -446
rect 2972 -460 2997 -446
rect 3096 -456 3121 -446
rect 2972 -488 3028 -460
rect 3058 -488 3092 -460
tri 3106 -463 3113 -456 ne
rect 3113 -488 3121 -456
rect 3151 -488 3199 -446
rect 3229 -456 3254 -446
rect 3229 -488 3237 -456
rect 3353 -460 3378 -446
rect 3258 -488 3292 -460
rect 3322 -488 3378 -460
rect 3408 -488 3436 -446
rect 3494 -488 3522 -446
rect 3552 -460 3577 -446
rect 3676 -456 3701 -446
rect 3552 -488 3608 -460
rect 3638 -488 3672 -460
tri 3686 -463 3693 -456 ne
rect 3693 -488 3701 -456
rect 3731 -488 3779 -446
rect 3809 -456 3834 -446
rect 3809 -488 3817 -456
rect 3933 -460 3958 -446
rect 3838 -488 3872 -460
rect 3902 -488 3958 -460
rect 3988 -488 4016 -446
rect 4074 -488 4102 -446
rect 4132 -460 4157 -446
rect 4256 -456 4281 -446
rect 4132 -488 4188 -460
rect 4218 -488 4252 -460
tri 4266 -463 4273 -456 ne
rect 4273 -488 4281 -456
rect 4311 -488 4359 -446
rect 4389 -456 4414 -446
rect 4389 -488 4397 -456
rect 4513 -460 4538 -446
rect 4418 -488 4452 -460
rect 4482 -488 4538 -460
rect 4568 -488 4596 -446
rect 5616 -343 5634 -315
rect 5664 -343 5683 -315
rect 5888 -343 5906 -315
rect 5936 -343 5954 -315
rect 6196 -343 6214 -315
rect 6244 -343 6263 -315
rect 6468 -343 6486 -315
rect 6516 -343 6534 -315
rect 6776 -343 6794 -315
rect 6824 -343 6843 -315
rect 165 -512 192 -488
rect 259 -510 291 -488
rect 259 -512 261 -510
rect 289 -512 291 -510
rect 358 -512 385 -488
rect 165 -526 259 -512
rect 291 -526 385 -512
rect 745 -512 772 -488
rect 839 -510 871 -488
rect 839 -512 841 -510
rect 869 -512 871 -510
rect 938 -512 965 -488
rect 745 -526 839 -512
rect 871 -526 965 -512
rect 1325 -512 1352 -488
rect 1419 -510 1451 -488
rect 1419 -512 1421 -510
rect 1449 -512 1451 -510
rect 1518 -512 1545 -488
rect 1325 -526 1419 -512
rect 1451 -526 1545 -512
rect 1905 -512 1932 -488
rect 1999 -510 2031 -488
rect 1999 -512 2001 -510
rect 2029 -512 2031 -510
rect 2098 -512 2125 -488
rect 1905 -526 1999 -512
rect 2031 -526 2125 -512
rect 2485 -512 2512 -488
rect 2579 -510 2611 -488
rect 2579 -512 2581 -510
rect 2609 -512 2611 -510
rect 2678 -512 2705 -488
rect 2485 -526 2579 -512
rect 2611 -526 2705 -512
rect 3065 -512 3092 -488
rect 3159 -510 3191 -488
rect 3159 -512 3161 -510
rect 3189 -512 3191 -510
rect 3258 -512 3285 -488
rect 3065 -526 3159 -512
rect 3191 -526 3285 -512
rect 3645 -512 3672 -488
rect 3739 -510 3771 -488
rect 3739 -512 3741 -510
rect 3769 -512 3771 -510
rect 3838 -512 3865 -488
rect 3645 -526 3739 -512
rect 3771 -526 3865 -512
rect 4225 -512 4252 -488
rect 4319 -510 4351 -488
rect 4319 -512 4321 -510
rect 4349 -512 4351 -510
rect 4418 -512 4445 -488
rect 4654 -489 4682 -447
rect 4712 -461 4737 -447
rect 4836 -457 4861 -447
rect 4712 -489 4768 -461
rect 4798 -489 4832 -461
tri 4846 -464 4853 -457 ne
rect 4853 -489 4861 -457
rect 4891 -489 4939 -447
rect 4969 -457 4994 -447
rect 4969 -489 4977 -457
rect 5093 -461 5118 -447
rect 4998 -489 5032 -461
rect 5062 -489 5118 -461
rect 5148 -489 5176 -447
rect 5234 -489 5262 -447
rect 5292 -461 5317 -447
rect 5416 -457 5441 -447
rect 5292 -489 5348 -461
rect 5378 -489 5412 -461
tri 5426 -464 5433 -457 ne
rect 5433 -489 5441 -457
rect 5471 -489 5519 -447
rect 5549 -457 5574 -447
rect 5549 -489 5557 -457
rect 5673 -461 5698 -447
rect 5578 -489 5612 -461
rect 5642 -489 5698 -461
rect 5728 -489 5756 -447
rect 5814 -489 5842 -447
rect 5872 -461 5897 -447
rect 5996 -457 6021 -447
rect 5872 -489 5928 -461
rect 5958 -489 5992 -461
tri 6006 -464 6013 -457 ne
rect 6013 -489 6021 -457
rect 6051 -489 6099 -447
rect 6129 -457 6154 -447
rect 6129 -489 6137 -457
rect 6253 -461 6278 -447
rect 6158 -489 6192 -461
rect 6222 -489 6278 -461
rect 6308 -489 6336 -447
rect 6394 -489 6422 -447
rect 6452 -461 6477 -447
rect 6576 -457 6601 -447
rect 6452 -489 6508 -461
rect 6538 -489 6572 -461
tri 6586 -464 6593 -457 ne
rect 6593 -489 6601 -457
rect 6631 -489 6679 -447
rect 6709 -457 6734 -447
rect 6709 -489 6717 -457
rect 6833 -461 6858 -447
rect 6738 -489 6772 -461
rect 6802 -489 6858 -461
rect 6888 -489 6916 -447
rect 4225 -526 4319 -512
rect 4351 -526 4445 -512
rect 4805 -513 4832 -489
rect 4899 -511 4931 -489
rect 4899 -513 4901 -511
rect 4929 -513 4931 -511
rect 4998 -513 5025 -489
rect 4805 -527 4899 -513
rect 4931 -527 5025 -513
rect 5385 -513 5412 -489
rect 5479 -511 5511 -489
rect 5479 -513 5481 -511
rect 5509 -513 5511 -511
rect 5578 -513 5605 -489
rect 5385 -527 5479 -513
rect 5511 -527 5605 -513
rect 5965 -513 5992 -489
rect 6059 -511 6091 -489
rect 6059 -513 6061 -511
rect 6089 -513 6091 -511
rect 6158 -513 6185 -489
rect 5965 -527 6059 -513
rect 6091 -527 6185 -513
rect 6545 -513 6572 -489
rect 6639 -511 6671 -489
rect 6639 -513 6641 -511
rect 6669 -513 6671 -511
rect 6738 -513 6765 -489
rect 6545 -527 6639 -513
rect 6671 -527 6765 -513
rect 88 -612 106 -584
rect 136 -612 154 -584
rect 396 -612 414 -584
rect 444 -612 463 -584
rect 668 -612 686 -584
rect 716 -612 734 -584
rect 976 -612 994 -584
rect 1024 -612 1043 -584
rect 1248 -612 1266 -584
rect 1296 -612 1314 -584
rect 1556 -612 1574 -584
rect 1604 -612 1623 -584
rect 1828 -612 1846 -584
rect 1876 -612 1894 -584
rect 2136 -612 2154 -584
rect 2184 -612 2203 -584
rect 2408 -612 2426 -584
rect 2456 -612 2474 -584
rect 2716 -612 2734 -584
rect 2764 -612 2783 -584
rect 2988 -612 3006 -584
rect 3036 -612 3054 -584
rect 3296 -612 3314 -584
rect 3344 -612 3363 -584
rect 3568 -612 3586 -584
rect 3616 -612 3634 -584
rect 3876 -612 3894 -584
rect 3924 -612 3943 -584
rect 4148 -612 4166 -584
rect 4196 -612 4214 -584
rect 4456 -612 4474 -584
rect 4504 -612 4523 -584
rect 4728 -613 4746 -585
rect 4776 -613 4794 -585
rect 5036 -613 5054 -585
rect 5084 -613 5103 -585
rect 5308 -613 5326 -585
rect 5356 -613 5374 -585
rect 14 -758 42 -716
rect 72 -730 97 -716
rect 196 -726 221 -716
rect 72 -758 128 -730
rect 158 -758 192 -730
tri 206 -733 213 -726 ne
rect 213 -758 221 -726
rect 251 -758 299 -716
rect 329 -726 354 -716
rect 329 -758 337 -726
rect 453 -730 478 -716
rect 358 -758 392 -730
rect 422 -758 478 -730
rect 508 -758 536 -716
rect 594 -758 622 -716
rect 652 -730 677 -716
rect 776 -726 801 -716
rect 652 -758 708 -730
rect 738 -758 772 -730
tri 786 -733 793 -726 ne
rect 793 -758 801 -726
rect 831 -758 879 -716
rect 909 -726 934 -716
rect 909 -758 917 -726
rect 1033 -730 1058 -716
rect 938 -758 972 -730
rect 1002 -758 1058 -730
rect 1088 -758 1116 -716
rect 1174 -758 1202 -716
rect 1232 -730 1257 -716
rect 1356 -726 1381 -716
rect 1232 -758 1288 -730
rect 1318 -758 1352 -730
tri 1366 -733 1373 -726 ne
rect 1373 -758 1381 -726
rect 1411 -758 1459 -716
rect 1489 -726 1514 -716
rect 1489 -758 1497 -726
rect 1613 -730 1638 -716
rect 1518 -758 1552 -730
rect 1582 -758 1638 -730
rect 1668 -758 1696 -716
rect 1754 -758 1782 -716
rect 1812 -730 1837 -716
rect 1936 -726 1961 -716
rect 1812 -758 1868 -730
rect 1898 -758 1932 -730
tri 1946 -733 1953 -726 ne
rect 1953 -758 1961 -726
rect 1991 -758 2039 -716
rect 2069 -726 2094 -716
rect 2069 -758 2077 -726
rect 2193 -730 2218 -716
rect 2098 -758 2132 -730
rect 2162 -758 2218 -730
rect 2248 -758 2276 -716
rect 2334 -758 2362 -716
rect 2392 -730 2417 -716
rect 2516 -726 2541 -716
rect 2392 -758 2448 -730
rect 2478 -758 2512 -730
tri 2526 -733 2533 -726 ne
rect 2533 -758 2541 -726
rect 2571 -758 2619 -716
rect 2649 -726 2674 -716
rect 2649 -758 2657 -726
rect 2773 -730 2798 -716
rect 2678 -758 2712 -730
rect 2742 -758 2798 -730
rect 2828 -758 2856 -716
rect 2914 -758 2942 -716
rect 2972 -730 2997 -716
rect 3096 -726 3121 -716
rect 2972 -758 3028 -730
rect 3058 -758 3092 -730
tri 3106 -733 3113 -726 ne
rect 3113 -758 3121 -726
rect 3151 -758 3199 -716
rect 3229 -726 3254 -716
rect 3229 -758 3237 -726
rect 3353 -730 3378 -716
rect 3258 -758 3292 -730
rect 3322 -758 3378 -730
rect 3408 -758 3436 -716
rect 3494 -758 3522 -716
rect 3552 -730 3577 -716
rect 3676 -726 3701 -716
rect 3552 -758 3608 -730
rect 3638 -758 3672 -730
tri 3686 -733 3693 -726 ne
rect 3693 -758 3701 -726
rect 3731 -758 3779 -716
rect 3809 -726 3834 -716
rect 3809 -758 3817 -726
rect 3933 -730 3958 -716
rect 3838 -758 3872 -730
rect 3902 -758 3958 -730
rect 3988 -758 4016 -716
rect 4074 -758 4102 -716
rect 4132 -730 4157 -716
rect 4256 -726 4281 -716
rect 4132 -758 4188 -730
rect 4218 -758 4252 -730
tri 4266 -733 4273 -726 ne
rect 4273 -758 4281 -726
rect 4311 -758 4359 -716
rect 4389 -726 4414 -716
rect 4389 -758 4397 -726
rect 4513 -730 4538 -716
rect 4418 -758 4452 -730
rect 4482 -758 4538 -730
rect 4568 -758 4596 -716
rect 5616 -613 5634 -585
rect 5664 -613 5683 -585
rect 5888 -613 5906 -585
rect 5936 -613 5954 -585
rect 6196 -613 6214 -585
rect 6244 -613 6263 -585
rect 6468 -613 6486 -585
rect 6516 -613 6534 -585
rect 6776 -613 6794 -585
rect 6824 -613 6843 -585
rect 165 -782 192 -758
rect 259 -780 291 -758
rect 259 -782 261 -780
rect 289 -782 291 -780
rect 358 -782 385 -758
rect 165 -796 259 -782
rect 291 -796 385 -782
rect 745 -782 772 -758
rect 839 -780 871 -758
rect 839 -782 841 -780
rect 869 -782 871 -780
rect 938 -782 965 -758
rect 745 -796 839 -782
rect 871 -796 965 -782
rect 1325 -782 1352 -758
rect 1419 -780 1451 -758
rect 1419 -782 1421 -780
rect 1449 -782 1451 -780
rect 1518 -782 1545 -758
rect 1325 -796 1419 -782
rect 1451 -796 1545 -782
rect 1905 -782 1932 -758
rect 1999 -780 2031 -758
rect 1999 -782 2001 -780
rect 2029 -782 2031 -780
rect 2098 -782 2125 -758
rect 1905 -796 1999 -782
rect 2031 -796 2125 -782
rect 2485 -782 2512 -758
rect 2579 -780 2611 -758
rect 2579 -782 2581 -780
rect 2609 -782 2611 -780
rect 2678 -782 2705 -758
rect 2485 -796 2579 -782
rect 2611 -796 2705 -782
rect 3065 -782 3092 -758
rect 3159 -780 3191 -758
rect 3159 -782 3161 -780
rect 3189 -782 3191 -780
rect 3258 -782 3285 -758
rect 3065 -796 3159 -782
rect 3191 -796 3285 -782
rect 3645 -782 3672 -758
rect 3739 -780 3771 -758
rect 3739 -782 3741 -780
rect 3769 -782 3771 -780
rect 3838 -782 3865 -758
rect 3645 -796 3739 -782
rect 3771 -796 3865 -782
rect 4225 -782 4252 -758
rect 4319 -780 4351 -758
rect 4319 -782 4321 -780
rect 4349 -782 4351 -780
rect 4418 -782 4445 -758
rect 4654 -759 4682 -717
rect 4712 -731 4737 -717
rect 4836 -727 4861 -717
rect 4712 -759 4768 -731
rect 4798 -759 4832 -731
tri 4846 -734 4853 -727 ne
rect 4853 -759 4861 -727
rect 4891 -759 4939 -717
rect 4969 -727 4994 -717
rect 4969 -759 4977 -727
rect 5093 -731 5118 -717
rect 4998 -759 5032 -731
rect 5062 -759 5118 -731
rect 5148 -759 5176 -717
rect 5234 -759 5262 -717
rect 5292 -731 5317 -717
rect 5416 -727 5441 -717
rect 5292 -759 5348 -731
rect 5378 -759 5412 -731
tri 5426 -734 5433 -727 ne
rect 5433 -759 5441 -727
rect 5471 -759 5519 -717
rect 5549 -727 5574 -717
rect 5549 -759 5557 -727
rect 5673 -731 5698 -717
rect 5578 -759 5612 -731
rect 5642 -759 5698 -731
rect 5728 -759 5756 -717
rect 5814 -759 5842 -717
rect 5872 -731 5897 -717
rect 5996 -727 6021 -717
rect 5872 -759 5928 -731
rect 5958 -759 5992 -731
tri 6006 -734 6013 -727 ne
rect 6013 -759 6021 -727
rect 6051 -759 6099 -717
rect 6129 -727 6154 -717
rect 6129 -759 6137 -727
rect 6253 -731 6278 -717
rect 6158 -759 6192 -731
rect 6222 -759 6278 -731
rect 6308 -759 6336 -717
rect 6394 -759 6422 -717
rect 6452 -731 6477 -717
rect 6576 -727 6601 -717
rect 6452 -759 6508 -731
rect 6538 -759 6572 -731
tri 6586 -734 6593 -727 ne
rect 6593 -759 6601 -727
rect 6631 -759 6679 -717
rect 6709 -727 6734 -717
rect 6709 -759 6717 -727
rect 6833 -731 6858 -717
rect 6738 -759 6772 -731
rect 6802 -759 6858 -731
rect 6888 -759 6916 -717
rect 4225 -796 4319 -782
rect 4351 -796 4445 -782
rect 4805 -783 4832 -759
rect 4899 -781 4931 -759
rect 4899 -783 4901 -781
rect 4929 -783 4931 -781
rect 4998 -783 5025 -759
rect 4805 -797 4899 -783
rect 4931 -797 5025 -783
rect 5385 -783 5412 -759
rect 5479 -781 5511 -759
rect 5479 -783 5481 -781
rect 5509 -783 5511 -781
rect 5578 -783 5605 -759
rect 5385 -797 5479 -783
rect 5511 -797 5605 -783
rect 5965 -783 5992 -759
rect 6059 -781 6091 -759
rect 6059 -783 6061 -781
rect 6089 -783 6091 -781
rect 6158 -783 6185 -759
rect 5965 -797 6059 -783
rect 6091 -797 6185 -783
rect 6545 -783 6572 -759
rect 6639 -781 6671 -759
rect 6639 -783 6641 -781
rect 6669 -783 6671 -781
rect 6738 -783 6765 -759
rect 6545 -797 6639 -783
rect 6671 -797 6765 -783
rect 88 -882 106 -854
rect 136 -882 154 -854
rect 396 -882 414 -854
rect 444 -882 463 -854
rect 668 -882 686 -854
rect 716 -882 734 -854
rect 976 -882 994 -854
rect 1024 -882 1043 -854
rect 1248 -882 1266 -854
rect 1296 -882 1314 -854
rect 1556 -882 1574 -854
rect 1604 -882 1623 -854
rect 1828 -882 1846 -854
rect 1876 -882 1894 -854
rect 2136 -882 2154 -854
rect 2184 -882 2203 -854
rect 2408 -882 2426 -854
rect 2456 -882 2474 -854
rect 2716 -882 2734 -854
rect 2764 -882 2783 -854
rect 2988 -882 3006 -854
rect 3036 -882 3054 -854
rect 3296 -882 3314 -854
rect 3344 -882 3363 -854
rect 3568 -882 3586 -854
rect 3616 -882 3634 -854
rect 3876 -882 3894 -854
rect 3924 -882 3943 -854
rect 4148 -882 4166 -854
rect 4196 -882 4214 -854
rect 4456 -882 4474 -854
rect 4504 -882 4523 -854
rect 4728 -883 4746 -855
rect 4776 -883 4794 -855
rect 5036 -883 5054 -855
rect 5084 -883 5103 -855
rect 5308 -883 5326 -855
rect 5356 -883 5374 -855
rect 14 -1028 42 -986
rect 72 -1000 97 -986
rect 196 -996 221 -986
rect 72 -1028 128 -1000
rect 158 -1028 192 -1000
tri 206 -1003 213 -996 ne
rect 213 -1028 221 -996
rect 251 -1028 299 -986
rect 329 -996 354 -986
rect 329 -1028 337 -996
rect 453 -1000 478 -986
rect 358 -1028 392 -1000
rect 422 -1028 478 -1000
rect 508 -1028 536 -986
rect 594 -1028 622 -986
rect 652 -1000 677 -986
rect 776 -996 801 -986
rect 652 -1028 708 -1000
rect 738 -1028 772 -1000
tri 786 -1003 793 -996 ne
rect 793 -1028 801 -996
rect 831 -1028 879 -986
rect 909 -996 934 -986
rect 909 -1028 917 -996
rect 1033 -1000 1058 -986
rect 938 -1028 972 -1000
rect 1002 -1028 1058 -1000
rect 1088 -1028 1116 -986
rect 1174 -1028 1202 -986
rect 1232 -1000 1257 -986
rect 1356 -996 1381 -986
rect 1232 -1028 1288 -1000
rect 1318 -1028 1352 -1000
tri 1366 -1003 1373 -996 ne
rect 1373 -1028 1381 -996
rect 1411 -1028 1459 -986
rect 1489 -996 1514 -986
rect 1489 -1028 1497 -996
rect 1613 -1000 1638 -986
rect 1518 -1028 1552 -1000
rect 1582 -1028 1638 -1000
rect 1668 -1028 1696 -986
rect 1754 -1028 1782 -986
rect 1812 -1000 1837 -986
rect 1936 -996 1961 -986
rect 1812 -1028 1868 -1000
rect 1898 -1028 1932 -1000
tri 1946 -1003 1953 -996 ne
rect 1953 -1028 1961 -996
rect 1991 -1028 2039 -986
rect 2069 -996 2094 -986
rect 2069 -1028 2077 -996
rect 2193 -1000 2218 -986
rect 2098 -1028 2132 -1000
rect 2162 -1028 2218 -1000
rect 2248 -1028 2276 -986
rect 2334 -1028 2362 -986
rect 2392 -1000 2417 -986
rect 2516 -996 2541 -986
rect 2392 -1028 2448 -1000
rect 2478 -1028 2512 -1000
tri 2526 -1003 2533 -996 ne
rect 2533 -1028 2541 -996
rect 2571 -1028 2619 -986
rect 2649 -996 2674 -986
rect 2649 -1028 2657 -996
rect 2773 -1000 2798 -986
rect 2678 -1028 2712 -1000
rect 2742 -1028 2798 -1000
rect 2828 -1028 2856 -986
rect 2914 -1028 2942 -986
rect 2972 -1000 2997 -986
rect 3096 -996 3121 -986
rect 2972 -1028 3028 -1000
rect 3058 -1028 3092 -1000
tri 3106 -1003 3113 -996 ne
rect 3113 -1028 3121 -996
rect 3151 -1028 3199 -986
rect 3229 -996 3254 -986
rect 3229 -1028 3237 -996
rect 3353 -1000 3378 -986
rect 3258 -1028 3292 -1000
rect 3322 -1028 3378 -1000
rect 3408 -1028 3436 -986
rect 3494 -1028 3522 -986
rect 3552 -1000 3577 -986
rect 3676 -996 3701 -986
rect 3552 -1028 3608 -1000
rect 3638 -1028 3672 -1000
tri 3686 -1003 3693 -996 ne
rect 3693 -1028 3701 -996
rect 3731 -1028 3779 -986
rect 3809 -996 3834 -986
rect 3809 -1028 3817 -996
rect 3933 -1000 3958 -986
rect 3838 -1028 3872 -1000
rect 3902 -1028 3958 -1000
rect 3988 -1028 4016 -986
rect 4074 -1028 4102 -986
rect 4132 -1000 4157 -986
rect 4256 -996 4281 -986
rect 4132 -1028 4188 -1000
rect 4218 -1028 4252 -1000
tri 4266 -1003 4273 -996 ne
rect 4273 -1028 4281 -996
rect 4311 -1028 4359 -986
rect 4389 -996 4414 -986
rect 4389 -1028 4397 -996
rect 4513 -1000 4538 -986
rect 4418 -1028 4452 -1000
rect 4482 -1028 4538 -1000
rect 4568 -1028 4596 -986
rect 5616 -883 5634 -855
rect 5664 -883 5683 -855
rect 5888 -883 5906 -855
rect 5936 -883 5954 -855
rect 6196 -883 6214 -855
rect 6244 -883 6263 -855
rect 6468 -883 6486 -855
rect 6516 -883 6534 -855
rect 6776 -883 6794 -855
rect 6824 -883 6843 -855
rect 165 -1052 192 -1028
rect 259 -1050 291 -1028
rect 259 -1052 261 -1050
rect 289 -1052 291 -1050
rect 358 -1052 385 -1028
rect 165 -1066 259 -1052
rect 291 -1066 385 -1052
rect 745 -1052 772 -1028
rect 839 -1050 871 -1028
rect 839 -1052 841 -1050
rect 869 -1052 871 -1050
rect 938 -1052 965 -1028
rect 745 -1066 839 -1052
rect 871 -1066 965 -1052
rect 1325 -1052 1352 -1028
rect 1419 -1050 1451 -1028
rect 1419 -1052 1421 -1050
rect 1449 -1052 1451 -1050
rect 1518 -1052 1545 -1028
rect 1325 -1066 1419 -1052
rect 1451 -1066 1545 -1052
rect 1905 -1052 1932 -1028
rect 1999 -1050 2031 -1028
rect 1999 -1052 2001 -1050
rect 2029 -1052 2031 -1050
rect 2098 -1052 2125 -1028
rect 1905 -1066 1999 -1052
rect 2031 -1066 2125 -1052
rect 2485 -1052 2512 -1028
rect 2579 -1050 2611 -1028
rect 2579 -1052 2581 -1050
rect 2609 -1052 2611 -1050
rect 2678 -1052 2705 -1028
rect 2485 -1066 2579 -1052
rect 2611 -1066 2705 -1052
rect 3065 -1052 3092 -1028
rect 3159 -1050 3191 -1028
rect 3159 -1052 3161 -1050
rect 3189 -1052 3191 -1050
rect 3258 -1052 3285 -1028
rect 3065 -1066 3159 -1052
rect 3191 -1066 3285 -1052
rect 3645 -1052 3672 -1028
rect 3739 -1050 3771 -1028
rect 3739 -1052 3741 -1050
rect 3769 -1052 3771 -1050
rect 3838 -1052 3865 -1028
rect 3645 -1066 3739 -1052
rect 3771 -1066 3865 -1052
rect 4225 -1052 4252 -1028
rect 4319 -1050 4351 -1028
rect 4319 -1052 4321 -1050
rect 4349 -1052 4351 -1050
rect 4418 -1052 4445 -1028
rect 4654 -1029 4682 -987
rect 4712 -1001 4737 -987
rect 4836 -997 4861 -987
rect 4712 -1029 4768 -1001
rect 4798 -1029 4832 -1001
tri 4846 -1004 4853 -997 ne
rect 4853 -1029 4861 -997
rect 4891 -1029 4939 -987
rect 4969 -997 4994 -987
rect 4969 -1029 4977 -997
rect 5093 -1001 5118 -987
rect 4998 -1029 5032 -1001
rect 5062 -1029 5118 -1001
rect 5148 -1029 5176 -987
rect 5234 -1029 5262 -987
rect 5292 -1001 5317 -987
rect 5416 -997 5441 -987
rect 5292 -1029 5348 -1001
rect 5378 -1029 5412 -1001
tri 5426 -1004 5433 -997 ne
rect 5433 -1029 5441 -997
rect 5471 -1029 5519 -987
rect 5549 -997 5574 -987
rect 5549 -1029 5557 -997
rect 5673 -1001 5698 -987
rect 5578 -1029 5612 -1001
rect 5642 -1029 5698 -1001
rect 5728 -1029 5756 -987
rect 5814 -1029 5842 -987
rect 5872 -1001 5897 -987
rect 5996 -997 6021 -987
rect 5872 -1029 5928 -1001
rect 5958 -1029 5992 -1001
tri 6006 -1004 6013 -997 ne
rect 6013 -1029 6021 -997
rect 6051 -1029 6099 -987
rect 6129 -997 6154 -987
rect 6129 -1029 6137 -997
rect 6253 -1001 6278 -987
rect 6158 -1029 6192 -1001
rect 6222 -1029 6278 -1001
rect 6308 -1029 6336 -987
rect 6394 -1029 6422 -987
rect 6452 -1001 6477 -987
rect 6576 -997 6601 -987
rect 6452 -1029 6508 -1001
rect 6538 -1029 6572 -1001
tri 6586 -1004 6593 -997 ne
rect 6593 -1029 6601 -997
rect 6631 -1029 6679 -987
rect 6709 -997 6734 -987
rect 6709 -1029 6717 -997
rect 6833 -1001 6858 -987
rect 6738 -1029 6772 -1001
rect 6802 -1029 6858 -1001
rect 6888 -1029 6916 -987
rect 4225 -1066 4319 -1052
rect 4351 -1066 4445 -1052
rect 4805 -1053 4832 -1029
rect 4899 -1051 4931 -1029
rect 4899 -1053 4901 -1051
rect 4929 -1053 4931 -1051
rect 4998 -1053 5025 -1029
rect 4805 -1067 4899 -1053
rect 4931 -1067 5025 -1053
rect 5385 -1053 5412 -1029
rect 5479 -1051 5511 -1029
rect 5479 -1053 5481 -1051
rect 5509 -1053 5511 -1051
rect 5578 -1053 5605 -1029
rect 5385 -1067 5479 -1053
rect 5511 -1067 5605 -1053
rect 5965 -1053 5992 -1029
rect 6059 -1051 6091 -1029
rect 6059 -1053 6061 -1051
rect 6089 -1053 6091 -1051
rect 6158 -1053 6185 -1029
rect 5965 -1067 6059 -1053
rect 6091 -1067 6185 -1053
rect 6545 -1053 6572 -1029
rect 6639 -1051 6671 -1029
rect 6639 -1053 6641 -1051
rect 6669 -1053 6671 -1051
rect 6738 -1053 6765 -1029
rect 6545 -1067 6639 -1053
rect 6671 -1067 6765 -1053
rect 88 -1152 106 -1124
rect 136 -1152 154 -1124
rect 396 -1152 414 -1124
rect 444 -1152 463 -1124
rect 668 -1152 686 -1124
rect 716 -1152 734 -1124
rect 976 -1152 994 -1124
rect 1024 -1152 1043 -1124
rect 1248 -1152 1266 -1124
rect 1296 -1152 1314 -1124
rect 1556 -1152 1574 -1124
rect 1604 -1152 1623 -1124
rect 1828 -1152 1846 -1124
rect 1876 -1152 1894 -1124
rect 2136 -1152 2154 -1124
rect 2184 -1152 2203 -1124
rect 2408 -1152 2426 -1124
rect 2456 -1152 2474 -1124
rect 2716 -1152 2734 -1124
rect 2764 -1152 2783 -1124
rect 2988 -1152 3006 -1124
rect 3036 -1152 3054 -1124
rect 3296 -1152 3314 -1124
rect 3344 -1152 3363 -1124
rect 3568 -1152 3586 -1124
rect 3616 -1152 3634 -1124
rect 3876 -1152 3894 -1124
rect 3924 -1152 3943 -1124
rect 4148 -1152 4166 -1124
rect 4196 -1152 4214 -1124
rect 4456 -1152 4474 -1124
rect 4504 -1152 4523 -1124
rect 4728 -1153 4746 -1125
rect 4776 -1153 4794 -1125
rect 5036 -1153 5054 -1125
rect 5084 -1153 5103 -1125
rect 5308 -1153 5326 -1125
rect 5356 -1153 5374 -1125
rect 14 -1298 42 -1256
rect 72 -1270 97 -1256
rect 196 -1266 221 -1256
rect 72 -1298 128 -1270
rect 158 -1298 192 -1270
tri 206 -1273 213 -1266 ne
rect 213 -1298 221 -1266
rect 251 -1298 299 -1256
rect 329 -1266 354 -1256
rect 329 -1298 337 -1266
rect 453 -1270 478 -1256
rect 358 -1298 392 -1270
rect 422 -1298 478 -1270
rect 508 -1298 536 -1256
rect 594 -1298 622 -1256
rect 652 -1270 677 -1256
rect 776 -1266 801 -1256
rect 652 -1298 708 -1270
rect 738 -1298 772 -1270
tri 786 -1273 793 -1266 ne
rect 793 -1298 801 -1266
rect 831 -1298 879 -1256
rect 909 -1266 934 -1256
rect 909 -1298 917 -1266
rect 1033 -1270 1058 -1256
rect 938 -1298 972 -1270
rect 1002 -1298 1058 -1270
rect 1088 -1298 1116 -1256
rect 1174 -1298 1202 -1256
rect 1232 -1270 1257 -1256
rect 1356 -1266 1381 -1256
rect 1232 -1298 1288 -1270
rect 1318 -1298 1352 -1270
tri 1366 -1273 1373 -1266 ne
rect 1373 -1298 1381 -1266
rect 1411 -1298 1459 -1256
rect 1489 -1266 1514 -1256
rect 1489 -1298 1497 -1266
rect 1613 -1270 1638 -1256
rect 1518 -1298 1552 -1270
rect 1582 -1298 1638 -1270
rect 1668 -1298 1696 -1256
rect 1754 -1298 1782 -1256
rect 1812 -1270 1837 -1256
rect 1936 -1266 1961 -1256
rect 1812 -1298 1868 -1270
rect 1898 -1298 1932 -1270
tri 1946 -1273 1953 -1266 ne
rect 1953 -1298 1961 -1266
rect 1991 -1298 2039 -1256
rect 2069 -1266 2094 -1256
rect 2069 -1298 2077 -1266
rect 2193 -1270 2218 -1256
rect 2098 -1298 2132 -1270
rect 2162 -1298 2218 -1270
rect 2248 -1298 2276 -1256
rect 2334 -1298 2362 -1256
rect 2392 -1270 2417 -1256
rect 2516 -1266 2541 -1256
rect 2392 -1298 2448 -1270
rect 2478 -1298 2512 -1270
tri 2526 -1273 2533 -1266 ne
rect 2533 -1298 2541 -1266
rect 2571 -1298 2619 -1256
rect 2649 -1266 2674 -1256
rect 2649 -1298 2657 -1266
rect 2773 -1270 2798 -1256
rect 2678 -1298 2712 -1270
rect 2742 -1298 2798 -1270
rect 2828 -1298 2856 -1256
rect 2914 -1298 2942 -1256
rect 2972 -1270 2997 -1256
rect 3096 -1266 3121 -1256
rect 2972 -1298 3028 -1270
rect 3058 -1298 3092 -1270
tri 3106 -1273 3113 -1266 ne
rect 3113 -1298 3121 -1266
rect 3151 -1298 3199 -1256
rect 3229 -1266 3254 -1256
rect 3229 -1298 3237 -1266
rect 3353 -1270 3378 -1256
rect 3258 -1298 3292 -1270
rect 3322 -1298 3378 -1270
rect 3408 -1298 3436 -1256
rect 3494 -1298 3522 -1256
rect 3552 -1270 3577 -1256
rect 3676 -1266 3701 -1256
rect 3552 -1298 3608 -1270
rect 3638 -1298 3672 -1270
tri 3686 -1273 3693 -1266 ne
rect 3693 -1298 3701 -1266
rect 3731 -1298 3779 -1256
rect 3809 -1266 3834 -1256
rect 3809 -1298 3817 -1266
rect 3933 -1270 3958 -1256
rect 3838 -1298 3872 -1270
rect 3902 -1298 3958 -1270
rect 3988 -1298 4016 -1256
rect 4074 -1298 4102 -1256
rect 4132 -1270 4157 -1256
rect 4256 -1266 4281 -1256
rect 4132 -1298 4188 -1270
rect 4218 -1298 4252 -1270
tri 4266 -1273 4273 -1266 ne
rect 4273 -1298 4281 -1266
rect 4311 -1298 4359 -1256
rect 4389 -1266 4414 -1256
rect 4389 -1298 4397 -1266
rect 4513 -1270 4538 -1256
rect 4418 -1298 4452 -1270
rect 4482 -1298 4538 -1270
rect 4568 -1298 4596 -1256
rect 5616 -1153 5634 -1125
rect 5664 -1153 5683 -1125
rect 5888 -1153 5906 -1125
rect 5936 -1153 5954 -1125
rect 6196 -1153 6214 -1125
rect 6244 -1153 6263 -1125
rect 6468 -1153 6486 -1125
rect 6516 -1153 6534 -1125
rect 6776 -1153 6794 -1125
rect 6824 -1153 6843 -1125
rect 165 -1322 192 -1298
rect 259 -1320 291 -1298
rect 259 -1322 261 -1320
rect 289 -1322 291 -1320
rect 358 -1322 385 -1298
rect 165 -1336 259 -1322
rect 291 -1336 385 -1322
rect 745 -1322 772 -1298
rect 839 -1320 871 -1298
rect 839 -1322 841 -1320
rect 869 -1322 871 -1320
rect 938 -1322 965 -1298
rect 745 -1336 839 -1322
rect 871 -1336 965 -1322
rect 1325 -1322 1352 -1298
rect 1419 -1320 1451 -1298
rect 1419 -1322 1421 -1320
rect 1449 -1322 1451 -1320
rect 1518 -1322 1545 -1298
rect 1325 -1336 1419 -1322
rect 1451 -1336 1545 -1322
rect 1905 -1322 1932 -1298
rect 1999 -1320 2031 -1298
rect 1999 -1322 2001 -1320
rect 2029 -1322 2031 -1320
rect 2098 -1322 2125 -1298
rect 1905 -1336 1999 -1322
rect 2031 -1336 2125 -1322
rect 2485 -1322 2512 -1298
rect 2579 -1320 2611 -1298
rect 2579 -1322 2581 -1320
rect 2609 -1322 2611 -1320
rect 2678 -1322 2705 -1298
rect 2485 -1336 2579 -1322
rect 2611 -1336 2705 -1322
rect 3065 -1322 3092 -1298
rect 3159 -1320 3191 -1298
rect 3159 -1322 3161 -1320
rect 3189 -1322 3191 -1320
rect 3258 -1322 3285 -1298
rect 3065 -1336 3159 -1322
rect 3191 -1336 3285 -1322
rect 3645 -1322 3672 -1298
rect 3739 -1320 3771 -1298
rect 3739 -1322 3741 -1320
rect 3769 -1322 3771 -1320
rect 3838 -1322 3865 -1298
rect 3645 -1336 3739 -1322
rect 3771 -1336 3865 -1322
rect 4225 -1322 4252 -1298
rect 4319 -1320 4351 -1298
rect 4319 -1322 4321 -1320
rect 4349 -1322 4351 -1320
rect 4418 -1322 4445 -1298
rect 4654 -1299 4682 -1257
rect 4712 -1271 4737 -1257
rect 4836 -1267 4861 -1257
rect 4712 -1299 4768 -1271
rect 4798 -1299 4832 -1271
tri 4846 -1274 4853 -1267 ne
rect 4853 -1299 4861 -1267
rect 4891 -1299 4939 -1257
rect 4969 -1267 4994 -1257
rect 4969 -1299 4977 -1267
rect 5093 -1271 5118 -1257
rect 4998 -1299 5032 -1271
rect 5062 -1299 5118 -1271
rect 5148 -1299 5176 -1257
rect 5234 -1299 5262 -1257
rect 5292 -1271 5317 -1257
rect 5416 -1267 5441 -1257
rect 5292 -1299 5348 -1271
rect 5378 -1299 5412 -1271
tri 5426 -1274 5433 -1267 ne
rect 5433 -1299 5441 -1267
rect 5471 -1299 5519 -1257
rect 5549 -1267 5574 -1257
rect 5549 -1299 5557 -1267
rect 5673 -1271 5698 -1257
rect 5578 -1299 5612 -1271
rect 5642 -1299 5698 -1271
rect 5728 -1299 5756 -1257
rect 5814 -1299 5842 -1257
rect 5872 -1271 5897 -1257
rect 5996 -1267 6021 -1257
rect 5872 -1299 5928 -1271
rect 5958 -1299 5992 -1271
tri 6006 -1274 6013 -1267 ne
rect 6013 -1299 6021 -1267
rect 6051 -1299 6099 -1257
rect 6129 -1267 6154 -1257
rect 6129 -1299 6137 -1267
rect 6253 -1271 6278 -1257
rect 6158 -1299 6192 -1271
rect 6222 -1299 6278 -1271
rect 6308 -1299 6336 -1257
rect 6394 -1299 6422 -1257
rect 6452 -1271 6477 -1257
rect 6576 -1267 6601 -1257
rect 6452 -1299 6508 -1271
rect 6538 -1299 6572 -1271
tri 6586 -1274 6593 -1267 ne
rect 6593 -1299 6601 -1267
rect 6631 -1299 6679 -1257
rect 6709 -1267 6734 -1257
rect 6709 -1299 6717 -1267
rect 6833 -1271 6858 -1257
rect 6738 -1299 6772 -1271
rect 6802 -1299 6858 -1271
rect 6888 -1299 6916 -1257
rect 4225 -1336 4319 -1322
rect 4351 -1336 4445 -1322
rect 4805 -1323 4832 -1299
rect 4899 -1321 4931 -1299
rect 4899 -1323 4901 -1321
rect 4929 -1323 4931 -1321
rect 4998 -1323 5025 -1299
rect 4805 -1337 4899 -1323
rect 4931 -1337 5025 -1323
rect 5385 -1323 5412 -1299
rect 5479 -1321 5511 -1299
rect 5479 -1323 5481 -1321
rect 5509 -1323 5511 -1321
rect 5578 -1323 5605 -1299
rect 5385 -1337 5479 -1323
rect 5511 -1337 5605 -1323
rect 5965 -1323 5992 -1299
rect 6059 -1321 6091 -1299
rect 6059 -1323 6061 -1321
rect 6089 -1323 6091 -1321
rect 6158 -1323 6185 -1299
rect 5965 -1337 6059 -1323
rect 6091 -1337 6185 -1323
rect 6545 -1323 6572 -1299
rect 6639 -1321 6671 -1299
rect 6639 -1323 6641 -1321
rect 6669 -1323 6671 -1321
rect 6738 -1323 6765 -1299
rect 6545 -1337 6639 -1323
rect 6671 -1337 6765 -1323
rect 88 -1422 106 -1394
rect 136 -1422 154 -1394
rect 396 -1422 414 -1394
rect 444 -1422 463 -1394
rect 668 -1422 686 -1394
rect 716 -1422 734 -1394
rect 976 -1422 994 -1394
rect 1024 -1422 1043 -1394
rect 1248 -1422 1266 -1394
rect 1296 -1422 1314 -1394
rect 1556 -1422 1574 -1394
rect 1604 -1422 1623 -1394
rect 1828 -1422 1846 -1394
rect 1876 -1422 1894 -1394
rect 2136 -1422 2154 -1394
rect 2184 -1422 2203 -1394
rect 2408 -1422 2426 -1394
rect 2456 -1422 2474 -1394
rect 2716 -1422 2734 -1394
rect 2764 -1422 2783 -1394
rect 2988 -1422 3006 -1394
rect 3036 -1422 3054 -1394
rect 3296 -1422 3314 -1394
rect 3344 -1422 3363 -1394
rect 3568 -1422 3586 -1394
rect 3616 -1422 3634 -1394
rect 3876 -1422 3894 -1394
rect 3924 -1422 3943 -1394
rect 4148 -1422 4166 -1394
rect 4196 -1422 4214 -1394
rect 4456 -1422 4474 -1394
rect 4504 -1422 4523 -1394
rect 4728 -1423 4746 -1395
rect 4776 -1423 4794 -1395
rect 5036 -1423 5054 -1395
rect 5084 -1423 5103 -1395
rect 5308 -1423 5326 -1395
rect 5356 -1423 5374 -1395
rect 14 -1568 42 -1526
rect 72 -1540 97 -1526
rect 196 -1536 221 -1526
rect 72 -1568 128 -1540
rect 158 -1568 192 -1540
tri 206 -1543 213 -1536 ne
rect 213 -1568 221 -1536
rect 251 -1568 299 -1526
rect 329 -1536 354 -1526
rect 329 -1568 337 -1536
rect 453 -1540 478 -1526
rect 358 -1568 392 -1540
rect 422 -1568 478 -1540
rect 508 -1568 536 -1526
rect 594 -1568 622 -1526
rect 652 -1540 677 -1526
rect 776 -1536 801 -1526
rect 652 -1568 708 -1540
rect 738 -1568 772 -1540
tri 786 -1543 793 -1536 ne
rect 793 -1568 801 -1536
rect 831 -1568 879 -1526
rect 909 -1536 934 -1526
rect 909 -1568 917 -1536
rect 1033 -1540 1058 -1526
rect 938 -1568 972 -1540
rect 1002 -1568 1058 -1540
rect 1088 -1568 1116 -1526
rect 1174 -1568 1202 -1526
rect 1232 -1540 1257 -1526
rect 1356 -1536 1381 -1526
rect 1232 -1568 1288 -1540
rect 1318 -1568 1352 -1540
tri 1366 -1543 1373 -1536 ne
rect 1373 -1568 1381 -1536
rect 1411 -1568 1459 -1526
rect 1489 -1536 1514 -1526
rect 1489 -1568 1497 -1536
rect 1613 -1540 1638 -1526
rect 1518 -1568 1552 -1540
rect 1582 -1568 1638 -1540
rect 1668 -1568 1696 -1526
rect 1754 -1568 1782 -1526
rect 1812 -1540 1837 -1526
rect 1936 -1536 1961 -1526
rect 1812 -1568 1868 -1540
rect 1898 -1568 1932 -1540
tri 1946 -1543 1953 -1536 ne
rect 1953 -1568 1961 -1536
rect 1991 -1568 2039 -1526
rect 2069 -1536 2094 -1526
rect 2069 -1568 2077 -1536
rect 2193 -1540 2218 -1526
rect 2098 -1568 2132 -1540
rect 2162 -1568 2218 -1540
rect 2248 -1568 2276 -1526
rect 2334 -1568 2362 -1526
rect 2392 -1540 2417 -1526
rect 2516 -1536 2541 -1526
rect 2392 -1568 2448 -1540
rect 2478 -1568 2512 -1540
tri 2526 -1543 2533 -1536 ne
rect 2533 -1568 2541 -1536
rect 2571 -1568 2619 -1526
rect 2649 -1536 2674 -1526
rect 2649 -1568 2657 -1536
rect 2773 -1540 2798 -1526
rect 2678 -1568 2712 -1540
rect 2742 -1568 2798 -1540
rect 2828 -1568 2856 -1526
rect 2914 -1568 2942 -1526
rect 2972 -1540 2997 -1526
rect 3096 -1536 3121 -1526
rect 2972 -1568 3028 -1540
rect 3058 -1568 3092 -1540
tri 3106 -1543 3113 -1536 ne
rect 3113 -1568 3121 -1536
rect 3151 -1568 3199 -1526
rect 3229 -1536 3254 -1526
rect 3229 -1568 3237 -1536
rect 3353 -1540 3378 -1526
rect 3258 -1568 3292 -1540
rect 3322 -1568 3378 -1540
rect 3408 -1568 3436 -1526
rect 3494 -1568 3522 -1526
rect 3552 -1540 3577 -1526
rect 3676 -1536 3701 -1526
rect 3552 -1568 3608 -1540
rect 3638 -1568 3672 -1540
tri 3686 -1543 3693 -1536 ne
rect 3693 -1568 3701 -1536
rect 3731 -1568 3779 -1526
rect 3809 -1536 3834 -1526
rect 3809 -1568 3817 -1536
rect 3933 -1540 3958 -1526
rect 3838 -1568 3872 -1540
rect 3902 -1568 3958 -1540
rect 3988 -1568 4016 -1526
rect 4074 -1568 4102 -1526
rect 4132 -1540 4157 -1526
rect 4256 -1536 4281 -1526
rect 4132 -1568 4188 -1540
rect 4218 -1568 4252 -1540
tri 4266 -1543 4273 -1536 ne
rect 4273 -1568 4281 -1536
rect 4311 -1568 4359 -1526
rect 4389 -1536 4414 -1526
rect 4389 -1568 4397 -1536
rect 4513 -1540 4538 -1526
rect 4418 -1568 4452 -1540
rect 4482 -1568 4538 -1540
rect 4568 -1568 4596 -1526
rect 5616 -1423 5634 -1395
rect 5664 -1423 5683 -1395
rect 5888 -1423 5906 -1395
rect 5936 -1423 5954 -1395
rect 6196 -1423 6214 -1395
rect 6244 -1423 6263 -1395
rect 6468 -1423 6486 -1395
rect 6516 -1423 6534 -1395
rect 6776 -1423 6794 -1395
rect 6824 -1423 6843 -1395
rect 165 -1592 192 -1568
rect 259 -1590 291 -1568
rect 259 -1592 261 -1590
rect 289 -1592 291 -1590
rect 358 -1592 385 -1568
rect 165 -1606 259 -1592
rect 291 -1606 385 -1592
rect 745 -1592 772 -1568
rect 839 -1590 871 -1568
rect 839 -1592 841 -1590
rect 869 -1592 871 -1590
rect 938 -1592 965 -1568
rect 745 -1606 839 -1592
rect 871 -1606 965 -1592
rect 1325 -1592 1352 -1568
rect 1419 -1590 1451 -1568
rect 1419 -1592 1421 -1590
rect 1449 -1592 1451 -1590
rect 1518 -1592 1545 -1568
rect 1325 -1606 1419 -1592
rect 1451 -1606 1545 -1592
rect 1905 -1592 1932 -1568
rect 1999 -1590 2031 -1568
rect 1999 -1592 2001 -1590
rect 2029 -1592 2031 -1590
rect 2098 -1592 2125 -1568
rect 1905 -1606 1999 -1592
rect 2031 -1606 2125 -1592
rect 2485 -1592 2512 -1568
rect 2579 -1590 2611 -1568
rect 2579 -1592 2581 -1590
rect 2609 -1592 2611 -1590
rect 2678 -1592 2705 -1568
rect 2485 -1606 2579 -1592
rect 2611 -1606 2705 -1592
rect 3065 -1592 3092 -1568
rect 3159 -1590 3191 -1568
rect 3159 -1592 3161 -1590
rect 3189 -1592 3191 -1590
rect 3258 -1592 3285 -1568
rect 3065 -1606 3159 -1592
rect 3191 -1606 3285 -1592
rect 3645 -1592 3672 -1568
rect 3739 -1590 3771 -1568
rect 3739 -1592 3741 -1590
rect 3769 -1592 3771 -1590
rect 3838 -1592 3865 -1568
rect 3645 -1606 3739 -1592
rect 3771 -1606 3865 -1592
rect 4225 -1592 4252 -1568
rect 4319 -1590 4351 -1568
rect 4319 -1592 4321 -1590
rect 4349 -1592 4351 -1590
rect 4418 -1592 4445 -1568
rect 4654 -1569 4682 -1527
rect 4712 -1541 4737 -1527
rect 4836 -1537 4861 -1527
rect 4712 -1569 4768 -1541
rect 4798 -1569 4832 -1541
tri 4846 -1544 4853 -1537 ne
rect 4853 -1569 4861 -1537
rect 4891 -1569 4939 -1527
rect 4969 -1537 4994 -1527
rect 4969 -1569 4977 -1537
rect 5093 -1541 5118 -1527
rect 4998 -1569 5032 -1541
rect 5062 -1569 5118 -1541
rect 5148 -1569 5176 -1527
rect 5234 -1569 5262 -1527
rect 5292 -1541 5317 -1527
rect 5416 -1537 5441 -1527
rect 5292 -1569 5348 -1541
rect 5378 -1569 5412 -1541
tri 5426 -1544 5433 -1537 ne
rect 5433 -1569 5441 -1537
rect 5471 -1569 5519 -1527
rect 5549 -1537 5574 -1527
rect 5549 -1569 5557 -1537
rect 5673 -1541 5698 -1527
rect 5578 -1569 5612 -1541
rect 5642 -1569 5698 -1541
rect 5728 -1569 5756 -1527
rect 5814 -1569 5842 -1527
rect 5872 -1541 5897 -1527
rect 5996 -1537 6021 -1527
rect 5872 -1569 5928 -1541
rect 5958 -1569 5992 -1541
tri 6006 -1544 6013 -1537 ne
rect 6013 -1569 6021 -1537
rect 6051 -1569 6099 -1527
rect 6129 -1537 6154 -1527
rect 6129 -1569 6137 -1537
rect 6253 -1541 6278 -1527
rect 6158 -1569 6192 -1541
rect 6222 -1569 6278 -1541
rect 6308 -1569 6336 -1527
rect 6394 -1569 6422 -1527
rect 6452 -1541 6477 -1527
rect 6576 -1537 6601 -1527
rect 6452 -1569 6508 -1541
rect 6538 -1569 6572 -1541
tri 6586 -1544 6593 -1537 ne
rect 6593 -1569 6601 -1537
rect 6631 -1569 6679 -1527
rect 6709 -1537 6734 -1527
rect 6709 -1569 6717 -1537
rect 6833 -1541 6858 -1527
rect 6738 -1569 6772 -1541
rect 6802 -1569 6858 -1541
rect 6888 -1569 6916 -1527
rect 4225 -1606 4319 -1592
rect 4351 -1606 4445 -1592
rect 4805 -1593 4832 -1569
rect 4899 -1591 4931 -1569
rect 4899 -1593 4901 -1591
rect 4929 -1593 4931 -1591
rect 4998 -1593 5025 -1569
rect 4805 -1607 4899 -1593
rect 4931 -1607 5025 -1593
rect 5385 -1593 5412 -1569
rect 5479 -1591 5511 -1569
rect 5479 -1593 5481 -1591
rect 5509 -1593 5511 -1591
rect 5578 -1593 5605 -1569
rect 5385 -1607 5479 -1593
rect 5511 -1607 5605 -1593
rect 5965 -1593 5992 -1569
rect 6059 -1591 6091 -1569
rect 6059 -1593 6061 -1591
rect 6089 -1593 6091 -1591
rect 6158 -1593 6185 -1569
rect 5965 -1607 6059 -1593
rect 6091 -1607 6185 -1593
rect 6545 -1593 6572 -1569
rect 6639 -1591 6671 -1569
rect 6639 -1593 6641 -1591
rect 6669 -1593 6671 -1591
rect 6738 -1593 6765 -1569
rect 6545 -1607 6639 -1593
rect 6671 -1607 6765 -1593
rect 88 -1692 106 -1664
rect 136 -1692 154 -1664
rect 396 -1692 414 -1664
rect 444 -1692 463 -1664
rect 668 -1692 686 -1664
rect 716 -1692 734 -1664
rect 976 -1692 994 -1664
rect 1024 -1692 1043 -1664
rect 1248 -1692 1266 -1664
rect 1296 -1692 1314 -1664
rect 1556 -1692 1574 -1664
rect 1604 -1692 1623 -1664
rect 1828 -1692 1846 -1664
rect 1876 -1692 1894 -1664
rect 2136 -1692 2154 -1664
rect 2184 -1692 2203 -1664
rect 2408 -1692 2426 -1664
rect 2456 -1692 2474 -1664
rect 2716 -1692 2734 -1664
rect 2764 -1692 2783 -1664
rect 2988 -1692 3006 -1664
rect 3036 -1692 3054 -1664
rect 3296 -1692 3314 -1664
rect 3344 -1692 3363 -1664
rect 3568 -1692 3586 -1664
rect 3616 -1692 3634 -1664
rect 3876 -1692 3894 -1664
rect 3924 -1692 3943 -1664
rect 4148 -1692 4166 -1664
rect 4196 -1692 4214 -1664
rect 4456 -1692 4474 -1664
rect 4504 -1692 4523 -1664
rect 4728 -1693 4746 -1665
rect 4776 -1693 4794 -1665
rect 5036 -1693 5054 -1665
rect 5084 -1693 5103 -1665
rect 5308 -1693 5326 -1665
rect 5356 -1693 5374 -1665
rect 14 -1838 42 -1796
rect 72 -1810 97 -1796
rect 196 -1806 221 -1796
rect 72 -1838 128 -1810
rect 158 -1838 192 -1810
tri 206 -1813 213 -1806 ne
rect 213 -1838 221 -1806
rect 251 -1838 299 -1796
rect 329 -1806 354 -1796
rect 329 -1838 337 -1806
rect 453 -1810 478 -1796
rect 358 -1838 392 -1810
rect 422 -1838 478 -1810
rect 508 -1838 536 -1796
rect 594 -1838 622 -1796
rect 652 -1810 677 -1796
rect 776 -1806 801 -1796
rect 652 -1838 708 -1810
rect 738 -1838 772 -1810
tri 786 -1813 793 -1806 ne
rect 793 -1838 801 -1806
rect 831 -1838 879 -1796
rect 909 -1806 934 -1796
rect 909 -1838 917 -1806
rect 1033 -1810 1058 -1796
rect 938 -1838 972 -1810
rect 1002 -1838 1058 -1810
rect 1088 -1838 1116 -1796
rect 1174 -1838 1202 -1796
rect 1232 -1810 1257 -1796
rect 1356 -1806 1381 -1796
rect 1232 -1838 1288 -1810
rect 1318 -1838 1352 -1810
tri 1366 -1813 1373 -1806 ne
rect 1373 -1838 1381 -1806
rect 1411 -1838 1459 -1796
rect 1489 -1806 1514 -1796
rect 1489 -1838 1497 -1806
rect 1613 -1810 1638 -1796
rect 1518 -1838 1552 -1810
rect 1582 -1838 1638 -1810
rect 1668 -1838 1696 -1796
rect 1754 -1838 1782 -1796
rect 1812 -1810 1837 -1796
rect 1936 -1806 1961 -1796
rect 1812 -1838 1868 -1810
rect 1898 -1838 1932 -1810
tri 1946 -1813 1953 -1806 ne
rect 1953 -1838 1961 -1806
rect 1991 -1838 2039 -1796
rect 2069 -1806 2094 -1796
rect 2069 -1838 2077 -1806
rect 2193 -1810 2218 -1796
rect 2098 -1838 2132 -1810
rect 2162 -1838 2218 -1810
rect 2248 -1838 2276 -1796
rect 2334 -1838 2362 -1796
rect 2392 -1810 2417 -1796
rect 2516 -1806 2541 -1796
rect 2392 -1838 2448 -1810
rect 2478 -1838 2512 -1810
tri 2526 -1813 2533 -1806 ne
rect 2533 -1838 2541 -1806
rect 2571 -1838 2619 -1796
rect 2649 -1806 2674 -1796
rect 2649 -1838 2657 -1806
rect 2773 -1810 2798 -1796
rect 2678 -1838 2712 -1810
rect 2742 -1838 2798 -1810
rect 2828 -1838 2856 -1796
rect 2914 -1838 2942 -1796
rect 2972 -1810 2997 -1796
rect 3096 -1806 3121 -1796
rect 2972 -1838 3028 -1810
rect 3058 -1838 3092 -1810
tri 3106 -1813 3113 -1806 ne
rect 3113 -1838 3121 -1806
rect 3151 -1838 3199 -1796
rect 3229 -1806 3254 -1796
rect 3229 -1838 3237 -1806
rect 3353 -1810 3378 -1796
rect 3258 -1838 3292 -1810
rect 3322 -1838 3378 -1810
rect 3408 -1838 3436 -1796
rect 3494 -1838 3522 -1796
rect 3552 -1810 3577 -1796
rect 3676 -1806 3701 -1796
rect 3552 -1838 3608 -1810
rect 3638 -1838 3672 -1810
tri 3686 -1813 3693 -1806 ne
rect 3693 -1838 3701 -1806
rect 3731 -1838 3779 -1796
rect 3809 -1806 3834 -1796
rect 3809 -1838 3817 -1806
rect 3933 -1810 3958 -1796
rect 3838 -1838 3872 -1810
rect 3902 -1838 3958 -1810
rect 3988 -1838 4016 -1796
rect 4074 -1838 4102 -1796
rect 4132 -1810 4157 -1796
rect 4256 -1806 4281 -1796
rect 4132 -1838 4188 -1810
rect 4218 -1838 4252 -1810
tri 4266 -1813 4273 -1806 ne
rect 4273 -1838 4281 -1806
rect 4311 -1838 4359 -1796
rect 4389 -1806 4414 -1796
rect 4389 -1838 4397 -1806
rect 4513 -1810 4538 -1796
rect 4418 -1838 4452 -1810
rect 4482 -1838 4538 -1810
rect 4568 -1838 4596 -1796
rect 5616 -1693 5634 -1665
rect 5664 -1693 5683 -1665
rect 5888 -1693 5906 -1665
rect 5936 -1693 5954 -1665
rect 6196 -1693 6214 -1665
rect 6244 -1693 6263 -1665
rect 6468 -1693 6486 -1665
rect 6516 -1693 6534 -1665
rect 6776 -1693 6794 -1665
rect 6824 -1693 6843 -1665
rect 165 -1862 192 -1838
rect 259 -1860 291 -1838
rect 259 -1862 261 -1860
rect 289 -1862 291 -1860
rect 358 -1862 385 -1838
rect 165 -1876 259 -1862
rect 291 -1876 385 -1862
rect 745 -1862 772 -1838
rect 839 -1860 871 -1838
rect 839 -1862 841 -1860
rect 869 -1862 871 -1860
rect 938 -1862 965 -1838
rect 745 -1876 839 -1862
rect 871 -1876 965 -1862
rect 1325 -1862 1352 -1838
rect 1419 -1860 1451 -1838
rect 1419 -1862 1421 -1860
rect 1449 -1862 1451 -1860
rect 1518 -1862 1545 -1838
rect 1325 -1876 1419 -1862
rect 1451 -1876 1545 -1862
rect 1905 -1862 1932 -1838
rect 1999 -1860 2031 -1838
rect 1999 -1862 2001 -1860
rect 2029 -1862 2031 -1860
rect 2098 -1862 2125 -1838
rect 1905 -1876 1999 -1862
rect 2031 -1876 2125 -1862
rect 2485 -1862 2512 -1838
rect 2579 -1860 2611 -1838
rect 2579 -1862 2581 -1860
rect 2609 -1862 2611 -1860
rect 2678 -1862 2705 -1838
rect 2485 -1876 2579 -1862
rect 2611 -1876 2705 -1862
rect 3065 -1862 3092 -1838
rect 3159 -1860 3191 -1838
rect 3159 -1862 3161 -1860
rect 3189 -1862 3191 -1860
rect 3258 -1862 3285 -1838
rect 3065 -1876 3159 -1862
rect 3191 -1876 3285 -1862
rect 3645 -1862 3672 -1838
rect 3739 -1860 3771 -1838
rect 3739 -1862 3741 -1860
rect 3769 -1862 3771 -1860
rect 3838 -1862 3865 -1838
rect 3645 -1876 3739 -1862
rect 3771 -1876 3865 -1862
rect 4225 -1862 4252 -1838
rect 4319 -1860 4351 -1838
rect 4319 -1862 4321 -1860
rect 4349 -1862 4351 -1860
rect 4418 -1862 4445 -1838
rect 4654 -1839 4682 -1797
rect 4712 -1811 4737 -1797
rect 4836 -1807 4861 -1797
rect 4712 -1839 4768 -1811
rect 4798 -1839 4832 -1811
tri 4846 -1814 4853 -1807 ne
rect 4853 -1839 4861 -1807
rect 4891 -1839 4939 -1797
rect 4969 -1807 4994 -1797
rect 4969 -1839 4977 -1807
rect 5093 -1811 5118 -1797
rect 4998 -1839 5032 -1811
rect 5062 -1839 5118 -1811
rect 5148 -1839 5176 -1797
rect 5234 -1839 5262 -1797
rect 5292 -1811 5317 -1797
rect 5416 -1807 5441 -1797
rect 5292 -1839 5348 -1811
rect 5378 -1839 5412 -1811
tri 5426 -1814 5433 -1807 ne
rect 5433 -1839 5441 -1807
rect 5471 -1839 5519 -1797
rect 5549 -1807 5574 -1797
rect 5549 -1839 5557 -1807
rect 5673 -1811 5698 -1797
rect 5578 -1839 5612 -1811
rect 5642 -1839 5698 -1811
rect 5728 -1839 5756 -1797
rect 5814 -1839 5842 -1797
rect 5872 -1811 5897 -1797
rect 5996 -1807 6021 -1797
rect 5872 -1839 5928 -1811
rect 5958 -1839 5992 -1811
tri 6006 -1814 6013 -1807 ne
rect 6013 -1839 6021 -1807
rect 6051 -1839 6099 -1797
rect 6129 -1807 6154 -1797
rect 6129 -1839 6137 -1807
rect 6253 -1811 6278 -1797
rect 6158 -1839 6192 -1811
rect 6222 -1839 6278 -1811
rect 6308 -1839 6336 -1797
rect 6394 -1839 6422 -1797
rect 6452 -1811 6477 -1797
rect 6576 -1807 6601 -1797
rect 6452 -1839 6508 -1811
rect 6538 -1839 6572 -1811
tri 6586 -1814 6593 -1807 ne
rect 6593 -1839 6601 -1807
rect 6631 -1839 6679 -1797
rect 6709 -1807 6734 -1797
rect 6709 -1839 6717 -1807
rect 6833 -1811 6858 -1797
rect 6738 -1839 6772 -1811
rect 6802 -1839 6858 -1811
rect 6888 -1839 6916 -1797
rect 4225 -1876 4319 -1862
rect 4351 -1876 4445 -1862
rect 4805 -1863 4832 -1839
rect 4899 -1861 4931 -1839
rect 4899 -1863 4901 -1861
rect 4929 -1863 4931 -1861
rect 4998 -1863 5025 -1839
rect 4805 -1877 4899 -1863
rect 4931 -1877 5025 -1863
rect 5385 -1863 5412 -1839
rect 5479 -1861 5511 -1839
rect 5479 -1863 5481 -1861
rect 5509 -1863 5511 -1861
rect 5578 -1863 5605 -1839
rect 5385 -1877 5479 -1863
rect 5511 -1877 5605 -1863
rect 5965 -1863 5992 -1839
rect 6059 -1861 6091 -1839
rect 6059 -1863 6061 -1861
rect 6089 -1863 6091 -1861
rect 6158 -1863 6185 -1839
rect 5965 -1877 6059 -1863
rect 6091 -1877 6185 -1863
rect 6545 -1863 6572 -1839
rect 6639 -1861 6671 -1839
rect 6639 -1863 6641 -1861
rect 6669 -1863 6671 -1861
rect 6738 -1863 6765 -1839
rect 6545 -1877 6639 -1863
rect 6671 -1877 6765 -1863
rect 88 -1962 106 -1934
rect 136 -1962 154 -1934
rect 396 -1962 414 -1934
rect 444 -1962 463 -1934
rect 668 -1962 686 -1934
rect 716 -1962 734 -1934
rect 976 -1962 994 -1934
rect 1024 -1962 1043 -1934
rect 1248 -1962 1266 -1934
rect 1296 -1962 1314 -1934
rect 1556 -1962 1574 -1934
rect 1604 -1962 1623 -1934
rect 1828 -1962 1846 -1934
rect 1876 -1962 1894 -1934
rect 2136 -1962 2154 -1934
rect 2184 -1962 2203 -1934
rect 2408 -1962 2426 -1934
rect 2456 -1962 2474 -1934
rect 2716 -1962 2734 -1934
rect 2764 -1962 2783 -1934
rect 2988 -1962 3006 -1934
rect 3036 -1962 3054 -1934
rect 3296 -1962 3314 -1934
rect 3344 -1962 3363 -1934
rect 3568 -1962 3586 -1934
rect 3616 -1962 3634 -1934
rect 3876 -1962 3894 -1934
rect 3924 -1962 3943 -1934
rect 4148 -1962 4166 -1934
rect 4196 -1962 4214 -1934
rect 4456 -1962 4474 -1934
rect 4504 -1962 4523 -1934
rect 4728 -1963 4746 -1935
rect 4776 -1963 4794 -1935
rect 5036 -1963 5054 -1935
rect 5084 -1963 5103 -1935
rect 5308 -1963 5326 -1935
rect 5356 -1963 5374 -1935
rect 14 -2108 42 -2066
rect 72 -2080 97 -2066
rect 196 -2076 221 -2066
rect 72 -2108 128 -2080
rect 158 -2108 192 -2080
tri 206 -2083 213 -2076 ne
rect 213 -2108 221 -2076
rect 251 -2108 299 -2066
rect 329 -2076 354 -2066
rect 329 -2108 337 -2076
rect 453 -2080 478 -2066
rect 358 -2108 392 -2080
rect 422 -2108 478 -2080
rect 508 -2108 536 -2066
rect 594 -2108 622 -2066
rect 652 -2080 677 -2066
rect 776 -2076 801 -2066
rect 652 -2108 708 -2080
rect 738 -2108 772 -2080
tri 786 -2083 793 -2076 ne
rect 793 -2108 801 -2076
rect 831 -2108 879 -2066
rect 909 -2076 934 -2066
rect 909 -2108 917 -2076
rect 1033 -2080 1058 -2066
rect 938 -2108 972 -2080
rect 1002 -2108 1058 -2080
rect 1088 -2108 1116 -2066
rect 1174 -2108 1202 -2066
rect 1232 -2080 1257 -2066
rect 1356 -2076 1381 -2066
rect 1232 -2108 1288 -2080
rect 1318 -2108 1352 -2080
tri 1366 -2083 1373 -2076 ne
rect 1373 -2108 1381 -2076
rect 1411 -2108 1459 -2066
rect 1489 -2076 1514 -2066
rect 1489 -2108 1497 -2076
rect 1613 -2080 1638 -2066
rect 1518 -2108 1552 -2080
rect 1582 -2108 1638 -2080
rect 1668 -2108 1696 -2066
rect 1754 -2108 1782 -2066
rect 1812 -2080 1837 -2066
rect 1936 -2076 1961 -2066
rect 1812 -2108 1868 -2080
rect 1898 -2108 1932 -2080
tri 1946 -2083 1953 -2076 ne
rect 1953 -2108 1961 -2076
rect 1991 -2108 2039 -2066
rect 2069 -2076 2094 -2066
rect 2069 -2108 2077 -2076
rect 2193 -2080 2218 -2066
rect 2098 -2108 2132 -2080
rect 2162 -2108 2218 -2080
rect 2248 -2108 2276 -2066
rect 2334 -2108 2362 -2066
rect 2392 -2080 2417 -2066
rect 2516 -2076 2541 -2066
rect 2392 -2108 2448 -2080
rect 2478 -2108 2512 -2080
tri 2526 -2083 2533 -2076 ne
rect 2533 -2108 2541 -2076
rect 2571 -2108 2619 -2066
rect 2649 -2076 2674 -2066
rect 2649 -2108 2657 -2076
rect 2773 -2080 2798 -2066
rect 2678 -2108 2712 -2080
rect 2742 -2108 2798 -2080
rect 2828 -2108 2856 -2066
rect 2914 -2108 2942 -2066
rect 2972 -2080 2997 -2066
rect 3096 -2076 3121 -2066
rect 2972 -2108 3028 -2080
rect 3058 -2108 3092 -2080
tri 3106 -2083 3113 -2076 ne
rect 3113 -2108 3121 -2076
rect 3151 -2108 3199 -2066
rect 3229 -2076 3254 -2066
rect 3229 -2108 3237 -2076
rect 3353 -2080 3378 -2066
rect 3258 -2108 3292 -2080
rect 3322 -2108 3378 -2080
rect 3408 -2108 3436 -2066
rect 3494 -2108 3522 -2066
rect 3552 -2080 3577 -2066
rect 3676 -2076 3701 -2066
rect 3552 -2108 3608 -2080
rect 3638 -2108 3672 -2080
tri 3686 -2083 3693 -2076 ne
rect 3693 -2108 3701 -2076
rect 3731 -2108 3779 -2066
rect 3809 -2076 3834 -2066
rect 3809 -2108 3817 -2076
rect 3933 -2080 3958 -2066
rect 3838 -2108 3872 -2080
rect 3902 -2108 3958 -2080
rect 3988 -2108 4016 -2066
rect 4074 -2108 4102 -2066
rect 4132 -2080 4157 -2066
rect 4256 -2076 4281 -2066
rect 4132 -2108 4188 -2080
rect 4218 -2108 4252 -2080
tri 4266 -2083 4273 -2076 ne
rect 4273 -2108 4281 -2076
rect 4311 -2108 4359 -2066
rect 4389 -2076 4414 -2066
rect 4389 -2108 4397 -2076
rect 4513 -2080 4538 -2066
rect 4418 -2108 4452 -2080
rect 4482 -2108 4538 -2080
rect 4568 -2108 4596 -2066
rect 5616 -1963 5634 -1935
rect 5664 -1963 5683 -1935
rect 5888 -1963 5906 -1935
rect 5936 -1963 5954 -1935
rect 6196 -1963 6214 -1935
rect 6244 -1963 6263 -1935
rect 6468 -1963 6486 -1935
rect 6516 -1963 6534 -1935
rect 6776 -1963 6794 -1935
rect 6824 -1963 6843 -1935
rect 165 -2132 192 -2108
rect 259 -2130 291 -2108
rect 259 -2132 261 -2130
rect 289 -2132 291 -2130
rect 358 -2132 385 -2108
rect 165 -2146 259 -2132
rect 291 -2146 385 -2132
rect 745 -2132 772 -2108
rect 839 -2130 871 -2108
rect 839 -2132 841 -2130
rect 869 -2132 871 -2130
rect 938 -2132 965 -2108
rect 745 -2146 839 -2132
rect 871 -2146 965 -2132
rect 1325 -2132 1352 -2108
rect 1419 -2130 1451 -2108
rect 1419 -2132 1421 -2130
rect 1449 -2132 1451 -2130
rect 1518 -2132 1545 -2108
rect 1325 -2146 1419 -2132
rect 1451 -2146 1545 -2132
rect 1905 -2132 1932 -2108
rect 1999 -2130 2031 -2108
rect 1999 -2132 2001 -2130
rect 2029 -2132 2031 -2130
rect 2098 -2132 2125 -2108
rect 1905 -2146 1999 -2132
rect 2031 -2146 2125 -2132
rect 2485 -2132 2512 -2108
rect 2579 -2130 2611 -2108
rect 2579 -2132 2581 -2130
rect 2609 -2132 2611 -2130
rect 2678 -2132 2705 -2108
rect 2485 -2146 2579 -2132
rect 2611 -2146 2705 -2132
rect 3065 -2132 3092 -2108
rect 3159 -2130 3191 -2108
rect 3159 -2132 3161 -2130
rect 3189 -2132 3191 -2130
rect 3258 -2132 3285 -2108
rect 3065 -2146 3159 -2132
rect 3191 -2146 3285 -2132
rect 3645 -2132 3672 -2108
rect 3739 -2130 3771 -2108
rect 3739 -2132 3741 -2130
rect 3769 -2132 3771 -2130
rect 3838 -2132 3865 -2108
rect 3645 -2146 3739 -2132
rect 3771 -2146 3865 -2132
rect 4225 -2132 4252 -2108
rect 4319 -2130 4351 -2108
rect 4319 -2132 4321 -2130
rect 4349 -2132 4351 -2130
rect 4418 -2132 4445 -2108
rect 4654 -2109 4682 -2067
rect 4712 -2081 4737 -2067
rect 4836 -2077 4861 -2067
rect 4712 -2109 4768 -2081
rect 4798 -2109 4832 -2081
tri 4846 -2084 4853 -2077 ne
rect 4853 -2109 4861 -2077
rect 4891 -2109 4939 -2067
rect 4969 -2077 4994 -2067
rect 4969 -2109 4977 -2077
rect 5093 -2081 5118 -2067
rect 4998 -2109 5032 -2081
rect 5062 -2109 5118 -2081
rect 5148 -2109 5176 -2067
rect 5234 -2109 5262 -2067
rect 5292 -2081 5317 -2067
rect 5416 -2077 5441 -2067
rect 5292 -2109 5348 -2081
rect 5378 -2109 5412 -2081
tri 5426 -2084 5433 -2077 ne
rect 5433 -2109 5441 -2077
rect 5471 -2109 5519 -2067
rect 5549 -2077 5574 -2067
rect 5549 -2109 5557 -2077
rect 5673 -2081 5698 -2067
rect 5578 -2109 5612 -2081
rect 5642 -2109 5698 -2081
rect 5728 -2109 5756 -2067
rect 5814 -2109 5842 -2067
rect 5872 -2081 5897 -2067
rect 5996 -2077 6021 -2067
rect 5872 -2109 5928 -2081
rect 5958 -2109 5992 -2081
tri 6006 -2084 6013 -2077 ne
rect 6013 -2109 6021 -2077
rect 6051 -2109 6099 -2067
rect 6129 -2077 6154 -2067
rect 6129 -2109 6137 -2077
rect 6253 -2081 6278 -2067
rect 6158 -2109 6192 -2081
rect 6222 -2109 6278 -2081
rect 6308 -2109 6336 -2067
rect 6394 -2109 6422 -2067
rect 6452 -2081 6477 -2067
rect 6576 -2077 6601 -2067
rect 6452 -2109 6508 -2081
rect 6538 -2109 6572 -2081
tri 6586 -2084 6593 -2077 ne
rect 6593 -2109 6601 -2077
rect 6631 -2109 6679 -2067
rect 6709 -2077 6734 -2067
rect 6709 -2109 6717 -2077
rect 6833 -2081 6858 -2067
rect 6738 -2109 6772 -2081
rect 6802 -2109 6858 -2081
rect 6888 -2109 6916 -2067
rect 4225 -2146 4319 -2132
rect 4351 -2146 4445 -2132
rect 4805 -2133 4832 -2109
rect 4899 -2131 4931 -2109
rect 4899 -2133 4901 -2131
rect 4929 -2133 4931 -2131
rect 4998 -2133 5025 -2109
rect 4805 -2147 4899 -2133
rect 4931 -2147 5025 -2133
rect 5385 -2133 5412 -2109
rect 5479 -2131 5511 -2109
rect 5479 -2133 5481 -2131
rect 5509 -2133 5511 -2131
rect 5578 -2133 5605 -2109
rect 5385 -2147 5479 -2133
rect 5511 -2147 5605 -2133
rect 5965 -2133 5992 -2109
rect 6059 -2131 6091 -2109
rect 6059 -2133 6061 -2131
rect 6089 -2133 6091 -2131
rect 6158 -2133 6185 -2109
rect 5965 -2147 6059 -2133
rect 6091 -2147 6185 -2133
rect 6545 -2133 6572 -2109
rect 6639 -2131 6671 -2109
rect 6639 -2133 6641 -2131
rect 6669 -2133 6671 -2131
rect 6738 -2133 6765 -2109
rect 6545 -2147 6639 -2133
rect 6671 -2147 6765 -2133
<< pdiff >>
rect 259 2128 261 2130
rect 289 2128 291 2130
rect 259 2106 291 2128
rect 212 2078 221 2106
rect 251 2078 299 2106
rect 329 2078 338 2106
tri 338 2078 350 2090 sw
rect 839 2128 841 2130
rect 869 2128 871 2130
rect 839 2106 871 2128
rect 792 2078 801 2106
rect 831 2078 879 2106
rect 909 2078 918 2106
tri 918 2078 930 2090 sw
rect 1419 2128 1421 2130
rect 1449 2128 1451 2130
rect 1419 2106 1451 2128
rect 1372 2078 1381 2106
rect 1411 2078 1459 2106
rect 1489 2078 1498 2106
tri 1498 2078 1510 2090 sw
rect 1999 2128 2001 2130
rect 2029 2128 2031 2130
rect 1999 2106 2031 2128
rect 1952 2078 1961 2106
rect 1991 2078 2039 2106
rect 2069 2078 2078 2106
tri 2078 2078 2090 2090 sw
rect 2579 2128 2581 2130
rect 2609 2128 2611 2130
rect 2579 2106 2611 2128
rect 2532 2078 2541 2106
rect 2571 2078 2619 2106
rect 2649 2078 2658 2106
tri 2658 2078 2670 2090 sw
rect 3159 2128 3161 2130
rect 3189 2128 3191 2130
rect 3159 2106 3191 2128
rect 3112 2078 3121 2106
rect 3151 2078 3199 2106
rect 3229 2078 3238 2106
tri 3238 2078 3250 2090 sw
rect 3739 2128 3741 2130
rect 3769 2128 3771 2130
rect 3739 2106 3771 2128
rect 3692 2078 3701 2106
rect 3731 2078 3779 2106
rect 3809 2078 3818 2106
tri 3818 2078 3830 2090 sw
rect 4319 2128 4321 2130
rect 4349 2128 4351 2130
rect 4319 2106 4351 2128
rect 4272 2078 4281 2106
rect 4311 2078 4359 2106
rect 4389 2078 4398 2106
tri 4398 2078 4410 2090 sw
rect 4899 2128 4901 2130
rect 4929 2128 4931 2130
rect 4899 2106 4931 2128
rect 4852 2078 4861 2106
rect 4891 2078 4939 2106
rect 4969 2078 4978 2106
tri 4978 2078 4990 2090 sw
rect 5479 2128 5481 2130
rect 5509 2128 5511 2130
rect 5479 2106 5511 2128
rect 5432 2078 5441 2106
rect 5471 2078 5519 2106
rect 5549 2078 5558 2106
tri 5558 2078 5570 2090 sw
rect 6059 2128 6061 2130
rect 6089 2128 6091 2130
rect 6059 2106 6091 2128
rect 6012 2078 6021 2106
rect 6051 2078 6099 2106
rect 6129 2078 6138 2106
tri 6138 2078 6150 2090 sw
rect 6639 2128 6641 2130
rect 6669 2128 6671 2130
rect 6639 2106 6671 2128
rect 6592 2078 6601 2106
rect 6631 2078 6679 2106
rect 6709 2078 6718 2106
tri 6718 2078 6730 2090 sw
rect 259 1858 261 1860
rect 289 1858 291 1860
rect 259 1836 291 1858
rect 212 1808 221 1836
rect 251 1808 299 1836
rect 329 1808 338 1836
tri 338 1808 350 1820 sw
rect 839 1858 841 1860
rect 869 1858 871 1860
rect 839 1836 871 1858
rect 792 1808 801 1836
rect 831 1808 879 1836
rect 909 1808 918 1836
tri 918 1808 930 1820 sw
rect 1419 1858 1421 1860
rect 1449 1858 1451 1860
rect 1419 1836 1451 1858
rect 1372 1808 1381 1836
rect 1411 1808 1459 1836
rect 1489 1808 1498 1836
tri 1498 1808 1510 1820 sw
rect 1999 1858 2001 1860
rect 2029 1858 2031 1860
rect 1999 1836 2031 1858
rect 1952 1808 1961 1836
rect 1991 1808 2039 1836
rect 2069 1808 2078 1836
tri 2078 1808 2090 1820 sw
rect 2579 1858 2581 1860
rect 2609 1858 2611 1860
rect 2579 1836 2611 1858
rect 2532 1808 2541 1836
rect 2571 1808 2619 1836
rect 2649 1808 2658 1836
tri 2658 1808 2670 1820 sw
rect 3159 1858 3161 1860
rect 3189 1858 3191 1860
rect 3159 1836 3191 1858
rect 3112 1808 3121 1836
rect 3151 1808 3199 1836
rect 3229 1808 3238 1836
tri 3238 1808 3250 1820 sw
rect 3739 1858 3741 1860
rect 3769 1858 3771 1860
rect 3739 1836 3771 1858
rect 3692 1808 3701 1836
rect 3731 1808 3779 1836
rect 3809 1808 3818 1836
tri 3818 1808 3830 1820 sw
rect 4319 1858 4321 1860
rect 4349 1858 4351 1860
rect 4319 1836 4351 1858
rect 4272 1808 4281 1836
rect 4311 1808 4359 1836
rect 4389 1808 4398 1836
tri 4398 1808 4410 1820 sw
rect 4899 1858 4901 1860
rect 4929 1858 4931 1860
rect 4899 1836 4931 1858
rect 4852 1808 4861 1836
rect 4891 1808 4939 1836
rect 4969 1808 4978 1836
tri 4978 1808 4990 1820 sw
rect 5479 1858 5481 1860
rect 5509 1858 5511 1860
rect 5479 1836 5511 1858
rect 5432 1808 5441 1836
rect 5471 1808 5519 1836
rect 5549 1808 5558 1836
tri 5558 1808 5570 1820 sw
rect 6059 1858 6061 1860
rect 6089 1858 6091 1860
rect 6059 1836 6091 1858
rect 6012 1808 6021 1836
rect 6051 1808 6099 1836
rect 6129 1808 6138 1836
tri 6138 1808 6150 1820 sw
rect 6639 1858 6641 1860
rect 6669 1858 6671 1860
rect 6639 1836 6671 1858
rect 6592 1808 6601 1836
rect 6631 1808 6679 1836
rect 6709 1808 6718 1836
tri 6718 1808 6730 1820 sw
rect 259 1588 261 1590
rect 289 1588 291 1590
rect 259 1566 291 1588
rect 212 1538 221 1566
rect 251 1538 299 1566
rect 329 1538 338 1566
tri 338 1538 350 1550 sw
rect 839 1588 841 1590
rect 869 1588 871 1590
rect 839 1566 871 1588
rect 792 1538 801 1566
rect 831 1538 879 1566
rect 909 1538 918 1566
tri 918 1538 930 1550 sw
rect 1419 1588 1421 1590
rect 1449 1588 1451 1590
rect 1419 1566 1451 1588
rect 1372 1538 1381 1566
rect 1411 1538 1459 1566
rect 1489 1538 1498 1566
tri 1498 1538 1510 1550 sw
rect 1999 1588 2001 1590
rect 2029 1588 2031 1590
rect 1999 1566 2031 1588
rect 1952 1538 1961 1566
rect 1991 1538 2039 1566
rect 2069 1538 2078 1566
tri 2078 1538 2090 1550 sw
rect 2579 1588 2581 1590
rect 2609 1588 2611 1590
rect 2579 1566 2611 1588
rect 2532 1538 2541 1566
rect 2571 1538 2619 1566
rect 2649 1538 2658 1566
tri 2658 1538 2670 1550 sw
rect 3159 1588 3161 1590
rect 3189 1588 3191 1590
rect 3159 1566 3191 1588
rect 3112 1538 3121 1566
rect 3151 1538 3199 1566
rect 3229 1538 3238 1566
tri 3238 1538 3250 1550 sw
rect 3739 1588 3741 1590
rect 3769 1588 3771 1590
rect 3739 1566 3771 1588
rect 3692 1538 3701 1566
rect 3731 1538 3779 1566
rect 3809 1538 3818 1566
tri 3818 1538 3830 1550 sw
rect 4319 1588 4321 1590
rect 4349 1588 4351 1590
rect 4319 1566 4351 1588
rect 4272 1538 4281 1566
rect 4311 1538 4359 1566
rect 4389 1538 4398 1566
tri 4398 1538 4410 1550 sw
rect 4899 1588 4901 1590
rect 4929 1588 4931 1590
rect 4899 1566 4931 1588
rect 4852 1538 4861 1566
rect 4891 1538 4939 1566
rect 4969 1538 4978 1566
tri 4978 1538 4990 1550 sw
rect 5479 1588 5481 1590
rect 5509 1588 5511 1590
rect 5479 1566 5511 1588
rect 5432 1538 5441 1566
rect 5471 1538 5519 1566
rect 5549 1538 5558 1566
tri 5558 1538 5570 1550 sw
rect 6059 1588 6061 1590
rect 6089 1588 6091 1590
rect 6059 1566 6091 1588
rect 6012 1538 6021 1566
rect 6051 1538 6099 1566
rect 6129 1538 6138 1566
tri 6138 1538 6150 1550 sw
rect 6639 1588 6641 1590
rect 6669 1588 6671 1590
rect 6639 1566 6671 1588
rect 6592 1538 6601 1566
rect 6631 1538 6679 1566
rect 6709 1538 6718 1566
tri 6718 1538 6730 1550 sw
rect 259 1318 261 1320
rect 289 1318 291 1320
rect 259 1296 291 1318
rect 212 1268 221 1296
rect 251 1268 299 1296
rect 329 1268 338 1296
tri 338 1268 350 1280 sw
rect 839 1318 841 1320
rect 869 1318 871 1320
rect 839 1296 871 1318
rect 792 1268 801 1296
rect 831 1268 879 1296
rect 909 1268 918 1296
tri 918 1268 930 1280 sw
rect 1419 1318 1421 1320
rect 1449 1318 1451 1320
rect 1419 1296 1451 1318
rect 1372 1268 1381 1296
rect 1411 1268 1459 1296
rect 1489 1268 1498 1296
tri 1498 1268 1510 1280 sw
rect 1999 1318 2001 1320
rect 2029 1318 2031 1320
rect 1999 1296 2031 1318
rect 1952 1268 1961 1296
rect 1991 1268 2039 1296
rect 2069 1268 2078 1296
tri 2078 1268 2090 1280 sw
rect 2579 1318 2581 1320
rect 2609 1318 2611 1320
rect 2579 1296 2611 1318
rect 2532 1268 2541 1296
rect 2571 1268 2619 1296
rect 2649 1268 2658 1296
tri 2658 1268 2670 1280 sw
rect 3159 1318 3161 1320
rect 3189 1318 3191 1320
rect 3159 1296 3191 1318
rect 3112 1268 3121 1296
rect 3151 1268 3199 1296
rect 3229 1268 3238 1296
tri 3238 1268 3250 1280 sw
rect 3739 1318 3741 1320
rect 3769 1318 3771 1320
rect 3739 1296 3771 1318
rect 3692 1268 3701 1296
rect 3731 1268 3779 1296
rect 3809 1268 3818 1296
tri 3818 1268 3830 1280 sw
rect 4319 1318 4321 1320
rect 4349 1318 4351 1320
rect 4319 1296 4351 1318
rect 4272 1268 4281 1296
rect 4311 1268 4359 1296
rect 4389 1268 4398 1296
tri 4398 1268 4410 1280 sw
rect 4899 1318 4901 1320
rect 4929 1318 4931 1320
rect 4899 1296 4931 1318
rect 4852 1268 4861 1296
rect 4891 1268 4939 1296
rect 4969 1268 4978 1296
tri 4978 1268 4990 1280 sw
rect 5479 1318 5481 1320
rect 5509 1318 5511 1320
rect 5479 1296 5511 1318
rect 5432 1268 5441 1296
rect 5471 1268 5519 1296
rect 5549 1268 5558 1296
tri 5558 1268 5570 1280 sw
rect 6059 1318 6061 1320
rect 6089 1318 6091 1320
rect 6059 1296 6091 1318
rect 6012 1268 6021 1296
rect 6051 1268 6099 1296
rect 6129 1268 6138 1296
tri 6138 1268 6150 1280 sw
rect 6639 1318 6641 1320
rect 6669 1318 6671 1320
rect 6639 1296 6671 1318
rect 6592 1268 6601 1296
rect 6631 1268 6679 1296
rect 6709 1268 6718 1296
tri 6718 1268 6730 1280 sw
rect 259 1048 261 1050
rect 289 1048 291 1050
rect 259 1026 291 1048
rect 212 998 221 1026
rect 251 998 299 1026
rect 329 998 338 1026
tri 338 998 350 1010 sw
rect 839 1048 841 1050
rect 869 1048 871 1050
rect 839 1026 871 1048
rect 792 998 801 1026
rect 831 998 879 1026
rect 909 998 918 1026
tri 918 998 930 1010 sw
rect 1419 1048 1421 1050
rect 1449 1048 1451 1050
rect 1419 1026 1451 1048
rect 1372 998 1381 1026
rect 1411 998 1459 1026
rect 1489 998 1498 1026
tri 1498 998 1510 1010 sw
rect 1999 1048 2001 1050
rect 2029 1048 2031 1050
rect 1999 1026 2031 1048
rect 1952 998 1961 1026
rect 1991 998 2039 1026
rect 2069 998 2078 1026
tri 2078 998 2090 1010 sw
rect 2579 1048 2581 1050
rect 2609 1048 2611 1050
rect 2579 1026 2611 1048
rect 2532 998 2541 1026
rect 2571 998 2619 1026
rect 2649 998 2658 1026
tri 2658 998 2670 1010 sw
rect 3159 1048 3161 1050
rect 3189 1048 3191 1050
rect 3159 1026 3191 1048
rect 3112 998 3121 1026
rect 3151 998 3199 1026
rect 3229 998 3238 1026
tri 3238 998 3250 1010 sw
rect 3739 1048 3741 1050
rect 3769 1048 3771 1050
rect 3739 1026 3771 1048
rect 3692 998 3701 1026
rect 3731 998 3779 1026
rect 3809 998 3818 1026
tri 3818 998 3830 1010 sw
rect 4319 1048 4321 1050
rect 4349 1048 4351 1050
rect 4319 1026 4351 1048
rect 4272 998 4281 1026
rect 4311 998 4359 1026
rect 4389 998 4398 1026
tri 4398 998 4410 1010 sw
rect 4899 1047 4901 1049
rect 4929 1047 4931 1049
rect 4899 1025 4931 1047
rect 4852 997 4861 1025
rect 4891 997 4939 1025
rect 4969 997 4978 1025
tri 4978 997 4990 1009 sw
rect 5479 1047 5481 1049
rect 5509 1047 5511 1049
rect 5479 1025 5511 1047
rect 5432 997 5441 1025
rect 5471 997 5519 1025
rect 5549 997 5558 1025
tri 5558 997 5570 1009 sw
rect 6059 1047 6061 1049
rect 6089 1047 6091 1049
rect 6059 1025 6091 1047
rect 6012 997 6021 1025
rect 6051 997 6099 1025
rect 6129 997 6138 1025
tri 6138 997 6150 1009 sw
rect 6639 1047 6641 1049
rect 6669 1047 6671 1049
rect 6639 1025 6671 1047
rect 6592 997 6601 1025
rect 6631 997 6679 1025
rect 6709 997 6718 1025
tri 6718 997 6730 1009 sw
rect 259 778 261 780
rect 289 778 291 780
rect 259 756 291 778
rect 212 728 221 756
rect 251 728 299 756
rect 329 728 338 756
tri 338 728 350 740 sw
rect 839 778 841 780
rect 869 778 871 780
rect 839 756 871 778
rect 792 728 801 756
rect 831 728 879 756
rect 909 728 918 756
tri 918 728 930 740 sw
rect 1419 778 1421 780
rect 1449 778 1451 780
rect 1419 756 1451 778
rect 1372 728 1381 756
rect 1411 728 1459 756
rect 1489 728 1498 756
tri 1498 728 1510 740 sw
rect 1999 778 2001 780
rect 2029 778 2031 780
rect 1999 756 2031 778
rect 1952 728 1961 756
rect 1991 728 2039 756
rect 2069 728 2078 756
tri 2078 728 2090 740 sw
rect 2579 778 2581 780
rect 2609 778 2611 780
rect 2579 756 2611 778
rect 2532 728 2541 756
rect 2571 728 2619 756
rect 2649 728 2658 756
tri 2658 728 2670 740 sw
rect 3159 778 3161 780
rect 3189 778 3191 780
rect 3159 756 3191 778
rect 3112 728 3121 756
rect 3151 728 3199 756
rect 3229 728 3238 756
tri 3238 728 3250 740 sw
rect 3739 778 3741 780
rect 3769 778 3771 780
rect 3739 756 3771 778
rect 3692 728 3701 756
rect 3731 728 3779 756
rect 3809 728 3818 756
tri 3818 728 3830 740 sw
rect 4319 778 4321 780
rect 4349 778 4351 780
rect 4319 756 4351 778
rect 4272 728 4281 756
rect 4311 728 4359 756
rect 4389 728 4398 756
tri 4398 728 4410 740 sw
rect 4899 777 4901 779
rect 4929 777 4931 779
rect 4899 755 4931 777
rect 4852 727 4861 755
rect 4891 727 4939 755
rect 4969 727 4978 755
tri 4978 727 4990 739 sw
rect 5479 777 5481 779
rect 5509 777 5511 779
rect 5479 755 5511 777
rect 5432 727 5441 755
rect 5471 727 5519 755
rect 5549 727 5558 755
tri 5558 727 5570 739 sw
rect 6059 777 6061 779
rect 6089 777 6091 779
rect 6059 755 6091 777
rect 6012 727 6021 755
rect 6051 727 6099 755
rect 6129 727 6138 755
tri 6138 727 6150 739 sw
rect 6639 777 6641 779
rect 6669 777 6671 779
rect 6639 755 6671 777
rect 6592 727 6601 755
rect 6631 727 6679 755
rect 6709 727 6718 755
tri 6718 727 6730 739 sw
rect 259 508 261 510
rect 289 508 291 510
rect 259 486 291 508
rect 212 458 221 486
rect 251 458 299 486
rect 329 458 338 486
tri 338 458 350 470 sw
rect 839 508 841 510
rect 869 508 871 510
rect 839 486 871 508
rect 792 458 801 486
rect 831 458 879 486
rect 909 458 918 486
tri 918 458 930 470 sw
rect 1419 508 1421 510
rect 1449 508 1451 510
rect 1419 486 1451 508
rect 1372 458 1381 486
rect 1411 458 1459 486
rect 1489 458 1498 486
tri 1498 458 1510 470 sw
rect 1999 508 2001 510
rect 2029 508 2031 510
rect 1999 486 2031 508
rect 1952 458 1961 486
rect 1991 458 2039 486
rect 2069 458 2078 486
tri 2078 458 2090 470 sw
rect 2579 508 2581 510
rect 2609 508 2611 510
rect 2579 486 2611 508
rect 2532 458 2541 486
rect 2571 458 2619 486
rect 2649 458 2658 486
tri 2658 458 2670 470 sw
rect 3159 508 3161 510
rect 3189 508 3191 510
rect 3159 486 3191 508
rect 3112 458 3121 486
rect 3151 458 3199 486
rect 3229 458 3238 486
tri 3238 458 3250 470 sw
rect 3739 508 3741 510
rect 3769 508 3771 510
rect 3739 486 3771 508
rect 3692 458 3701 486
rect 3731 458 3779 486
rect 3809 458 3818 486
tri 3818 458 3830 470 sw
rect 4319 508 4321 510
rect 4349 508 4351 510
rect 4319 486 4351 508
rect 4272 458 4281 486
rect 4311 458 4359 486
rect 4389 458 4398 486
tri 4398 458 4410 470 sw
rect 4899 507 4901 509
rect 4929 507 4931 509
rect 4899 485 4931 507
rect 4852 457 4861 485
rect 4891 457 4939 485
rect 4969 457 4978 485
tri 4978 457 4990 469 sw
rect 5479 507 5481 509
rect 5509 507 5511 509
rect 5479 485 5511 507
rect 5432 457 5441 485
rect 5471 457 5519 485
rect 5549 457 5558 485
tri 5558 457 5570 469 sw
rect 6059 507 6061 509
rect 6089 507 6091 509
rect 6059 485 6091 507
rect 6012 457 6021 485
rect 6051 457 6099 485
rect 6129 457 6138 485
tri 6138 457 6150 469 sw
rect 6639 507 6641 509
rect 6669 507 6671 509
rect 6639 485 6671 507
rect 6592 457 6601 485
rect 6631 457 6679 485
rect 6709 457 6718 485
tri 6718 457 6730 469 sw
rect 259 238 261 240
rect 289 238 291 240
rect 259 216 291 238
rect 212 188 221 216
rect 251 188 299 216
rect 329 188 338 216
tri 338 188 350 200 sw
rect 839 238 841 240
rect 869 238 871 240
rect 839 216 871 238
rect 792 188 801 216
rect 831 188 879 216
rect 909 188 918 216
tri 918 188 930 200 sw
rect 1419 238 1421 240
rect 1449 238 1451 240
rect 1419 216 1451 238
rect 1372 188 1381 216
rect 1411 188 1459 216
rect 1489 188 1498 216
tri 1498 188 1510 200 sw
rect 1999 238 2001 240
rect 2029 238 2031 240
rect 1999 216 2031 238
rect 1952 188 1961 216
rect 1991 188 2039 216
rect 2069 188 2078 216
tri 2078 188 2090 200 sw
rect 2579 238 2581 240
rect 2609 238 2611 240
rect 2579 216 2611 238
rect 2532 188 2541 216
rect 2571 188 2619 216
rect 2649 188 2658 216
tri 2658 188 2670 200 sw
rect 3159 238 3161 240
rect 3189 238 3191 240
rect 3159 216 3191 238
rect 3112 188 3121 216
rect 3151 188 3199 216
rect 3229 188 3238 216
tri 3238 188 3250 200 sw
rect 3739 238 3741 240
rect 3769 238 3771 240
rect 3739 216 3771 238
rect 3692 188 3701 216
rect 3731 188 3779 216
rect 3809 188 3818 216
tri 3818 188 3830 200 sw
rect 4319 238 4321 240
rect 4349 238 4351 240
rect 4319 216 4351 238
rect 4272 188 4281 216
rect 4311 188 4359 216
rect 4389 188 4398 216
tri 4398 188 4410 200 sw
rect 4899 237 4901 239
rect 4929 237 4931 239
rect 4899 215 4931 237
rect 4852 187 4861 215
rect 4891 187 4939 215
rect 4969 187 4978 215
tri 4978 187 4990 199 sw
rect 5479 237 5481 239
rect 5509 237 5511 239
rect 5479 215 5511 237
rect 5432 187 5441 215
rect 5471 187 5519 215
rect 5549 187 5558 215
tri 5558 187 5570 199 sw
rect 6059 237 6061 239
rect 6089 237 6091 239
rect 6059 215 6091 237
rect 6012 187 6021 215
rect 6051 187 6099 215
rect 6129 187 6138 215
tri 6138 187 6150 199 sw
rect 6639 237 6641 239
rect 6669 237 6671 239
rect 6639 215 6671 237
rect 6592 187 6601 215
rect 6631 187 6679 215
rect 6709 187 6718 215
tri 6718 187 6730 199 sw
rect 259 -32 261 -30
rect 289 -32 291 -30
rect 259 -54 291 -32
rect 212 -82 221 -54
rect 251 -82 299 -54
rect 329 -82 338 -54
tri 338 -82 350 -70 sw
rect 839 -32 841 -30
rect 869 -32 871 -30
rect 839 -54 871 -32
rect 792 -82 801 -54
rect 831 -82 879 -54
rect 909 -82 918 -54
tri 918 -82 930 -70 sw
rect 1419 -32 1421 -30
rect 1449 -32 1451 -30
rect 1419 -54 1451 -32
rect 1372 -82 1381 -54
rect 1411 -82 1459 -54
rect 1489 -82 1498 -54
tri 1498 -82 1510 -70 sw
rect 1999 -32 2001 -30
rect 2029 -32 2031 -30
rect 1999 -54 2031 -32
rect 1952 -82 1961 -54
rect 1991 -82 2039 -54
rect 2069 -82 2078 -54
tri 2078 -82 2090 -70 sw
rect 2579 -32 2581 -30
rect 2609 -32 2611 -30
rect 2579 -54 2611 -32
rect 2532 -82 2541 -54
rect 2571 -82 2619 -54
rect 2649 -82 2658 -54
tri 2658 -82 2670 -70 sw
rect 3159 -32 3161 -30
rect 3189 -32 3191 -30
rect 3159 -54 3191 -32
rect 3112 -82 3121 -54
rect 3151 -82 3199 -54
rect 3229 -82 3238 -54
tri 3238 -82 3250 -70 sw
rect 3739 -32 3741 -30
rect 3769 -32 3771 -30
rect 3739 -54 3771 -32
rect 3692 -82 3701 -54
rect 3731 -82 3779 -54
rect 3809 -82 3818 -54
tri 3818 -82 3830 -70 sw
rect 4319 -32 4321 -30
rect 4349 -32 4351 -30
rect 4319 -54 4351 -32
rect 4272 -82 4281 -54
rect 4311 -82 4359 -54
rect 4389 -82 4398 -54
tri 4398 -82 4410 -70 sw
rect 4899 -33 4901 -31
rect 4929 -33 4931 -31
rect 4899 -55 4931 -33
rect 4852 -83 4861 -55
rect 4891 -83 4939 -55
rect 4969 -83 4978 -55
tri 4978 -83 4990 -71 sw
rect 5479 -33 5481 -31
rect 5509 -33 5511 -31
rect 5479 -55 5511 -33
rect 5432 -83 5441 -55
rect 5471 -83 5519 -55
rect 5549 -83 5558 -55
tri 5558 -83 5570 -71 sw
rect 6059 -33 6061 -31
rect 6089 -33 6091 -31
rect 6059 -55 6091 -33
rect 6012 -83 6021 -55
rect 6051 -83 6099 -55
rect 6129 -83 6138 -55
tri 6138 -83 6150 -71 sw
rect 6639 -33 6641 -31
rect 6669 -33 6671 -31
rect 6639 -55 6671 -33
rect 6592 -83 6601 -55
rect 6631 -83 6679 -55
rect 6709 -83 6718 -55
tri 6718 -83 6730 -71 sw
rect 259 -302 261 -300
rect 289 -302 291 -300
rect 259 -324 291 -302
rect 212 -352 221 -324
rect 251 -352 299 -324
rect 329 -352 338 -324
tri 338 -352 350 -340 sw
rect 839 -302 841 -300
rect 869 -302 871 -300
rect 839 -324 871 -302
rect 792 -352 801 -324
rect 831 -352 879 -324
rect 909 -352 918 -324
tri 918 -352 930 -340 sw
rect 1419 -302 1421 -300
rect 1449 -302 1451 -300
rect 1419 -324 1451 -302
rect 1372 -352 1381 -324
rect 1411 -352 1459 -324
rect 1489 -352 1498 -324
tri 1498 -352 1510 -340 sw
rect 1999 -302 2001 -300
rect 2029 -302 2031 -300
rect 1999 -324 2031 -302
rect 1952 -352 1961 -324
rect 1991 -352 2039 -324
rect 2069 -352 2078 -324
tri 2078 -352 2090 -340 sw
rect 2579 -302 2581 -300
rect 2609 -302 2611 -300
rect 2579 -324 2611 -302
rect 2532 -352 2541 -324
rect 2571 -352 2619 -324
rect 2649 -352 2658 -324
tri 2658 -352 2670 -340 sw
rect 3159 -302 3161 -300
rect 3189 -302 3191 -300
rect 3159 -324 3191 -302
rect 3112 -352 3121 -324
rect 3151 -352 3199 -324
rect 3229 -352 3238 -324
tri 3238 -352 3250 -340 sw
rect 3739 -302 3741 -300
rect 3769 -302 3771 -300
rect 3739 -324 3771 -302
rect 3692 -352 3701 -324
rect 3731 -352 3779 -324
rect 3809 -352 3818 -324
tri 3818 -352 3830 -340 sw
rect 4319 -302 4321 -300
rect 4349 -302 4351 -300
rect 4319 -324 4351 -302
rect 4272 -352 4281 -324
rect 4311 -352 4359 -324
rect 4389 -352 4398 -324
tri 4398 -352 4410 -340 sw
rect 4899 -303 4901 -301
rect 4929 -303 4931 -301
rect 4899 -325 4931 -303
rect 4852 -353 4861 -325
rect 4891 -353 4939 -325
rect 4969 -353 4978 -325
tri 4978 -353 4990 -341 sw
rect 5479 -303 5481 -301
rect 5509 -303 5511 -301
rect 5479 -325 5511 -303
rect 5432 -353 5441 -325
rect 5471 -353 5519 -325
rect 5549 -353 5558 -325
tri 5558 -353 5570 -341 sw
rect 6059 -303 6061 -301
rect 6089 -303 6091 -301
rect 6059 -325 6091 -303
rect 6012 -353 6021 -325
rect 6051 -353 6099 -325
rect 6129 -353 6138 -325
tri 6138 -353 6150 -341 sw
rect 6639 -303 6641 -301
rect 6669 -303 6671 -301
rect 6639 -325 6671 -303
rect 6592 -353 6601 -325
rect 6631 -353 6679 -325
rect 6709 -353 6718 -325
tri 6718 -353 6730 -341 sw
rect 259 -572 261 -570
rect 289 -572 291 -570
rect 259 -594 291 -572
rect 212 -622 221 -594
rect 251 -622 299 -594
rect 329 -622 338 -594
tri 338 -622 350 -610 sw
rect 839 -572 841 -570
rect 869 -572 871 -570
rect 839 -594 871 -572
rect 792 -622 801 -594
rect 831 -622 879 -594
rect 909 -622 918 -594
tri 918 -622 930 -610 sw
rect 1419 -572 1421 -570
rect 1449 -572 1451 -570
rect 1419 -594 1451 -572
rect 1372 -622 1381 -594
rect 1411 -622 1459 -594
rect 1489 -622 1498 -594
tri 1498 -622 1510 -610 sw
rect 1999 -572 2001 -570
rect 2029 -572 2031 -570
rect 1999 -594 2031 -572
rect 1952 -622 1961 -594
rect 1991 -622 2039 -594
rect 2069 -622 2078 -594
tri 2078 -622 2090 -610 sw
rect 2579 -572 2581 -570
rect 2609 -572 2611 -570
rect 2579 -594 2611 -572
rect 2532 -622 2541 -594
rect 2571 -622 2619 -594
rect 2649 -622 2658 -594
tri 2658 -622 2670 -610 sw
rect 3159 -572 3161 -570
rect 3189 -572 3191 -570
rect 3159 -594 3191 -572
rect 3112 -622 3121 -594
rect 3151 -622 3199 -594
rect 3229 -622 3238 -594
tri 3238 -622 3250 -610 sw
rect 3739 -572 3741 -570
rect 3769 -572 3771 -570
rect 3739 -594 3771 -572
rect 3692 -622 3701 -594
rect 3731 -622 3779 -594
rect 3809 -622 3818 -594
tri 3818 -622 3830 -610 sw
rect 4319 -572 4321 -570
rect 4349 -572 4351 -570
rect 4319 -594 4351 -572
rect 4272 -622 4281 -594
rect 4311 -622 4359 -594
rect 4389 -622 4398 -594
tri 4398 -622 4410 -610 sw
rect 4899 -573 4901 -571
rect 4929 -573 4931 -571
rect 4899 -595 4931 -573
rect 4852 -623 4861 -595
rect 4891 -623 4939 -595
rect 4969 -623 4978 -595
tri 4978 -623 4990 -611 sw
rect 5479 -573 5481 -571
rect 5509 -573 5511 -571
rect 5479 -595 5511 -573
rect 5432 -623 5441 -595
rect 5471 -623 5519 -595
rect 5549 -623 5558 -595
tri 5558 -623 5570 -611 sw
rect 6059 -573 6061 -571
rect 6089 -573 6091 -571
rect 6059 -595 6091 -573
rect 6012 -623 6021 -595
rect 6051 -623 6099 -595
rect 6129 -623 6138 -595
tri 6138 -623 6150 -611 sw
rect 6639 -573 6641 -571
rect 6669 -573 6671 -571
rect 6639 -595 6671 -573
rect 6592 -623 6601 -595
rect 6631 -623 6679 -595
rect 6709 -623 6718 -595
tri 6718 -623 6730 -611 sw
rect 259 -842 261 -840
rect 289 -842 291 -840
rect 259 -864 291 -842
rect 212 -892 221 -864
rect 251 -892 299 -864
rect 329 -892 338 -864
tri 338 -892 350 -880 sw
rect 839 -842 841 -840
rect 869 -842 871 -840
rect 839 -864 871 -842
rect 792 -892 801 -864
rect 831 -892 879 -864
rect 909 -892 918 -864
tri 918 -892 930 -880 sw
rect 1419 -842 1421 -840
rect 1449 -842 1451 -840
rect 1419 -864 1451 -842
rect 1372 -892 1381 -864
rect 1411 -892 1459 -864
rect 1489 -892 1498 -864
tri 1498 -892 1510 -880 sw
rect 1999 -842 2001 -840
rect 2029 -842 2031 -840
rect 1999 -864 2031 -842
rect 1952 -892 1961 -864
rect 1991 -892 2039 -864
rect 2069 -892 2078 -864
tri 2078 -892 2090 -880 sw
rect 2579 -842 2581 -840
rect 2609 -842 2611 -840
rect 2579 -864 2611 -842
rect 2532 -892 2541 -864
rect 2571 -892 2619 -864
rect 2649 -892 2658 -864
tri 2658 -892 2670 -880 sw
rect 3159 -842 3161 -840
rect 3189 -842 3191 -840
rect 3159 -864 3191 -842
rect 3112 -892 3121 -864
rect 3151 -892 3199 -864
rect 3229 -892 3238 -864
tri 3238 -892 3250 -880 sw
rect 3739 -842 3741 -840
rect 3769 -842 3771 -840
rect 3739 -864 3771 -842
rect 3692 -892 3701 -864
rect 3731 -892 3779 -864
rect 3809 -892 3818 -864
tri 3818 -892 3830 -880 sw
rect 4319 -842 4321 -840
rect 4349 -842 4351 -840
rect 4319 -864 4351 -842
rect 4272 -892 4281 -864
rect 4311 -892 4359 -864
rect 4389 -892 4398 -864
tri 4398 -892 4410 -880 sw
rect 4899 -843 4901 -841
rect 4929 -843 4931 -841
rect 4899 -865 4931 -843
rect 4852 -893 4861 -865
rect 4891 -893 4939 -865
rect 4969 -893 4978 -865
tri 4978 -893 4990 -881 sw
rect 5479 -843 5481 -841
rect 5509 -843 5511 -841
rect 5479 -865 5511 -843
rect 5432 -893 5441 -865
rect 5471 -893 5519 -865
rect 5549 -893 5558 -865
tri 5558 -893 5570 -881 sw
rect 6059 -843 6061 -841
rect 6089 -843 6091 -841
rect 6059 -865 6091 -843
rect 6012 -893 6021 -865
rect 6051 -893 6099 -865
rect 6129 -893 6138 -865
tri 6138 -893 6150 -881 sw
rect 6639 -843 6641 -841
rect 6669 -843 6671 -841
rect 6639 -865 6671 -843
rect 6592 -893 6601 -865
rect 6631 -893 6679 -865
rect 6709 -893 6718 -865
tri 6718 -893 6730 -881 sw
rect 259 -1112 261 -1110
rect 289 -1112 291 -1110
rect 259 -1134 291 -1112
rect 212 -1162 221 -1134
rect 251 -1162 299 -1134
rect 329 -1162 338 -1134
tri 338 -1162 350 -1150 sw
rect 839 -1112 841 -1110
rect 869 -1112 871 -1110
rect 839 -1134 871 -1112
rect 792 -1162 801 -1134
rect 831 -1162 879 -1134
rect 909 -1162 918 -1134
tri 918 -1162 930 -1150 sw
rect 1419 -1112 1421 -1110
rect 1449 -1112 1451 -1110
rect 1419 -1134 1451 -1112
rect 1372 -1162 1381 -1134
rect 1411 -1162 1459 -1134
rect 1489 -1162 1498 -1134
tri 1498 -1162 1510 -1150 sw
rect 1999 -1112 2001 -1110
rect 2029 -1112 2031 -1110
rect 1999 -1134 2031 -1112
rect 1952 -1162 1961 -1134
rect 1991 -1162 2039 -1134
rect 2069 -1162 2078 -1134
tri 2078 -1162 2090 -1150 sw
rect 2579 -1112 2581 -1110
rect 2609 -1112 2611 -1110
rect 2579 -1134 2611 -1112
rect 2532 -1162 2541 -1134
rect 2571 -1162 2619 -1134
rect 2649 -1162 2658 -1134
tri 2658 -1162 2670 -1150 sw
rect 3159 -1112 3161 -1110
rect 3189 -1112 3191 -1110
rect 3159 -1134 3191 -1112
rect 3112 -1162 3121 -1134
rect 3151 -1162 3199 -1134
rect 3229 -1162 3238 -1134
tri 3238 -1162 3250 -1150 sw
rect 3739 -1112 3741 -1110
rect 3769 -1112 3771 -1110
rect 3739 -1134 3771 -1112
rect 3692 -1162 3701 -1134
rect 3731 -1162 3779 -1134
rect 3809 -1162 3818 -1134
tri 3818 -1162 3830 -1150 sw
rect 4319 -1112 4321 -1110
rect 4349 -1112 4351 -1110
rect 4319 -1134 4351 -1112
rect 4272 -1162 4281 -1134
rect 4311 -1162 4359 -1134
rect 4389 -1162 4398 -1134
tri 4398 -1162 4410 -1150 sw
rect 4899 -1113 4901 -1111
rect 4929 -1113 4931 -1111
rect 4899 -1135 4931 -1113
rect 4852 -1163 4861 -1135
rect 4891 -1163 4939 -1135
rect 4969 -1163 4978 -1135
tri 4978 -1163 4990 -1151 sw
rect 5479 -1113 5481 -1111
rect 5509 -1113 5511 -1111
rect 5479 -1135 5511 -1113
rect 5432 -1163 5441 -1135
rect 5471 -1163 5519 -1135
rect 5549 -1163 5558 -1135
tri 5558 -1163 5570 -1151 sw
rect 6059 -1113 6061 -1111
rect 6089 -1113 6091 -1111
rect 6059 -1135 6091 -1113
rect 6012 -1163 6021 -1135
rect 6051 -1163 6099 -1135
rect 6129 -1163 6138 -1135
tri 6138 -1163 6150 -1151 sw
rect 6639 -1113 6641 -1111
rect 6669 -1113 6671 -1111
rect 6639 -1135 6671 -1113
rect 6592 -1163 6601 -1135
rect 6631 -1163 6679 -1135
rect 6709 -1163 6718 -1135
tri 6718 -1163 6730 -1151 sw
rect 259 -1382 261 -1380
rect 289 -1382 291 -1380
rect 259 -1404 291 -1382
rect 212 -1432 221 -1404
rect 251 -1432 299 -1404
rect 329 -1432 338 -1404
tri 338 -1432 350 -1420 sw
rect 839 -1382 841 -1380
rect 869 -1382 871 -1380
rect 839 -1404 871 -1382
rect 792 -1432 801 -1404
rect 831 -1432 879 -1404
rect 909 -1432 918 -1404
tri 918 -1432 930 -1420 sw
rect 1419 -1382 1421 -1380
rect 1449 -1382 1451 -1380
rect 1419 -1404 1451 -1382
rect 1372 -1432 1381 -1404
rect 1411 -1432 1459 -1404
rect 1489 -1432 1498 -1404
tri 1498 -1432 1510 -1420 sw
rect 1999 -1382 2001 -1380
rect 2029 -1382 2031 -1380
rect 1999 -1404 2031 -1382
rect 1952 -1432 1961 -1404
rect 1991 -1432 2039 -1404
rect 2069 -1432 2078 -1404
tri 2078 -1432 2090 -1420 sw
rect 2579 -1382 2581 -1380
rect 2609 -1382 2611 -1380
rect 2579 -1404 2611 -1382
rect 2532 -1432 2541 -1404
rect 2571 -1432 2619 -1404
rect 2649 -1432 2658 -1404
tri 2658 -1432 2670 -1420 sw
rect 3159 -1382 3161 -1380
rect 3189 -1382 3191 -1380
rect 3159 -1404 3191 -1382
rect 3112 -1432 3121 -1404
rect 3151 -1432 3199 -1404
rect 3229 -1432 3238 -1404
tri 3238 -1432 3250 -1420 sw
rect 3739 -1382 3741 -1380
rect 3769 -1382 3771 -1380
rect 3739 -1404 3771 -1382
rect 3692 -1432 3701 -1404
rect 3731 -1432 3779 -1404
rect 3809 -1432 3818 -1404
tri 3818 -1432 3830 -1420 sw
rect 4319 -1382 4321 -1380
rect 4349 -1382 4351 -1380
rect 4319 -1404 4351 -1382
rect 4272 -1432 4281 -1404
rect 4311 -1432 4359 -1404
rect 4389 -1432 4398 -1404
tri 4398 -1432 4410 -1420 sw
rect 4899 -1383 4901 -1381
rect 4929 -1383 4931 -1381
rect 4899 -1405 4931 -1383
rect 4852 -1433 4861 -1405
rect 4891 -1433 4939 -1405
rect 4969 -1433 4978 -1405
tri 4978 -1433 4990 -1421 sw
rect 5479 -1383 5481 -1381
rect 5509 -1383 5511 -1381
rect 5479 -1405 5511 -1383
rect 5432 -1433 5441 -1405
rect 5471 -1433 5519 -1405
rect 5549 -1433 5558 -1405
tri 5558 -1433 5570 -1421 sw
rect 6059 -1383 6061 -1381
rect 6089 -1383 6091 -1381
rect 6059 -1405 6091 -1383
rect 6012 -1433 6021 -1405
rect 6051 -1433 6099 -1405
rect 6129 -1433 6138 -1405
tri 6138 -1433 6150 -1421 sw
rect 6639 -1383 6641 -1381
rect 6669 -1383 6671 -1381
rect 6639 -1405 6671 -1383
rect 6592 -1433 6601 -1405
rect 6631 -1433 6679 -1405
rect 6709 -1433 6718 -1405
tri 6718 -1433 6730 -1421 sw
rect 259 -1652 261 -1650
rect 289 -1652 291 -1650
rect 259 -1674 291 -1652
rect 212 -1702 221 -1674
rect 251 -1702 299 -1674
rect 329 -1702 338 -1674
tri 338 -1702 350 -1690 sw
rect 839 -1652 841 -1650
rect 869 -1652 871 -1650
rect 839 -1674 871 -1652
rect 792 -1702 801 -1674
rect 831 -1702 879 -1674
rect 909 -1702 918 -1674
tri 918 -1702 930 -1690 sw
rect 1419 -1652 1421 -1650
rect 1449 -1652 1451 -1650
rect 1419 -1674 1451 -1652
rect 1372 -1702 1381 -1674
rect 1411 -1702 1459 -1674
rect 1489 -1702 1498 -1674
tri 1498 -1702 1510 -1690 sw
rect 1999 -1652 2001 -1650
rect 2029 -1652 2031 -1650
rect 1999 -1674 2031 -1652
rect 1952 -1702 1961 -1674
rect 1991 -1702 2039 -1674
rect 2069 -1702 2078 -1674
tri 2078 -1702 2090 -1690 sw
rect 2579 -1652 2581 -1650
rect 2609 -1652 2611 -1650
rect 2579 -1674 2611 -1652
rect 2532 -1702 2541 -1674
rect 2571 -1702 2619 -1674
rect 2649 -1702 2658 -1674
tri 2658 -1702 2670 -1690 sw
rect 3159 -1652 3161 -1650
rect 3189 -1652 3191 -1650
rect 3159 -1674 3191 -1652
rect 3112 -1702 3121 -1674
rect 3151 -1702 3199 -1674
rect 3229 -1702 3238 -1674
tri 3238 -1702 3250 -1690 sw
rect 3739 -1652 3741 -1650
rect 3769 -1652 3771 -1650
rect 3739 -1674 3771 -1652
rect 3692 -1702 3701 -1674
rect 3731 -1702 3779 -1674
rect 3809 -1702 3818 -1674
tri 3818 -1702 3830 -1690 sw
rect 4319 -1652 4321 -1650
rect 4349 -1652 4351 -1650
rect 4319 -1674 4351 -1652
rect 4272 -1702 4281 -1674
rect 4311 -1702 4359 -1674
rect 4389 -1702 4398 -1674
tri 4398 -1702 4410 -1690 sw
rect 4899 -1653 4901 -1651
rect 4929 -1653 4931 -1651
rect 4899 -1675 4931 -1653
rect 4852 -1703 4861 -1675
rect 4891 -1703 4939 -1675
rect 4969 -1703 4978 -1675
tri 4978 -1703 4990 -1691 sw
rect 5479 -1653 5481 -1651
rect 5509 -1653 5511 -1651
rect 5479 -1675 5511 -1653
rect 5432 -1703 5441 -1675
rect 5471 -1703 5519 -1675
rect 5549 -1703 5558 -1675
tri 5558 -1703 5570 -1691 sw
rect 6059 -1653 6061 -1651
rect 6089 -1653 6091 -1651
rect 6059 -1675 6091 -1653
rect 6012 -1703 6021 -1675
rect 6051 -1703 6099 -1675
rect 6129 -1703 6138 -1675
tri 6138 -1703 6150 -1691 sw
rect 6639 -1653 6641 -1651
rect 6669 -1653 6671 -1651
rect 6639 -1675 6671 -1653
rect 6592 -1703 6601 -1675
rect 6631 -1703 6679 -1675
rect 6709 -1703 6718 -1675
tri 6718 -1703 6730 -1691 sw
rect 259 -1922 261 -1920
rect 289 -1922 291 -1920
rect 259 -1944 291 -1922
rect 212 -1972 221 -1944
rect 251 -1972 299 -1944
rect 329 -1972 338 -1944
tri 338 -1972 350 -1960 sw
rect 839 -1922 841 -1920
rect 869 -1922 871 -1920
rect 839 -1944 871 -1922
rect 792 -1972 801 -1944
rect 831 -1972 879 -1944
rect 909 -1972 918 -1944
tri 918 -1972 930 -1960 sw
rect 1419 -1922 1421 -1920
rect 1449 -1922 1451 -1920
rect 1419 -1944 1451 -1922
rect 1372 -1972 1381 -1944
rect 1411 -1972 1459 -1944
rect 1489 -1972 1498 -1944
tri 1498 -1972 1510 -1960 sw
rect 1999 -1922 2001 -1920
rect 2029 -1922 2031 -1920
rect 1999 -1944 2031 -1922
rect 1952 -1972 1961 -1944
rect 1991 -1972 2039 -1944
rect 2069 -1972 2078 -1944
tri 2078 -1972 2090 -1960 sw
rect 2579 -1922 2581 -1920
rect 2609 -1922 2611 -1920
rect 2579 -1944 2611 -1922
rect 2532 -1972 2541 -1944
rect 2571 -1972 2619 -1944
rect 2649 -1972 2658 -1944
tri 2658 -1972 2670 -1960 sw
rect 3159 -1922 3161 -1920
rect 3189 -1922 3191 -1920
rect 3159 -1944 3191 -1922
rect 3112 -1972 3121 -1944
rect 3151 -1972 3199 -1944
rect 3229 -1972 3238 -1944
tri 3238 -1972 3250 -1960 sw
rect 3739 -1922 3741 -1920
rect 3769 -1922 3771 -1920
rect 3739 -1944 3771 -1922
rect 3692 -1972 3701 -1944
rect 3731 -1972 3779 -1944
rect 3809 -1972 3818 -1944
tri 3818 -1972 3830 -1960 sw
rect 4319 -1922 4321 -1920
rect 4349 -1922 4351 -1920
rect 4319 -1944 4351 -1922
rect 4272 -1972 4281 -1944
rect 4311 -1972 4359 -1944
rect 4389 -1972 4398 -1944
tri 4398 -1972 4410 -1960 sw
rect 4899 -1923 4901 -1921
rect 4929 -1923 4931 -1921
rect 4899 -1945 4931 -1923
rect 4852 -1973 4861 -1945
rect 4891 -1973 4939 -1945
rect 4969 -1973 4978 -1945
tri 4978 -1973 4990 -1961 sw
rect 5479 -1923 5481 -1921
rect 5509 -1923 5511 -1921
rect 5479 -1945 5511 -1923
rect 5432 -1973 5441 -1945
rect 5471 -1973 5519 -1945
rect 5549 -1973 5558 -1945
tri 5558 -1973 5570 -1961 sw
rect 6059 -1923 6061 -1921
rect 6089 -1923 6091 -1921
rect 6059 -1945 6091 -1923
rect 6012 -1973 6021 -1945
rect 6051 -1973 6099 -1945
rect 6129 -1973 6138 -1945
tri 6138 -1973 6150 -1961 sw
rect 6639 -1923 6641 -1921
rect 6669 -1923 6671 -1921
rect 6639 -1945 6671 -1923
rect 6592 -1973 6601 -1945
rect 6631 -1973 6679 -1945
rect 6709 -1973 6718 -1945
tri 6718 -1973 6730 -1961 sw
<< ndiffc >>
rect 73 2088 88 2116
rect 154 2088 169 2116
rect 381 2088 396 2116
rect 463 2088 478 2117
rect 653 2088 668 2116
rect 734 2088 749 2116
rect 961 2088 976 2116
rect 1043 2088 1058 2117
rect 1233 2088 1248 2116
rect 1314 2088 1329 2116
rect 1541 2088 1556 2116
rect 1623 2088 1638 2117
rect 1813 2088 1828 2116
rect 1894 2088 1909 2116
rect 2121 2088 2136 2116
rect 2203 2088 2218 2117
rect 2393 2088 2408 2116
rect 2474 2088 2489 2116
rect 2701 2088 2716 2116
rect 2783 2088 2798 2117
rect 2973 2088 2988 2116
rect 3054 2088 3069 2116
rect 3281 2088 3296 2116
rect 3363 2088 3378 2117
rect 3553 2088 3568 2116
rect 3634 2088 3649 2116
rect 3861 2088 3876 2116
rect 3943 2088 3958 2117
rect 4133 2088 4148 2116
rect 4214 2088 4229 2116
rect 4441 2088 4456 2116
rect 4523 2088 4538 2117
rect 4713 2088 4728 2116
rect 4794 2088 4809 2116
rect 5021 2088 5036 2116
rect 5103 2088 5118 2117
rect 5293 2088 5308 2116
rect 5374 2088 5389 2116
rect 5601 2088 5616 2116
rect 5683 2088 5698 2117
rect 5873 2088 5888 2116
rect 5954 2088 5969 2116
rect 6181 2088 6196 2116
rect 6263 2088 6278 2117
rect 6453 2088 6468 2116
rect 6534 2088 6549 2116
rect 6761 2088 6776 2116
rect 6843 2088 6858 2117
rect -1 1942 14 1984
rect 196 1967 206 1974
tri 206 1967 213 1974 sw
rect 196 1942 213 1967
rect 337 1942 354 1974
rect 536 1942 551 1984
rect 579 1942 594 1984
rect 776 1967 786 1974
tri 786 1967 793 1974 sw
rect 776 1942 793 1967
rect 917 1942 934 1974
rect 1116 1942 1131 1984
rect 1159 1942 1174 1984
rect 1356 1967 1366 1974
tri 1366 1967 1373 1974 sw
rect 1356 1942 1373 1967
rect 1497 1942 1514 1974
rect 1696 1942 1711 1984
rect 1739 1942 1754 1984
rect 1936 1967 1946 1974
tri 1946 1967 1953 1974 sw
rect 1936 1942 1953 1967
rect 2077 1942 2094 1974
rect 2276 1942 2291 1984
rect 2319 1942 2334 1984
rect 2516 1967 2526 1974
tri 2526 1967 2533 1974 sw
rect 2516 1942 2533 1967
rect 2657 1942 2674 1974
rect 2856 1942 2871 1984
rect 2899 1942 2914 1984
rect 3096 1967 3106 1974
tri 3106 1967 3113 1974 sw
rect 3096 1942 3113 1967
rect 3237 1942 3254 1974
rect 3436 1942 3451 1984
rect 3479 1942 3494 1984
rect 3676 1967 3686 1974
tri 3686 1967 3693 1974 sw
rect 3676 1942 3693 1967
rect 3817 1942 3834 1974
rect 4016 1942 4031 1984
rect 4059 1942 4074 1984
rect 4256 1967 4266 1974
tri 4266 1967 4273 1974 sw
rect 4256 1942 4273 1967
rect 4397 1942 4414 1974
rect 4596 1942 4611 1984
rect 4639 1942 4654 1984
rect 4836 1967 4846 1974
tri 4846 1967 4853 1974 sw
rect 4836 1942 4853 1967
rect 4977 1942 4994 1974
rect 5176 1942 5191 1984
rect 5219 1942 5234 1984
rect 5416 1967 5426 1974
tri 5426 1967 5433 1974 sw
rect 5416 1942 5433 1967
rect 5557 1942 5574 1974
rect 5756 1942 5771 1984
rect 5799 1942 5814 1984
rect 5996 1967 6006 1974
tri 6006 1967 6013 1974 sw
rect 5996 1942 6013 1967
rect 6137 1942 6154 1974
rect 6336 1942 6351 1984
rect 6379 1942 6394 1984
rect 6576 1967 6586 1974
tri 6586 1967 6593 1974 sw
rect 6576 1942 6593 1967
rect 6717 1942 6734 1974
rect 6916 1942 6931 1984
rect 259 1904 291 1918
rect 839 1904 871 1918
rect 1419 1904 1451 1918
rect 1999 1904 2031 1918
rect 2579 1904 2611 1918
rect 3159 1904 3191 1918
rect 3739 1904 3771 1918
rect 4319 1904 4351 1918
rect 4899 1904 4931 1918
rect 5479 1904 5511 1918
rect 6059 1904 6091 1918
rect 6639 1904 6671 1918
rect 73 1818 88 1846
rect 154 1818 169 1846
rect 381 1818 396 1846
rect 463 1818 478 1847
rect 653 1818 668 1846
rect 734 1818 749 1846
rect 961 1818 976 1846
rect 1043 1818 1058 1847
rect 1233 1818 1248 1846
rect 1314 1818 1329 1846
rect 1541 1818 1556 1846
rect 1623 1818 1638 1847
rect 1813 1818 1828 1846
rect 1894 1818 1909 1846
rect 2121 1818 2136 1846
rect 2203 1818 2218 1847
rect 2393 1818 2408 1846
rect 2474 1818 2489 1846
rect 2701 1818 2716 1846
rect 2783 1818 2798 1847
rect 2973 1818 2988 1846
rect 3054 1818 3069 1846
rect 3281 1818 3296 1846
rect 3363 1818 3378 1847
rect 3553 1818 3568 1846
rect 3634 1818 3649 1846
rect 3861 1818 3876 1846
rect 3943 1818 3958 1847
rect 4133 1818 4148 1846
rect 4214 1818 4229 1846
rect 4441 1818 4456 1846
rect 4523 1818 4538 1847
rect 4713 1818 4728 1846
rect 4794 1818 4809 1846
rect 5021 1818 5036 1846
rect 5103 1818 5118 1847
rect 5293 1818 5308 1846
rect 5374 1818 5389 1846
rect 5601 1818 5616 1846
rect 5683 1818 5698 1847
rect 5873 1818 5888 1846
rect 5954 1818 5969 1846
rect 6181 1818 6196 1846
rect 6263 1818 6278 1847
rect 6453 1818 6468 1846
rect 6534 1818 6549 1846
rect 6761 1818 6776 1846
rect 6843 1818 6858 1847
rect -1 1672 14 1714
rect 196 1697 206 1704
tri 206 1697 213 1704 sw
rect 196 1672 213 1697
rect 337 1672 354 1704
rect 536 1672 551 1714
rect 579 1672 594 1714
rect 776 1697 786 1704
tri 786 1697 793 1704 sw
rect 776 1672 793 1697
rect 917 1672 934 1704
rect 1116 1672 1131 1714
rect 1159 1672 1174 1714
rect 1356 1697 1366 1704
tri 1366 1697 1373 1704 sw
rect 1356 1672 1373 1697
rect 1497 1672 1514 1704
rect 1696 1672 1711 1714
rect 1739 1672 1754 1714
rect 1936 1697 1946 1704
tri 1946 1697 1953 1704 sw
rect 1936 1672 1953 1697
rect 2077 1672 2094 1704
rect 2276 1672 2291 1714
rect 2319 1672 2334 1714
rect 2516 1697 2526 1704
tri 2526 1697 2533 1704 sw
rect 2516 1672 2533 1697
rect 2657 1672 2674 1704
rect 2856 1672 2871 1714
rect 2899 1672 2914 1714
rect 3096 1697 3106 1704
tri 3106 1697 3113 1704 sw
rect 3096 1672 3113 1697
rect 3237 1672 3254 1704
rect 3436 1672 3451 1714
rect 3479 1672 3494 1714
rect 3676 1697 3686 1704
tri 3686 1697 3693 1704 sw
rect 3676 1672 3693 1697
rect 3817 1672 3834 1704
rect 4016 1672 4031 1714
rect 4059 1672 4074 1714
rect 4256 1697 4266 1704
tri 4266 1697 4273 1704 sw
rect 4256 1672 4273 1697
rect 4397 1672 4414 1704
rect 4596 1672 4611 1714
rect 4639 1672 4654 1714
rect 4836 1697 4846 1704
tri 4846 1697 4853 1704 sw
rect 4836 1672 4853 1697
rect 4977 1672 4994 1704
rect 5176 1672 5191 1714
rect 5219 1672 5234 1714
rect 5416 1697 5426 1704
tri 5426 1697 5433 1704 sw
rect 5416 1672 5433 1697
rect 5557 1672 5574 1704
rect 5756 1672 5771 1714
rect 5799 1672 5814 1714
rect 5996 1697 6006 1704
tri 6006 1697 6013 1704 sw
rect 5996 1672 6013 1697
rect 6137 1672 6154 1704
rect 6336 1672 6351 1714
rect 6379 1672 6394 1714
rect 6576 1697 6586 1704
tri 6586 1697 6593 1704 sw
rect 6576 1672 6593 1697
rect 6717 1672 6734 1704
rect 6916 1672 6931 1714
rect 259 1634 291 1648
rect 839 1634 871 1648
rect 1419 1634 1451 1648
rect 1999 1634 2031 1648
rect 2579 1634 2611 1648
rect 3159 1634 3191 1648
rect 3739 1634 3771 1648
rect 4319 1634 4351 1648
rect 4899 1634 4931 1648
rect 5479 1634 5511 1648
rect 6059 1634 6091 1648
rect 6639 1634 6671 1648
rect 73 1548 88 1576
rect 154 1548 169 1576
rect 381 1548 396 1576
rect 463 1548 478 1577
rect 653 1548 668 1576
rect 734 1548 749 1576
rect 961 1548 976 1576
rect 1043 1548 1058 1577
rect 1233 1548 1248 1576
rect 1314 1548 1329 1576
rect 1541 1548 1556 1576
rect 1623 1548 1638 1577
rect 1813 1548 1828 1576
rect 1894 1548 1909 1576
rect 2121 1548 2136 1576
rect 2203 1548 2218 1577
rect 2393 1548 2408 1576
rect 2474 1548 2489 1576
rect 2701 1548 2716 1576
rect 2783 1548 2798 1577
rect 2973 1548 2988 1576
rect 3054 1548 3069 1576
rect 3281 1548 3296 1576
rect 3363 1548 3378 1577
rect 3553 1548 3568 1576
rect 3634 1548 3649 1576
rect 3861 1548 3876 1576
rect 3943 1548 3958 1577
rect 4133 1548 4148 1576
rect 4214 1548 4229 1576
rect 4441 1548 4456 1576
rect 4523 1548 4538 1577
rect 4713 1548 4728 1576
rect 4794 1548 4809 1576
rect 5021 1548 5036 1576
rect 5103 1548 5118 1577
rect 5293 1548 5308 1576
rect 5374 1548 5389 1576
rect 5601 1548 5616 1576
rect 5683 1548 5698 1577
rect 5873 1548 5888 1576
rect 5954 1548 5969 1576
rect 6181 1548 6196 1576
rect 6263 1548 6278 1577
rect 6453 1548 6468 1576
rect 6534 1548 6549 1576
rect 6761 1548 6776 1576
rect 6843 1548 6858 1577
rect -1 1402 14 1444
rect 196 1427 206 1434
tri 206 1427 213 1434 sw
rect 196 1402 213 1427
rect 337 1402 354 1434
rect 536 1402 551 1444
rect 579 1402 594 1444
rect 776 1427 786 1434
tri 786 1427 793 1434 sw
rect 776 1402 793 1427
rect 917 1402 934 1434
rect 1116 1402 1131 1444
rect 1159 1402 1174 1444
rect 1356 1427 1366 1434
tri 1366 1427 1373 1434 sw
rect 1356 1402 1373 1427
rect 1497 1402 1514 1434
rect 1696 1402 1711 1444
rect 1739 1402 1754 1444
rect 1936 1427 1946 1434
tri 1946 1427 1953 1434 sw
rect 1936 1402 1953 1427
rect 2077 1402 2094 1434
rect 2276 1402 2291 1444
rect 2319 1402 2334 1444
rect 2516 1427 2526 1434
tri 2526 1427 2533 1434 sw
rect 2516 1402 2533 1427
rect 2657 1402 2674 1434
rect 2856 1402 2871 1444
rect 2899 1402 2914 1444
rect 3096 1427 3106 1434
tri 3106 1427 3113 1434 sw
rect 3096 1402 3113 1427
rect 3237 1402 3254 1434
rect 3436 1402 3451 1444
rect 3479 1402 3494 1444
rect 3676 1427 3686 1434
tri 3686 1427 3693 1434 sw
rect 3676 1402 3693 1427
rect 3817 1402 3834 1434
rect 4016 1402 4031 1444
rect 4059 1402 4074 1444
rect 4256 1427 4266 1434
tri 4266 1427 4273 1434 sw
rect 4256 1402 4273 1427
rect 4397 1402 4414 1434
rect 4596 1402 4611 1444
rect 4639 1402 4654 1444
rect 4836 1427 4846 1434
tri 4846 1427 4853 1434 sw
rect 4836 1402 4853 1427
rect 4977 1402 4994 1434
rect 5176 1402 5191 1444
rect 5219 1402 5234 1444
rect 5416 1427 5426 1434
tri 5426 1427 5433 1434 sw
rect 5416 1402 5433 1427
rect 5557 1402 5574 1434
rect 5756 1402 5771 1444
rect 5799 1402 5814 1444
rect 5996 1427 6006 1434
tri 6006 1427 6013 1434 sw
rect 5996 1402 6013 1427
rect 6137 1402 6154 1434
rect 6336 1402 6351 1444
rect 6379 1402 6394 1444
rect 6576 1427 6586 1434
tri 6586 1427 6593 1434 sw
rect 6576 1402 6593 1427
rect 6717 1402 6734 1434
rect 6916 1402 6931 1444
rect 259 1364 291 1378
rect 839 1364 871 1378
rect 1419 1364 1451 1378
rect 1999 1364 2031 1378
rect 2579 1364 2611 1378
rect 3159 1364 3191 1378
rect 3739 1364 3771 1378
rect 4319 1364 4351 1378
rect 4899 1364 4931 1378
rect 5479 1364 5511 1378
rect 6059 1364 6091 1378
rect 6639 1364 6671 1378
rect 73 1278 88 1306
rect 154 1278 169 1306
rect 381 1278 396 1306
rect 463 1278 478 1307
rect 653 1278 668 1306
rect 734 1278 749 1306
rect 961 1278 976 1306
rect 1043 1278 1058 1307
rect 1233 1278 1248 1306
rect 1314 1278 1329 1306
rect 1541 1278 1556 1306
rect 1623 1278 1638 1307
rect 1813 1278 1828 1306
rect 1894 1278 1909 1306
rect 2121 1278 2136 1306
rect 2203 1278 2218 1307
rect 2393 1278 2408 1306
rect 2474 1278 2489 1306
rect 2701 1278 2716 1306
rect 2783 1278 2798 1307
rect 2973 1278 2988 1306
rect 3054 1278 3069 1306
rect 3281 1278 3296 1306
rect 3363 1278 3378 1307
rect 3553 1278 3568 1306
rect 3634 1278 3649 1306
rect 3861 1278 3876 1306
rect 3943 1278 3958 1307
rect 4133 1278 4148 1306
rect 4214 1278 4229 1306
rect 4441 1278 4456 1306
rect 4523 1278 4538 1307
rect 4713 1278 4728 1306
rect 4794 1278 4809 1306
rect 5021 1278 5036 1306
rect 5103 1278 5118 1307
rect 5293 1278 5308 1306
rect 5374 1278 5389 1306
rect 5601 1278 5616 1306
rect 5683 1278 5698 1307
rect 5873 1278 5888 1306
rect 5954 1278 5969 1306
rect 6181 1278 6196 1306
rect 6263 1278 6278 1307
rect 6453 1278 6468 1306
rect 6534 1278 6549 1306
rect 6761 1278 6776 1306
rect 6843 1278 6858 1307
rect -1 1132 14 1174
rect 196 1157 206 1164
tri 206 1157 213 1164 sw
rect 196 1132 213 1157
rect 337 1132 354 1164
rect 536 1132 551 1174
rect 579 1132 594 1174
rect 776 1157 786 1164
tri 786 1157 793 1164 sw
rect 776 1132 793 1157
rect 917 1132 934 1164
rect 1116 1132 1131 1174
rect 1159 1132 1174 1174
rect 1356 1157 1366 1164
tri 1366 1157 1373 1164 sw
rect 1356 1132 1373 1157
rect 1497 1132 1514 1164
rect 1696 1132 1711 1174
rect 1739 1132 1754 1174
rect 1936 1157 1946 1164
tri 1946 1157 1953 1164 sw
rect 1936 1132 1953 1157
rect 2077 1132 2094 1164
rect 2276 1132 2291 1174
rect 2319 1132 2334 1174
rect 2516 1157 2526 1164
tri 2526 1157 2533 1164 sw
rect 2516 1132 2533 1157
rect 2657 1132 2674 1164
rect 2856 1132 2871 1174
rect 2899 1132 2914 1174
rect 3096 1157 3106 1164
tri 3106 1157 3113 1164 sw
rect 3096 1132 3113 1157
rect 3237 1132 3254 1164
rect 3436 1132 3451 1174
rect 3479 1132 3494 1174
rect 3676 1157 3686 1164
tri 3686 1157 3693 1164 sw
rect 3676 1132 3693 1157
rect 3817 1132 3834 1164
rect 4016 1132 4031 1174
rect 4059 1132 4074 1174
rect 4256 1157 4266 1164
tri 4266 1157 4273 1164 sw
rect 4256 1132 4273 1157
rect 4397 1132 4414 1164
rect 4596 1132 4611 1174
rect 4639 1132 4654 1174
rect 4836 1157 4846 1164
tri 4846 1157 4853 1164 sw
rect 4836 1132 4853 1157
rect 4977 1132 4994 1164
rect 5176 1132 5191 1174
rect 5219 1132 5234 1174
rect 5416 1157 5426 1164
tri 5426 1157 5433 1164 sw
rect 5416 1132 5433 1157
rect 5557 1132 5574 1164
rect 5756 1132 5771 1174
rect 5799 1132 5814 1174
rect 5996 1157 6006 1164
tri 6006 1157 6013 1164 sw
rect 5996 1132 6013 1157
rect 6137 1132 6154 1164
rect 6336 1132 6351 1174
rect 6379 1132 6394 1174
rect 6576 1157 6586 1164
tri 6586 1157 6593 1164 sw
rect 6576 1132 6593 1157
rect 6717 1132 6734 1164
rect 6916 1132 6931 1174
rect 259 1094 291 1108
rect 839 1094 871 1108
rect 1419 1094 1451 1108
rect 1999 1094 2031 1108
rect 2579 1094 2611 1108
rect 3159 1094 3191 1108
rect 3739 1094 3771 1108
rect 4319 1094 4351 1108
rect 4899 1094 4931 1108
rect 5479 1094 5511 1108
rect 6059 1094 6091 1108
rect 6639 1094 6671 1108
rect 73 1008 88 1036
rect 154 1008 169 1036
rect 381 1008 396 1036
rect 463 1008 478 1037
rect 653 1008 668 1036
rect 734 1008 749 1036
rect 961 1008 976 1036
rect 1043 1008 1058 1037
rect 1233 1008 1248 1036
rect 1314 1008 1329 1036
rect 1541 1008 1556 1036
rect 1623 1008 1638 1037
rect 1813 1008 1828 1036
rect 1894 1008 1909 1036
rect 2121 1008 2136 1036
rect 2203 1008 2218 1037
rect 2393 1008 2408 1036
rect 2474 1008 2489 1036
rect 2701 1008 2716 1036
rect 2783 1008 2798 1037
rect 2973 1008 2988 1036
rect 3054 1008 3069 1036
rect 3281 1008 3296 1036
rect 3363 1008 3378 1037
rect 3553 1008 3568 1036
rect 3634 1008 3649 1036
rect 3861 1008 3876 1036
rect 3943 1008 3958 1037
rect 4133 1008 4148 1036
rect 4214 1008 4229 1036
rect 4441 1008 4456 1036
rect 4523 1008 4538 1037
rect 4713 1007 4728 1035
rect 4794 1007 4809 1035
rect 5021 1007 5036 1035
rect 5103 1007 5118 1036
rect 5293 1007 5308 1035
rect 5374 1007 5389 1035
rect -1 862 14 904
rect 196 887 206 894
tri 206 887 213 894 sw
rect 196 862 213 887
rect 337 862 354 894
rect 536 862 551 904
rect 579 862 594 904
rect 776 887 786 894
tri 786 887 793 894 sw
rect 776 862 793 887
rect 917 862 934 894
rect 1116 862 1131 904
rect 1159 862 1174 904
rect 1356 887 1366 894
tri 1366 887 1373 894 sw
rect 1356 862 1373 887
rect 1497 862 1514 894
rect 1696 862 1711 904
rect 1739 862 1754 904
rect 1936 887 1946 894
tri 1946 887 1953 894 sw
rect 1936 862 1953 887
rect 2077 862 2094 894
rect 2276 862 2291 904
rect 2319 862 2334 904
rect 2516 887 2526 894
tri 2526 887 2533 894 sw
rect 2516 862 2533 887
rect 2657 862 2674 894
rect 2856 862 2871 904
rect 2899 862 2914 904
rect 3096 887 3106 894
tri 3106 887 3113 894 sw
rect 3096 862 3113 887
rect 3237 862 3254 894
rect 3436 862 3451 904
rect 3479 862 3494 904
rect 3676 887 3686 894
tri 3686 887 3693 894 sw
rect 3676 862 3693 887
rect 3817 862 3834 894
rect 4016 862 4031 904
rect 4059 862 4074 904
rect 4256 887 4266 894
tri 4266 887 4273 894 sw
rect 4256 862 4273 887
rect 4397 862 4414 894
rect 4596 862 4611 904
rect 5601 1007 5616 1035
rect 5683 1007 5698 1036
rect 5873 1007 5888 1035
rect 5954 1007 5969 1035
rect 6181 1007 6196 1035
rect 6263 1007 6278 1036
rect 6453 1007 6468 1035
rect 6534 1007 6549 1035
rect 6761 1007 6776 1035
rect 6843 1007 6858 1036
rect 259 824 291 838
rect 839 824 871 838
rect 1419 824 1451 838
rect 1999 824 2031 838
rect 2579 824 2611 838
rect 3159 824 3191 838
rect 3739 824 3771 838
rect 4639 861 4654 903
rect 4836 886 4846 893
tri 4846 886 4853 893 sw
rect 4836 861 4853 886
rect 4977 861 4994 893
rect 5176 861 5191 903
rect 5219 861 5234 903
rect 5416 886 5426 893
tri 5426 886 5433 893 sw
rect 5416 861 5433 886
rect 5557 861 5574 893
rect 5756 861 5771 903
rect 5799 861 5814 903
rect 5996 886 6006 893
tri 6006 886 6013 893 sw
rect 5996 861 6013 886
rect 6137 861 6154 893
rect 6336 861 6351 903
rect 6379 861 6394 903
rect 6576 886 6586 893
tri 6586 886 6593 893 sw
rect 6576 861 6593 886
rect 6717 861 6734 893
rect 6916 861 6931 903
rect 4319 824 4351 838
rect 4899 823 4931 837
rect 5479 823 5511 837
rect 6059 823 6091 837
rect 6639 823 6671 837
rect 73 738 88 766
rect 154 738 169 766
rect 381 738 396 766
rect 463 738 478 767
rect 653 738 668 766
rect 734 738 749 766
rect 961 738 976 766
rect 1043 738 1058 767
rect 1233 738 1248 766
rect 1314 738 1329 766
rect 1541 738 1556 766
rect 1623 738 1638 767
rect 1813 738 1828 766
rect 1894 738 1909 766
rect 2121 738 2136 766
rect 2203 738 2218 767
rect 2393 738 2408 766
rect 2474 738 2489 766
rect 2701 738 2716 766
rect 2783 738 2798 767
rect 2973 738 2988 766
rect 3054 738 3069 766
rect 3281 738 3296 766
rect 3363 738 3378 767
rect 3553 738 3568 766
rect 3634 738 3649 766
rect 3861 738 3876 766
rect 3943 738 3958 767
rect 4133 738 4148 766
rect 4214 738 4229 766
rect 4441 738 4456 766
rect 4523 738 4538 767
rect 4713 737 4728 765
rect 4794 737 4809 765
rect 5021 737 5036 765
rect 5103 737 5118 766
rect 5293 737 5308 765
rect 5374 737 5389 765
rect -1 592 14 634
rect 196 617 206 624
tri 206 617 213 624 sw
rect 196 592 213 617
rect 337 592 354 624
rect 536 592 551 634
rect 579 592 594 634
rect 776 617 786 624
tri 786 617 793 624 sw
rect 776 592 793 617
rect 917 592 934 624
rect 1116 592 1131 634
rect 1159 592 1174 634
rect 1356 617 1366 624
tri 1366 617 1373 624 sw
rect 1356 592 1373 617
rect 1497 592 1514 624
rect 1696 592 1711 634
rect 1739 592 1754 634
rect 1936 617 1946 624
tri 1946 617 1953 624 sw
rect 1936 592 1953 617
rect 2077 592 2094 624
rect 2276 592 2291 634
rect 2319 592 2334 634
rect 2516 617 2526 624
tri 2526 617 2533 624 sw
rect 2516 592 2533 617
rect 2657 592 2674 624
rect 2856 592 2871 634
rect 2899 592 2914 634
rect 3096 617 3106 624
tri 3106 617 3113 624 sw
rect 3096 592 3113 617
rect 3237 592 3254 624
rect 3436 592 3451 634
rect 3479 592 3494 634
rect 3676 617 3686 624
tri 3686 617 3693 624 sw
rect 3676 592 3693 617
rect 3817 592 3834 624
rect 4016 592 4031 634
rect 4059 592 4074 634
rect 4256 617 4266 624
tri 4266 617 4273 624 sw
rect 4256 592 4273 617
rect 4397 592 4414 624
rect 4596 592 4611 634
rect 5601 737 5616 765
rect 5683 737 5698 766
rect 5873 737 5888 765
rect 5954 737 5969 765
rect 6181 737 6196 765
rect 6263 737 6278 766
rect 6453 737 6468 765
rect 6534 737 6549 765
rect 6761 737 6776 765
rect 6843 737 6858 766
rect 259 554 291 568
rect 839 554 871 568
rect 1419 554 1451 568
rect 1999 554 2031 568
rect 2579 554 2611 568
rect 3159 554 3191 568
rect 3739 554 3771 568
rect 4639 591 4654 633
rect 4836 616 4846 623
tri 4846 616 4853 623 sw
rect 4836 591 4853 616
rect 4977 591 4994 623
rect 5176 591 5191 633
rect 5219 591 5234 633
rect 5416 616 5426 623
tri 5426 616 5433 623 sw
rect 5416 591 5433 616
rect 5557 591 5574 623
rect 5756 591 5771 633
rect 5799 591 5814 633
rect 5996 616 6006 623
tri 6006 616 6013 623 sw
rect 5996 591 6013 616
rect 6137 591 6154 623
rect 6336 591 6351 633
rect 6379 591 6394 633
rect 6576 616 6586 623
tri 6586 616 6593 623 sw
rect 6576 591 6593 616
rect 6717 591 6734 623
rect 6916 591 6931 633
rect 4319 554 4351 568
rect 4899 553 4931 567
rect 5479 553 5511 567
rect 6059 553 6091 567
rect 6639 553 6671 567
rect 73 468 88 496
rect 154 468 169 496
rect 381 468 396 496
rect 463 468 478 497
rect 653 468 668 496
rect 734 468 749 496
rect 961 468 976 496
rect 1043 468 1058 497
rect 1233 468 1248 496
rect 1314 468 1329 496
rect 1541 468 1556 496
rect 1623 468 1638 497
rect 1813 468 1828 496
rect 1894 468 1909 496
rect 2121 468 2136 496
rect 2203 468 2218 497
rect 2393 468 2408 496
rect 2474 468 2489 496
rect 2701 468 2716 496
rect 2783 468 2798 497
rect 2973 468 2988 496
rect 3054 468 3069 496
rect 3281 468 3296 496
rect 3363 468 3378 497
rect 3553 468 3568 496
rect 3634 468 3649 496
rect 3861 468 3876 496
rect 3943 468 3958 497
rect 4133 468 4148 496
rect 4214 468 4229 496
rect 4441 468 4456 496
rect 4523 468 4538 497
rect 4713 467 4728 495
rect 4794 467 4809 495
rect 5021 467 5036 495
rect 5103 467 5118 496
rect 5293 467 5308 495
rect 5374 467 5389 495
rect -1 322 14 364
rect 196 347 206 354
tri 206 347 213 354 sw
rect 196 322 213 347
rect 337 322 354 354
rect 536 322 551 364
rect 579 322 594 364
rect 776 347 786 354
tri 786 347 793 354 sw
rect 776 322 793 347
rect 917 322 934 354
rect 1116 322 1131 364
rect 1159 322 1174 364
rect 1356 347 1366 354
tri 1366 347 1373 354 sw
rect 1356 322 1373 347
rect 1497 322 1514 354
rect 1696 322 1711 364
rect 1739 322 1754 364
rect 1936 347 1946 354
tri 1946 347 1953 354 sw
rect 1936 322 1953 347
rect 2077 322 2094 354
rect 2276 322 2291 364
rect 2319 322 2334 364
rect 2516 347 2526 354
tri 2526 347 2533 354 sw
rect 2516 322 2533 347
rect 2657 322 2674 354
rect 2856 322 2871 364
rect 2899 322 2914 364
rect 3096 347 3106 354
tri 3106 347 3113 354 sw
rect 3096 322 3113 347
rect 3237 322 3254 354
rect 3436 322 3451 364
rect 3479 322 3494 364
rect 3676 347 3686 354
tri 3686 347 3693 354 sw
rect 3676 322 3693 347
rect 3817 322 3834 354
rect 4016 322 4031 364
rect 4059 322 4074 364
rect 4256 347 4266 354
tri 4266 347 4273 354 sw
rect 4256 322 4273 347
rect 4397 322 4414 354
rect 4596 322 4611 364
rect 5601 467 5616 495
rect 5683 467 5698 496
rect 5873 467 5888 495
rect 5954 467 5969 495
rect 6181 467 6196 495
rect 6263 467 6278 496
rect 6453 467 6468 495
rect 6534 467 6549 495
rect 6761 467 6776 495
rect 6843 467 6858 496
rect 259 284 291 298
rect 839 284 871 298
rect 1419 284 1451 298
rect 1999 284 2031 298
rect 2579 284 2611 298
rect 3159 284 3191 298
rect 3739 284 3771 298
rect 4639 321 4654 363
rect 4836 346 4846 353
tri 4846 346 4853 353 sw
rect 4836 321 4853 346
rect 4977 321 4994 353
rect 5176 321 5191 363
rect 5219 321 5234 363
rect 5416 346 5426 353
tri 5426 346 5433 353 sw
rect 5416 321 5433 346
rect 5557 321 5574 353
rect 5756 321 5771 363
rect 5799 321 5814 363
rect 5996 346 6006 353
tri 6006 346 6013 353 sw
rect 5996 321 6013 346
rect 6137 321 6154 353
rect 6336 321 6351 363
rect 6379 321 6394 363
rect 6576 346 6586 353
tri 6586 346 6593 353 sw
rect 6576 321 6593 346
rect 6717 321 6734 353
rect 6916 321 6931 363
rect 4319 284 4351 298
rect 4899 283 4931 297
rect 5479 283 5511 297
rect 6059 283 6091 297
rect 6639 283 6671 297
rect 73 198 88 226
rect 154 198 169 226
rect 381 198 396 226
rect 463 198 478 227
rect 653 198 668 226
rect 734 198 749 226
rect 961 198 976 226
rect 1043 198 1058 227
rect 1233 198 1248 226
rect 1314 198 1329 226
rect 1541 198 1556 226
rect 1623 198 1638 227
rect 1813 198 1828 226
rect 1894 198 1909 226
rect 2121 198 2136 226
rect 2203 198 2218 227
rect 2393 198 2408 226
rect 2474 198 2489 226
rect 2701 198 2716 226
rect 2783 198 2798 227
rect 2973 198 2988 226
rect 3054 198 3069 226
rect 3281 198 3296 226
rect 3363 198 3378 227
rect 3553 198 3568 226
rect 3634 198 3649 226
rect 3861 198 3876 226
rect 3943 198 3958 227
rect 4133 198 4148 226
rect 4214 198 4229 226
rect 4441 198 4456 226
rect 4523 198 4538 227
rect 4713 197 4728 225
rect 4794 197 4809 225
rect 5021 197 5036 225
rect 5103 197 5118 226
rect 5293 197 5308 225
rect 5374 197 5389 225
rect -1 52 14 94
rect 196 77 206 84
tri 206 77 213 84 sw
rect 196 52 213 77
rect 337 52 354 84
rect 536 52 551 94
rect 579 52 594 94
rect 776 77 786 84
tri 786 77 793 84 sw
rect 776 52 793 77
rect 917 52 934 84
rect 1116 52 1131 94
rect 1159 52 1174 94
rect 1356 77 1366 84
tri 1366 77 1373 84 sw
rect 1356 52 1373 77
rect 1497 52 1514 84
rect 1696 52 1711 94
rect 1739 52 1754 94
rect 1936 77 1946 84
tri 1946 77 1953 84 sw
rect 1936 52 1953 77
rect 2077 52 2094 84
rect 2276 52 2291 94
rect 2319 52 2334 94
rect 2516 77 2526 84
tri 2526 77 2533 84 sw
rect 2516 52 2533 77
rect 2657 52 2674 84
rect 2856 52 2871 94
rect 2899 52 2914 94
rect 3096 77 3106 84
tri 3106 77 3113 84 sw
rect 3096 52 3113 77
rect 3237 52 3254 84
rect 3436 52 3451 94
rect 3479 52 3494 94
rect 3676 77 3686 84
tri 3686 77 3693 84 sw
rect 3676 52 3693 77
rect 3817 52 3834 84
rect 4016 52 4031 94
rect 4059 52 4074 94
rect 4256 77 4266 84
tri 4266 77 4273 84 sw
rect 4256 52 4273 77
rect 4397 52 4414 84
rect 4596 52 4611 94
rect 5601 197 5616 225
rect 5683 197 5698 226
rect 5873 197 5888 225
rect 5954 197 5969 225
rect 6181 197 6196 225
rect 6263 197 6278 226
rect 6453 197 6468 225
rect 6534 197 6549 225
rect 6761 197 6776 225
rect 6843 197 6858 226
rect 259 14 291 28
rect 839 14 871 28
rect 1419 14 1451 28
rect 1999 14 2031 28
rect 2579 14 2611 28
rect 3159 14 3191 28
rect 3739 14 3771 28
rect 4639 51 4654 93
rect 4836 76 4846 83
tri 4846 76 4853 83 sw
rect 4836 51 4853 76
rect 4977 51 4994 83
rect 5176 51 5191 93
rect 5219 51 5234 93
rect 5416 76 5426 83
tri 5426 76 5433 83 sw
rect 5416 51 5433 76
rect 5557 51 5574 83
rect 5756 51 5771 93
rect 5799 51 5814 93
rect 5996 76 6006 83
tri 6006 76 6013 83 sw
rect 5996 51 6013 76
rect 6137 51 6154 83
rect 6336 51 6351 93
rect 6379 51 6394 93
rect 6576 76 6586 83
tri 6586 76 6593 83 sw
rect 6576 51 6593 76
rect 6717 51 6734 83
rect 6916 51 6931 93
rect 4319 14 4351 28
rect 4899 13 4931 27
rect 5479 13 5511 27
rect 6059 13 6091 27
rect 6639 13 6671 27
rect 73 -72 88 -44
rect 154 -72 169 -44
rect 381 -72 396 -44
rect 463 -72 478 -43
rect 653 -72 668 -44
rect 734 -72 749 -44
rect 961 -72 976 -44
rect 1043 -72 1058 -43
rect 1233 -72 1248 -44
rect 1314 -72 1329 -44
rect 1541 -72 1556 -44
rect 1623 -72 1638 -43
rect 1813 -72 1828 -44
rect 1894 -72 1909 -44
rect 2121 -72 2136 -44
rect 2203 -72 2218 -43
rect 2393 -72 2408 -44
rect 2474 -72 2489 -44
rect 2701 -72 2716 -44
rect 2783 -72 2798 -43
rect 2973 -72 2988 -44
rect 3054 -72 3069 -44
rect 3281 -72 3296 -44
rect 3363 -72 3378 -43
rect 3553 -72 3568 -44
rect 3634 -72 3649 -44
rect 3861 -72 3876 -44
rect 3943 -72 3958 -43
rect 4133 -72 4148 -44
rect 4214 -72 4229 -44
rect 4441 -72 4456 -44
rect 4523 -72 4538 -43
rect 4713 -73 4728 -45
rect 4794 -73 4809 -45
rect 5021 -73 5036 -45
rect 5103 -73 5118 -44
rect 5293 -73 5308 -45
rect 5374 -73 5389 -45
rect -1 -218 14 -176
rect 196 -193 206 -186
tri 206 -193 213 -186 sw
rect 196 -218 213 -193
rect 337 -218 354 -186
rect 536 -218 551 -176
rect 579 -218 594 -176
rect 776 -193 786 -186
tri 786 -193 793 -186 sw
rect 776 -218 793 -193
rect 917 -218 934 -186
rect 1116 -218 1131 -176
rect 1159 -218 1174 -176
rect 1356 -193 1366 -186
tri 1366 -193 1373 -186 sw
rect 1356 -218 1373 -193
rect 1497 -218 1514 -186
rect 1696 -218 1711 -176
rect 1739 -218 1754 -176
rect 1936 -193 1946 -186
tri 1946 -193 1953 -186 sw
rect 1936 -218 1953 -193
rect 2077 -218 2094 -186
rect 2276 -218 2291 -176
rect 2319 -218 2334 -176
rect 2516 -193 2526 -186
tri 2526 -193 2533 -186 sw
rect 2516 -218 2533 -193
rect 2657 -218 2674 -186
rect 2856 -218 2871 -176
rect 2899 -218 2914 -176
rect 3096 -193 3106 -186
tri 3106 -193 3113 -186 sw
rect 3096 -218 3113 -193
rect 3237 -218 3254 -186
rect 3436 -218 3451 -176
rect 3479 -218 3494 -176
rect 3676 -193 3686 -186
tri 3686 -193 3693 -186 sw
rect 3676 -218 3693 -193
rect 3817 -218 3834 -186
rect 4016 -218 4031 -176
rect 4059 -218 4074 -176
rect 4256 -193 4266 -186
tri 4266 -193 4273 -186 sw
rect 4256 -218 4273 -193
rect 4397 -218 4414 -186
rect 4596 -218 4611 -176
rect 5601 -73 5616 -45
rect 5683 -73 5698 -44
rect 5873 -73 5888 -45
rect 5954 -73 5969 -45
rect 6181 -73 6196 -45
rect 6263 -73 6278 -44
rect 6453 -73 6468 -45
rect 6534 -73 6549 -45
rect 6761 -73 6776 -45
rect 6843 -73 6858 -44
rect 259 -256 291 -242
rect 839 -256 871 -242
rect 1419 -256 1451 -242
rect 1999 -256 2031 -242
rect 2579 -256 2611 -242
rect 3159 -256 3191 -242
rect 3739 -256 3771 -242
rect 4639 -219 4654 -177
rect 4836 -194 4846 -187
tri 4846 -194 4853 -187 sw
rect 4836 -219 4853 -194
rect 4977 -219 4994 -187
rect 5176 -219 5191 -177
rect 5219 -219 5234 -177
rect 5416 -194 5426 -187
tri 5426 -194 5433 -187 sw
rect 5416 -219 5433 -194
rect 5557 -219 5574 -187
rect 5756 -219 5771 -177
rect 5799 -219 5814 -177
rect 5996 -194 6006 -187
tri 6006 -194 6013 -187 sw
rect 5996 -219 6013 -194
rect 6137 -219 6154 -187
rect 6336 -219 6351 -177
rect 6379 -219 6394 -177
rect 6576 -194 6586 -187
tri 6586 -194 6593 -187 sw
rect 6576 -219 6593 -194
rect 6717 -219 6734 -187
rect 6916 -219 6931 -177
rect 4319 -256 4351 -242
rect 4899 -257 4931 -243
rect 5479 -257 5511 -243
rect 6059 -257 6091 -243
rect 6639 -257 6671 -243
rect 73 -342 88 -314
rect 154 -342 169 -314
rect 381 -342 396 -314
rect 463 -342 478 -313
rect 653 -342 668 -314
rect 734 -342 749 -314
rect 961 -342 976 -314
rect 1043 -342 1058 -313
rect 1233 -342 1248 -314
rect 1314 -342 1329 -314
rect 1541 -342 1556 -314
rect 1623 -342 1638 -313
rect 1813 -342 1828 -314
rect 1894 -342 1909 -314
rect 2121 -342 2136 -314
rect 2203 -342 2218 -313
rect 2393 -342 2408 -314
rect 2474 -342 2489 -314
rect 2701 -342 2716 -314
rect 2783 -342 2798 -313
rect 2973 -342 2988 -314
rect 3054 -342 3069 -314
rect 3281 -342 3296 -314
rect 3363 -342 3378 -313
rect 3553 -342 3568 -314
rect 3634 -342 3649 -314
rect 3861 -342 3876 -314
rect 3943 -342 3958 -313
rect 4133 -342 4148 -314
rect 4214 -342 4229 -314
rect 4441 -342 4456 -314
rect 4523 -342 4538 -313
rect 4713 -343 4728 -315
rect 4794 -343 4809 -315
rect 5021 -343 5036 -315
rect 5103 -343 5118 -314
rect 5293 -343 5308 -315
rect 5374 -343 5389 -315
rect -1 -488 14 -446
rect 196 -463 206 -456
tri 206 -463 213 -456 sw
rect 196 -488 213 -463
rect 337 -488 354 -456
rect 536 -488 551 -446
rect 579 -488 594 -446
rect 776 -463 786 -456
tri 786 -463 793 -456 sw
rect 776 -488 793 -463
rect 917 -488 934 -456
rect 1116 -488 1131 -446
rect 1159 -488 1174 -446
rect 1356 -463 1366 -456
tri 1366 -463 1373 -456 sw
rect 1356 -488 1373 -463
rect 1497 -488 1514 -456
rect 1696 -488 1711 -446
rect 1739 -488 1754 -446
rect 1936 -463 1946 -456
tri 1946 -463 1953 -456 sw
rect 1936 -488 1953 -463
rect 2077 -488 2094 -456
rect 2276 -488 2291 -446
rect 2319 -488 2334 -446
rect 2516 -463 2526 -456
tri 2526 -463 2533 -456 sw
rect 2516 -488 2533 -463
rect 2657 -488 2674 -456
rect 2856 -488 2871 -446
rect 2899 -488 2914 -446
rect 3096 -463 3106 -456
tri 3106 -463 3113 -456 sw
rect 3096 -488 3113 -463
rect 3237 -488 3254 -456
rect 3436 -488 3451 -446
rect 3479 -488 3494 -446
rect 3676 -463 3686 -456
tri 3686 -463 3693 -456 sw
rect 3676 -488 3693 -463
rect 3817 -488 3834 -456
rect 4016 -488 4031 -446
rect 4059 -488 4074 -446
rect 4256 -463 4266 -456
tri 4266 -463 4273 -456 sw
rect 4256 -488 4273 -463
rect 4397 -488 4414 -456
rect 4596 -488 4611 -446
rect 5601 -343 5616 -315
rect 5683 -343 5698 -314
rect 5873 -343 5888 -315
rect 5954 -343 5969 -315
rect 6181 -343 6196 -315
rect 6263 -343 6278 -314
rect 6453 -343 6468 -315
rect 6534 -343 6549 -315
rect 6761 -343 6776 -315
rect 6843 -343 6858 -314
rect 259 -526 291 -512
rect 839 -526 871 -512
rect 1419 -526 1451 -512
rect 1999 -526 2031 -512
rect 2579 -526 2611 -512
rect 3159 -526 3191 -512
rect 3739 -526 3771 -512
rect 4639 -489 4654 -447
rect 4836 -464 4846 -457
tri 4846 -464 4853 -457 sw
rect 4836 -489 4853 -464
rect 4977 -489 4994 -457
rect 5176 -489 5191 -447
rect 5219 -489 5234 -447
rect 5416 -464 5426 -457
tri 5426 -464 5433 -457 sw
rect 5416 -489 5433 -464
rect 5557 -489 5574 -457
rect 5756 -489 5771 -447
rect 5799 -489 5814 -447
rect 5996 -464 6006 -457
tri 6006 -464 6013 -457 sw
rect 5996 -489 6013 -464
rect 6137 -489 6154 -457
rect 6336 -489 6351 -447
rect 6379 -489 6394 -447
rect 6576 -464 6586 -457
tri 6586 -464 6593 -457 sw
rect 6576 -489 6593 -464
rect 6717 -489 6734 -457
rect 6916 -489 6931 -447
rect 4319 -526 4351 -512
rect 4899 -527 4931 -513
rect 5479 -527 5511 -513
rect 6059 -527 6091 -513
rect 6639 -527 6671 -513
rect 73 -612 88 -584
rect 154 -612 169 -584
rect 381 -612 396 -584
rect 463 -612 478 -583
rect 653 -612 668 -584
rect 734 -612 749 -584
rect 961 -612 976 -584
rect 1043 -612 1058 -583
rect 1233 -612 1248 -584
rect 1314 -612 1329 -584
rect 1541 -612 1556 -584
rect 1623 -612 1638 -583
rect 1813 -612 1828 -584
rect 1894 -612 1909 -584
rect 2121 -612 2136 -584
rect 2203 -612 2218 -583
rect 2393 -612 2408 -584
rect 2474 -612 2489 -584
rect 2701 -612 2716 -584
rect 2783 -612 2798 -583
rect 2973 -612 2988 -584
rect 3054 -612 3069 -584
rect 3281 -612 3296 -584
rect 3363 -612 3378 -583
rect 3553 -612 3568 -584
rect 3634 -612 3649 -584
rect 3861 -612 3876 -584
rect 3943 -612 3958 -583
rect 4133 -612 4148 -584
rect 4214 -612 4229 -584
rect 4441 -612 4456 -584
rect 4523 -612 4538 -583
rect 4713 -613 4728 -585
rect 4794 -613 4809 -585
rect 5021 -613 5036 -585
rect 5103 -613 5118 -584
rect 5293 -613 5308 -585
rect 5374 -613 5389 -585
rect -1 -758 14 -716
rect 196 -733 206 -726
tri 206 -733 213 -726 sw
rect 196 -758 213 -733
rect 337 -758 354 -726
rect 536 -758 551 -716
rect 579 -758 594 -716
rect 776 -733 786 -726
tri 786 -733 793 -726 sw
rect 776 -758 793 -733
rect 917 -758 934 -726
rect 1116 -758 1131 -716
rect 1159 -758 1174 -716
rect 1356 -733 1366 -726
tri 1366 -733 1373 -726 sw
rect 1356 -758 1373 -733
rect 1497 -758 1514 -726
rect 1696 -758 1711 -716
rect 1739 -758 1754 -716
rect 1936 -733 1946 -726
tri 1946 -733 1953 -726 sw
rect 1936 -758 1953 -733
rect 2077 -758 2094 -726
rect 2276 -758 2291 -716
rect 2319 -758 2334 -716
rect 2516 -733 2526 -726
tri 2526 -733 2533 -726 sw
rect 2516 -758 2533 -733
rect 2657 -758 2674 -726
rect 2856 -758 2871 -716
rect 2899 -758 2914 -716
rect 3096 -733 3106 -726
tri 3106 -733 3113 -726 sw
rect 3096 -758 3113 -733
rect 3237 -758 3254 -726
rect 3436 -758 3451 -716
rect 3479 -758 3494 -716
rect 3676 -733 3686 -726
tri 3686 -733 3693 -726 sw
rect 3676 -758 3693 -733
rect 3817 -758 3834 -726
rect 4016 -758 4031 -716
rect 4059 -758 4074 -716
rect 4256 -733 4266 -726
tri 4266 -733 4273 -726 sw
rect 4256 -758 4273 -733
rect 4397 -758 4414 -726
rect 4596 -758 4611 -716
rect 5601 -613 5616 -585
rect 5683 -613 5698 -584
rect 5873 -613 5888 -585
rect 5954 -613 5969 -585
rect 6181 -613 6196 -585
rect 6263 -613 6278 -584
rect 6453 -613 6468 -585
rect 6534 -613 6549 -585
rect 6761 -613 6776 -585
rect 6843 -613 6858 -584
rect 259 -796 291 -782
rect 839 -796 871 -782
rect 1419 -796 1451 -782
rect 1999 -796 2031 -782
rect 2579 -796 2611 -782
rect 3159 -796 3191 -782
rect 3739 -796 3771 -782
rect 4639 -759 4654 -717
rect 4836 -734 4846 -727
tri 4846 -734 4853 -727 sw
rect 4836 -759 4853 -734
rect 4977 -759 4994 -727
rect 5176 -759 5191 -717
rect 5219 -759 5234 -717
rect 5416 -734 5426 -727
tri 5426 -734 5433 -727 sw
rect 5416 -759 5433 -734
rect 5557 -759 5574 -727
rect 5756 -759 5771 -717
rect 5799 -759 5814 -717
rect 5996 -734 6006 -727
tri 6006 -734 6013 -727 sw
rect 5996 -759 6013 -734
rect 6137 -759 6154 -727
rect 6336 -759 6351 -717
rect 6379 -759 6394 -717
rect 6576 -734 6586 -727
tri 6586 -734 6593 -727 sw
rect 6576 -759 6593 -734
rect 6717 -759 6734 -727
rect 6916 -759 6931 -717
rect 4319 -796 4351 -782
rect 4899 -797 4931 -783
rect 5479 -797 5511 -783
rect 6059 -797 6091 -783
rect 6639 -797 6671 -783
rect 73 -882 88 -854
rect 154 -882 169 -854
rect 381 -882 396 -854
rect 463 -882 478 -853
rect 653 -882 668 -854
rect 734 -882 749 -854
rect 961 -882 976 -854
rect 1043 -882 1058 -853
rect 1233 -882 1248 -854
rect 1314 -882 1329 -854
rect 1541 -882 1556 -854
rect 1623 -882 1638 -853
rect 1813 -882 1828 -854
rect 1894 -882 1909 -854
rect 2121 -882 2136 -854
rect 2203 -882 2218 -853
rect 2393 -882 2408 -854
rect 2474 -882 2489 -854
rect 2701 -882 2716 -854
rect 2783 -882 2798 -853
rect 2973 -882 2988 -854
rect 3054 -882 3069 -854
rect 3281 -882 3296 -854
rect 3363 -882 3378 -853
rect 3553 -882 3568 -854
rect 3634 -882 3649 -854
rect 3861 -882 3876 -854
rect 3943 -882 3958 -853
rect 4133 -882 4148 -854
rect 4214 -882 4229 -854
rect 4441 -882 4456 -854
rect 4523 -882 4538 -853
rect 4713 -883 4728 -855
rect 4794 -883 4809 -855
rect 5021 -883 5036 -855
rect 5103 -883 5118 -854
rect 5293 -883 5308 -855
rect 5374 -883 5389 -855
rect -1 -1028 14 -986
rect 196 -1003 206 -996
tri 206 -1003 213 -996 sw
rect 196 -1028 213 -1003
rect 337 -1028 354 -996
rect 536 -1028 551 -986
rect 579 -1028 594 -986
rect 776 -1003 786 -996
tri 786 -1003 793 -996 sw
rect 776 -1028 793 -1003
rect 917 -1028 934 -996
rect 1116 -1028 1131 -986
rect 1159 -1028 1174 -986
rect 1356 -1003 1366 -996
tri 1366 -1003 1373 -996 sw
rect 1356 -1028 1373 -1003
rect 1497 -1028 1514 -996
rect 1696 -1028 1711 -986
rect 1739 -1028 1754 -986
rect 1936 -1003 1946 -996
tri 1946 -1003 1953 -996 sw
rect 1936 -1028 1953 -1003
rect 2077 -1028 2094 -996
rect 2276 -1028 2291 -986
rect 2319 -1028 2334 -986
rect 2516 -1003 2526 -996
tri 2526 -1003 2533 -996 sw
rect 2516 -1028 2533 -1003
rect 2657 -1028 2674 -996
rect 2856 -1028 2871 -986
rect 2899 -1028 2914 -986
rect 3096 -1003 3106 -996
tri 3106 -1003 3113 -996 sw
rect 3096 -1028 3113 -1003
rect 3237 -1028 3254 -996
rect 3436 -1028 3451 -986
rect 3479 -1028 3494 -986
rect 3676 -1003 3686 -996
tri 3686 -1003 3693 -996 sw
rect 3676 -1028 3693 -1003
rect 3817 -1028 3834 -996
rect 4016 -1028 4031 -986
rect 4059 -1028 4074 -986
rect 4256 -1003 4266 -996
tri 4266 -1003 4273 -996 sw
rect 4256 -1028 4273 -1003
rect 4397 -1028 4414 -996
rect 4596 -1028 4611 -986
rect 5601 -883 5616 -855
rect 5683 -883 5698 -854
rect 5873 -883 5888 -855
rect 5954 -883 5969 -855
rect 6181 -883 6196 -855
rect 6263 -883 6278 -854
rect 6453 -883 6468 -855
rect 6534 -883 6549 -855
rect 6761 -883 6776 -855
rect 6843 -883 6858 -854
rect 259 -1066 291 -1052
rect 839 -1066 871 -1052
rect 1419 -1066 1451 -1052
rect 1999 -1066 2031 -1052
rect 2579 -1066 2611 -1052
rect 3159 -1066 3191 -1052
rect 3739 -1066 3771 -1052
rect 4639 -1029 4654 -987
rect 4836 -1004 4846 -997
tri 4846 -1004 4853 -997 sw
rect 4836 -1029 4853 -1004
rect 4977 -1029 4994 -997
rect 5176 -1029 5191 -987
rect 5219 -1029 5234 -987
rect 5416 -1004 5426 -997
tri 5426 -1004 5433 -997 sw
rect 5416 -1029 5433 -1004
rect 5557 -1029 5574 -997
rect 5756 -1029 5771 -987
rect 5799 -1029 5814 -987
rect 5996 -1004 6006 -997
tri 6006 -1004 6013 -997 sw
rect 5996 -1029 6013 -1004
rect 6137 -1029 6154 -997
rect 6336 -1029 6351 -987
rect 6379 -1029 6394 -987
rect 6576 -1004 6586 -997
tri 6586 -1004 6593 -997 sw
rect 6576 -1029 6593 -1004
rect 6717 -1029 6734 -997
rect 6916 -1029 6931 -987
rect 4319 -1066 4351 -1052
rect 4899 -1067 4931 -1053
rect 5479 -1067 5511 -1053
rect 6059 -1067 6091 -1053
rect 6639 -1067 6671 -1053
rect 73 -1152 88 -1124
rect 154 -1152 169 -1124
rect 381 -1152 396 -1124
rect 463 -1152 478 -1123
rect 653 -1152 668 -1124
rect 734 -1152 749 -1124
rect 961 -1152 976 -1124
rect 1043 -1152 1058 -1123
rect 1233 -1152 1248 -1124
rect 1314 -1152 1329 -1124
rect 1541 -1152 1556 -1124
rect 1623 -1152 1638 -1123
rect 1813 -1152 1828 -1124
rect 1894 -1152 1909 -1124
rect 2121 -1152 2136 -1124
rect 2203 -1152 2218 -1123
rect 2393 -1152 2408 -1124
rect 2474 -1152 2489 -1124
rect 2701 -1152 2716 -1124
rect 2783 -1152 2798 -1123
rect 2973 -1152 2988 -1124
rect 3054 -1152 3069 -1124
rect 3281 -1152 3296 -1124
rect 3363 -1152 3378 -1123
rect 3553 -1152 3568 -1124
rect 3634 -1152 3649 -1124
rect 3861 -1152 3876 -1124
rect 3943 -1152 3958 -1123
rect 4133 -1152 4148 -1124
rect 4214 -1152 4229 -1124
rect 4441 -1152 4456 -1124
rect 4523 -1152 4538 -1123
rect 4713 -1153 4728 -1125
rect 4794 -1153 4809 -1125
rect 5021 -1153 5036 -1125
rect 5103 -1153 5118 -1124
rect 5293 -1153 5308 -1125
rect 5374 -1153 5389 -1125
rect -1 -1298 14 -1256
rect 196 -1273 206 -1266
tri 206 -1273 213 -1266 sw
rect 196 -1298 213 -1273
rect 337 -1298 354 -1266
rect 536 -1298 551 -1256
rect 579 -1298 594 -1256
rect 776 -1273 786 -1266
tri 786 -1273 793 -1266 sw
rect 776 -1298 793 -1273
rect 917 -1298 934 -1266
rect 1116 -1298 1131 -1256
rect 1159 -1298 1174 -1256
rect 1356 -1273 1366 -1266
tri 1366 -1273 1373 -1266 sw
rect 1356 -1298 1373 -1273
rect 1497 -1298 1514 -1266
rect 1696 -1298 1711 -1256
rect 1739 -1298 1754 -1256
rect 1936 -1273 1946 -1266
tri 1946 -1273 1953 -1266 sw
rect 1936 -1298 1953 -1273
rect 2077 -1298 2094 -1266
rect 2276 -1298 2291 -1256
rect 2319 -1298 2334 -1256
rect 2516 -1273 2526 -1266
tri 2526 -1273 2533 -1266 sw
rect 2516 -1298 2533 -1273
rect 2657 -1298 2674 -1266
rect 2856 -1298 2871 -1256
rect 2899 -1298 2914 -1256
rect 3096 -1273 3106 -1266
tri 3106 -1273 3113 -1266 sw
rect 3096 -1298 3113 -1273
rect 3237 -1298 3254 -1266
rect 3436 -1298 3451 -1256
rect 3479 -1298 3494 -1256
rect 3676 -1273 3686 -1266
tri 3686 -1273 3693 -1266 sw
rect 3676 -1298 3693 -1273
rect 3817 -1298 3834 -1266
rect 4016 -1298 4031 -1256
rect 4059 -1298 4074 -1256
rect 4256 -1273 4266 -1266
tri 4266 -1273 4273 -1266 sw
rect 4256 -1298 4273 -1273
rect 4397 -1298 4414 -1266
rect 4596 -1298 4611 -1256
rect 5601 -1153 5616 -1125
rect 5683 -1153 5698 -1124
rect 5873 -1153 5888 -1125
rect 5954 -1153 5969 -1125
rect 6181 -1153 6196 -1125
rect 6263 -1153 6278 -1124
rect 6453 -1153 6468 -1125
rect 6534 -1153 6549 -1125
rect 6761 -1153 6776 -1125
rect 6843 -1153 6858 -1124
rect 259 -1336 291 -1322
rect 839 -1336 871 -1322
rect 1419 -1336 1451 -1322
rect 1999 -1336 2031 -1322
rect 2579 -1336 2611 -1322
rect 3159 -1336 3191 -1322
rect 3739 -1336 3771 -1322
rect 4639 -1299 4654 -1257
rect 4836 -1274 4846 -1267
tri 4846 -1274 4853 -1267 sw
rect 4836 -1299 4853 -1274
rect 4977 -1299 4994 -1267
rect 5176 -1299 5191 -1257
rect 5219 -1299 5234 -1257
rect 5416 -1274 5426 -1267
tri 5426 -1274 5433 -1267 sw
rect 5416 -1299 5433 -1274
rect 5557 -1299 5574 -1267
rect 5756 -1299 5771 -1257
rect 5799 -1299 5814 -1257
rect 5996 -1274 6006 -1267
tri 6006 -1274 6013 -1267 sw
rect 5996 -1299 6013 -1274
rect 6137 -1299 6154 -1267
rect 6336 -1299 6351 -1257
rect 6379 -1299 6394 -1257
rect 6576 -1274 6586 -1267
tri 6586 -1274 6593 -1267 sw
rect 6576 -1299 6593 -1274
rect 6717 -1299 6734 -1267
rect 6916 -1299 6931 -1257
rect 4319 -1336 4351 -1322
rect 4899 -1337 4931 -1323
rect 5479 -1337 5511 -1323
rect 6059 -1337 6091 -1323
rect 6639 -1337 6671 -1323
rect 73 -1422 88 -1394
rect 154 -1422 169 -1394
rect 381 -1422 396 -1394
rect 463 -1422 478 -1393
rect 653 -1422 668 -1394
rect 734 -1422 749 -1394
rect 961 -1422 976 -1394
rect 1043 -1422 1058 -1393
rect 1233 -1422 1248 -1394
rect 1314 -1422 1329 -1394
rect 1541 -1422 1556 -1394
rect 1623 -1422 1638 -1393
rect 1813 -1422 1828 -1394
rect 1894 -1422 1909 -1394
rect 2121 -1422 2136 -1394
rect 2203 -1422 2218 -1393
rect 2393 -1422 2408 -1394
rect 2474 -1422 2489 -1394
rect 2701 -1422 2716 -1394
rect 2783 -1422 2798 -1393
rect 2973 -1422 2988 -1394
rect 3054 -1422 3069 -1394
rect 3281 -1422 3296 -1394
rect 3363 -1422 3378 -1393
rect 3553 -1422 3568 -1394
rect 3634 -1422 3649 -1394
rect 3861 -1422 3876 -1394
rect 3943 -1422 3958 -1393
rect 4133 -1422 4148 -1394
rect 4214 -1422 4229 -1394
rect 4441 -1422 4456 -1394
rect 4523 -1422 4538 -1393
rect 4713 -1423 4728 -1395
rect 4794 -1423 4809 -1395
rect 5021 -1423 5036 -1395
rect 5103 -1423 5118 -1394
rect 5293 -1423 5308 -1395
rect 5374 -1423 5389 -1395
rect -1 -1568 14 -1526
rect 196 -1543 206 -1536
tri 206 -1543 213 -1536 sw
rect 196 -1568 213 -1543
rect 337 -1568 354 -1536
rect 536 -1568 551 -1526
rect 579 -1568 594 -1526
rect 776 -1543 786 -1536
tri 786 -1543 793 -1536 sw
rect 776 -1568 793 -1543
rect 917 -1568 934 -1536
rect 1116 -1568 1131 -1526
rect 1159 -1568 1174 -1526
rect 1356 -1543 1366 -1536
tri 1366 -1543 1373 -1536 sw
rect 1356 -1568 1373 -1543
rect 1497 -1568 1514 -1536
rect 1696 -1568 1711 -1526
rect 1739 -1568 1754 -1526
rect 1936 -1543 1946 -1536
tri 1946 -1543 1953 -1536 sw
rect 1936 -1568 1953 -1543
rect 2077 -1568 2094 -1536
rect 2276 -1568 2291 -1526
rect 2319 -1568 2334 -1526
rect 2516 -1543 2526 -1536
tri 2526 -1543 2533 -1536 sw
rect 2516 -1568 2533 -1543
rect 2657 -1568 2674 -1536
rect 2856 -1568 2871 -1526
rect 2899 -1568 2914 -1526
rect 3096 -1543 3106 -1536
tri 3106 -1543 3113 -1536 sw
rect 3096 -1568 3113 -1543
rect 3237 -1568 3254 -1536
rect 3436 -1568 3451 -1526
rect 3479 -1568 3494 -1526
rect 3676 -1543 3686 -1536
tri 3686 -1543 3693 -1536 sw
rect 3676 -1568 3693 -1543
rect 3817 -1568 3834 -1536
rect 4016 -1568 4031 -1526
rect 4059 -1568 4074 -1526
rect 4256 -1543 4266 -1536
tri 4266 -1543 4273 -1536 sw
rect 4256 -1568 4273 -1543
rect 4397 -1568 4414 -1536
rect 4596 -1568 4611 -1526
rect 5601 -1423 5616 -1395
rect 5683 -1423 5698 -1394
rect 5873 -1423 5888 -1395
rect 5954 -1423 5969 -1395
rect 6181 -1423 6196 -1395
rect 6263 -1423 6278 -1394
rect 6453 -1423 6468 -1395
rect 6534 -1423 6549 -1395
rect 6761 -1423 6776 -1395
rect 6843 -1423 6858 -1394
rect 259 -1606 291 -1592
rect 839 -1606 871 -1592
rect 1419 -1606 1451 -1592
rect 1999 -1606 2031 -1592
rect 2579 -1606 2611 -1592
rect 3159 -1606 3191 -1592
rect 3739 -1606 3771 -1592
rect 4639 -1569 4654 -1527
rect 4836 -1544 4846 -1537
tri 4846 -1544 4853 -1537 sw
rect 4836 -1569 4853 -1544
rect 4977 -1569 4994 -1537
rect 5176 -1569 5191 -1527
rect 5219 -1569 5234 -1527
rect 5416 -1544 5426 -1537
tri 5426 -1544 5433 -1537 sw
rect 5416 -1569 5433 -1544
rect 5557 -1569 5574 -1537
rect 5756 -1569 5771 -1527
rect 5799 -1569 5814 -1527
rect 5996 -1544 6006 -1537
tri 6006 -1544 6013 -1537 sw
rect 5996 -1569 6013 -1544
rect 6137 -1569 6154 -1537
rect 6336 -1569 6351 -1527
rect 6379 -1569 6394 -1527
rect 6576 -1544 6586 -1537
tri 6586 -1544 6593 -1537 sw
rect 6576 -1569 6593 -1544
rect 6717 -1569 6734 -1537
rect 6916 -1569 6931 -1527
rect 4319 -1606 4351 -1592
rect 4899 -1607 4931 -1593
rect 5479 -1607 5511 -1593
rect 6059 -1607 6091 -1593
rect 6639 -1607 6671 -1593
rect 73 -1692 88 -1664
rect 154 -1692 169 -1664
rect 381 -1692 396 -1664
rect 463 -1692 478 -1663
rect 653 -1692 668 -1664
rect 734 -1692 749 -1664
rect 961 -1692 976 -1664
rect 1043 -1692 1058 -1663
rect 1233 -1692 1248 -1664
rect 1314 -1692 1329 -1664
rect 1541 -1692 1556 -1664
rect 1623 -1692 1638 -1663
rect 1813 -1692 1828 -1664
rect 1894 -1692 1909 -1664
rect 2121 -1692 2136 -1664
rect 2203 -1692 2218 -1663
rect 2393 -1692 2408 -1664
rect 2474 -1692 2489 -1664
rect 2701 -1692 2716 -1664
rect 2783 -1692 2798 -1663
rect 2973 -1692 2988 -1664
rect 3054 -1692 3069 -1664
rect 3281 -1692 3296 -1664
rect 3363 -1692 3378 -1663
rect 3553 -1692 3568 -1664
rect 3634 -1692 3649 -1664
rect 3861 -1692 3876 -1664
rect 3943 -1692 3958 -1663
rect 4133 -1692 4148 -1664
rect 4214 -1692 4229 -1664
rect 4441 -1692 4456 -1664
rect 4523 -1692 4538 -1663
rect 4713 -1693 4728 -1665
rect 4794 -1693 4809 -1665
rect 5021 -1693 5036 -1665
rect 5103 -1693 5118 -1664
rect 5293 -1693 5308 -1665
rect 5374 -1693 5389 -1665
rect -1 -1838 14 -1796
rect 196 -1813 206 -1806
tri 206 -1813 213 -1806 sw
rect 196 -1838 213 -1813
rect 337 -1838 354 -1806
rect 536 -1838 551 -1796
rect 579 -1838 594 -1796
rect 776 -1813 786 -1806
tri 786 -1813 793 -1806 sw
rect 776 -1838 793 -1813
rect 917 -1838 934 -1806
rect 1116 -1838 1131 -1796
rect 1159 -1838 1174 -1796
rect 1356 -1813 1366 -1806
tri 1366 -1813 1373 -1806 sw
rect 1356 -1838 1373 -1813
rect 1497 -1838 1514 -1806
rect 1696 -1838 1711 -1796
rect 1739 -1838 1754 -1796
rect 1936 -1813 1946 -1806
tri 1946 -1813 1953 -1806 sw
rect 1936 -1838 1953 -1813
rect 2077 -1838 2094 -1806
rect 2276 -1838 2291 -1796
rect 2319 -1838 2334 -1796
rect 2516 -1813 2526 -1806
tri 2526 -1813 2533 -1806 sw
rect 2516 -1838 2533 -1813
rect 2657 -1838 2674 -1806
rect 2856 -1838 2871 -1796
rect 2899 -1838 2914 -1796
rect 3096 -1813 3106 -1806
tri 3106 -1813 3113 -1806 sw
rect 3096 -1838 3113 -1813
rect 3237 -1838 3254 -1806
rect 3436 -1838 3451 -1796
rect 3479 -1838 3494 -1796
rect 3676 -1813 3686 -1806
tri 3686 -1813 3693 -1806 sw
rect 3676 -1838 3693 -1813
rect 3817 -1838 3834 -1806
rect 4016 -1838 4031 -1796
rect 4059 -1838 4074 -1796
rect 4256 -1813 4266 -1806
tri 4266 -1813 4273 -1806 sw
rect 4256 -1838 4273 -1813
rect 4397 -1838 4414 -1806
rect 4596 -1838 4611 -1796
rect 5601 -1693 5616 -1665
rect 5683 -1693 5698 -1664
rect 5873 -1693 5888 -1665
rect 5954 -1693 5969 -1665
rect 6181 -1693 6196 -1665
rect 6263 -1693 6278 -1664
rect 6453 -1693 6468 -1665
rect 6534 -1693 6549 -1665
rect 6761 -1693 6776 -1665
rect 6843 -1693 6858 -1664
rect 259 -1876 291 -1862
rect 839 -1876 871 -1862
rect 1419 -1876 1451 -1862
rect 1999 -1876 2031 -1862
rect 2579 -1876 2611 -1862
rect 3159 -1876 3191 -1862
rect 3739 -1876 3771 -1862
rect 4639 -1839 4654 -1797
rect 4836 -1814 4846 -1807
tri 4846 -1814 4853 -1807 sw
rect 4836 -1839 4853 -1814
rect 4977 -1839 4994 -1807
rect 5176 -1839 5191 -1797
rect 5219 -1839 5234 -1797
rect 5416 -1814 5426 -1807
tri 5426 -1814 5433 -1807 sw
rect 5416 -1839 5433 -1814
rect 5557 -1839 5574 -1807
rect 5756 -1839 5771 -1797
rect 5799 -1839 5814 -1797
rect 5996 -1814 6006 -1807
tri 6006 -1814 6013 -1807 sw
rect 5996 -1839 6013 -1814
rect 6137 -1839 6154 -1807
rect 6336 -1839 6351 -1797
rect 6379 -1839 6394 -1797
rect 6576 -1814 6586 -1807
tri 6586 -1814 6593 -1807 sw
rect 6576 -1839 6593 -1814
rect 6717 -1839 6734 -1807
rect 6916 -1839 6931 -1797
rect 4319 -1876 4351 -1862
rect 4899 -1877 4931 -1863
rect 5479 -1877 5511 -1863
rect 6059 -1877 6091 -1863
rect 6639 -1877 6671 -1863
rect 73 -1962 88 -1934
rect 154 -1962 169 -1934
rect 381 -1962 396 -1934
rect 463 -1962 478 -1933
rect 653 -1962 668 -1934
rect 734 -1962 749 -1934
rect 961 -1962 976 -1934
rect 1043 -1962 1058 -1933
rect 1233 -1962 1248 -1934
rect 1314 -1962 1329 -1934
rect 1541 -1962 1556 -1934
rect 1623 -1962 1638 -1933
rect 1813 -1962 1828 -1934
rect 1894 -1962 1909 -1934
rect 2121 -1962 2136 -1934
rect 2203 -1962 2218 -1933
rect 2393 -1962 2408 -1934
rect 2474 -1962 2489 -1934
rect 2701 -1962 2716 -1934
rect 2783 -1962 2798 -1933
rect 2973 -1962 2988 -1934
rect 3054 -1962 3069 -1934
rect 3281 -1962 3296 -1934
rect 3363 -1962 3378 -1933
rect 3553 -1962 3568 -1934
rect 3634 -1962 3649 -1934
rect 3861 -1962 3876 -1934
rect 3943 -1962 3958 -1933
rect 4133 -1962 4148 -1934
rect 4214 -1962 4229 -1934
rect 4441 -1962 4456 -1934
rect 4523 -1962 4538 -1933
rect 4713 -1963 4728 -1935
rect 4794 -1963 4809 -1935
rect 5021 -1963 5036 -1935
rect 5103 -1963 5118 -1934
rect 5293 -1963 5308 -1935
rect 5374 -1963 5389 -1935
rect -1 -2108 14 -2066
rect 196 -2083 206 -2076
tri 206 -2083 213 -2076 sw
rect 196 -2108 213 -2083
rect 337 -2108 354 -2076
rect 536 -2108 551 -2066
rect 579 -2108 594 -2066
rect 776 -2083 786 -2076
tri 786 -2083 793 -2076 sw
rect 776 -2108 793 -2083
rect 917 -2108 934 -2076
rect 1116 -2108 1131 -2066
rect 1159 -2108 1174 -2066
rect 1356 -2083 1366 -2076
tri 1366 -2083 1373 -2076 sw
rect 1356 -2108 1373 -2083
rect 1497 -2108 1514 -2076
rect 1696 -2108 1711 -2066
rect 1739 -2108 1754 -2066
rect 1936 -2083 1946 -2076
tri 1946 -2083 1953 -2076 sw
rect 1936 -2108 1953 -2083
rect 2077 -2108 2094 -2076
rect 2276 -2108 2291 -2066
rect 2319 -2108 2334 -2066
rect 2516 -2083 2526 -2076
tri 2526 -2083 2533 -2076 sw
rect 2516 -2108 2533 -2083
rect 2657 -2108 2674 -2076
rect 2856 -2108 2871 -2066
rect 2899 -2108 2914 -2066
rect 3096 -2083 3106 -2076
tri 3106 -2083 3113 -2076 sw
rect 3096 -2108 3113 -2083
rect 3237 -2108 3254 -2076
rect 3436 -2108 3451 -2066
rect 3479 -2108 3494 -2066
rect 3676 -2083 3686 -2076
tri 3686 -2083 3693 -2076 sw
rect 3676 -2108 3693 -2083
rect 3817 -2108 3834 -2076
rect 4016 -2108 4031 -2066
rect 4059 -2108 4074 -2066
rect 4256 -2083 4266 -2076
tri 4266 -2083 4273 -2076 sw
rect 4256 -2108 4273 -2083
rect 4397 -2108 4414 -2076
rect 4596 -2108 4611 -2066
rect 5601 -1963 5616 -1935
rect 5683 -1963 5698 -1934
rect 5873 -1963 5888 -1935
rect 5954 -1963 5969 -1935
rect 6181 -1963 6196 -1935
rect 6263 -1963 6278 -1934
rect 6453 -1963 6468 -1935
rect 6534 -1963 6549 -1935
rect 6761 -1963 6776 -1935
rect 6843 -1963 6858 -1934
rect 259 -2146 291 -2132
rect 839 -2146 871 -2132
rect 1419 -2146 1451 -2132
rect 1999 -2146 2031 -2132
rect 2579 -2146 2611 -2132
rect 3159 -2146 3191 -2132
rect 3739 -2146 3771 -2132
rect 4639 -2109 4654 -2067
rect 4836 -2084 4846 -2077
tri 4846 -2084 4853 -2077 sw
rect 4836 -2109 4853 -2084
rect 4977 -2109 4994 -2077
rect 5176 -2109 5191 -2067
rect 5219 -2109 5234 -2067
rect 5416 -2084 5426 -2077
tri 5426 -2084 5433 -2077 sw
rect 5416 -2109 5433 -2084
rect 5557 -2109 5574 -2077
rect 5756 -2109 5771 -2067
rect 5799 -2109 5814 -2067
rect 5996 -2084 6006 -2077
tri 6006 -2084 6013 -2077 sw
rect 5996 -2109 6013 -2084
rect 6137 -2109 6154 -2077
rect 6336 -2109 6351 -2067
rect 6379 -2109 6394 -2067
rect 6576 -2084 6586 -2077
tri 6586 -2084 6593 -2077 sw
rect 6576 -2109 6593 -2084
rect 6717 -2109 6734 -2077
rect 6916 -2109 6931 -2067
rect 4319 -2146 4351 -2132
rect 4899 -2147 4931 -2133
rect 5479 -2147 5511 -2133
rect 6059 -2147 6091 -2133
rect 6639 -2147 6671 -2133
<< pdiffc >>
rect 259 2130 291 2144
rect 197 2078 212 2106
rect 338 2090 350 2106
tri 338 2078 350 2090 ne
rect 839 2130 871 2144
rect 777 2078 792 2106
rect 918 2090 930 2106
tri 918 2078 930 2090 ne
rect 1419 2130 1451 2144
rect 1357 2078 1372 2106
rect 1498 2090 1510 2106
tri 1498 2078 1510 2090 ne
rect 1999 2130 2031 2144
rect 1937 2078 1952 2106
rect 2078 2090 2090 2106
tri 2078 2078 2090 2090 ne
rect 2579 2130 2611 2144
rect 2517 2078 2532 2106
rect 2658 2090 2670 2106
tri 2658 2078 2670 2090 ne
rect 3159 2130 3191 2144
rect 3097 2078 3112 2106
rect 3238 2090 3250 2106
tri 3238 2078 3250 2090 ne
rect 3739 2130 3771 2144
rect 3677 2078 3692 2106
rect 3818 2090 3830 2106
tri 3818 2078 3830 2090 ne
rect 4319 2130 4351 2144
rect 4257 2078 4272 2106
rect 4398 2090 4410 2106
tri 4398 2078 4410 2090 ne
rect 4899 2130 4931 2144
rect 4837 2078 4852 2106
rect 4978 2090 4990 2106
tri 4978 2078 4990 2090 ne
rect 5479 2130 5511 2144
rect 5417 2078 5432 2106
rect 5558 2090 5570 2106
tri 5558 2078 5570 2090 ne
rect 6059 2130 6091 2144
rect 5997 2078 6012 2106
rect 6138 2090 6150 2106
tri 6138 2078 6150 2090 ne
rect 6639 2130 6671 2144
rect 6577 2078 6592 2106
rect 6718 2090 6730 2106
tri 6718 2078 6730 2090 ne
rect 259 1860 291 1874
rect 197 1808 212 1836
rect 338 1820 350 1836
tri 338 1808 350 1820 ne
rect 839 1860 871 1874
rect 777 1808 792 1836
rect 918 1820 930 1836
tri 918 1808 930 1820 ne
rect 1419 1860 1451 1874
rect 1357 1808 1372 1836
rect 1498 1820 1510 1836
tri 1498 1808 1510 1820 ne
rect 1999 1860 2031 1874
rect 1937 1808 1952 1836
rect 2078 1820 2090 1836
tri 2078 1808 2090 1820 ne
rect 2579 1860 2611 1874
rect 2517 1808 2532 1836
rect 2658 1820 2670 1836
tri 2658 1808 2670 1820 ne
rect 3159 1860 3191 1874
rect 3097 1808 3112 1836
rect 3238 1820 3250 1836
tri 3238 1808 3250 1820 ne
rect 3739 1860 3771 1874
rect 3677 1808 3692 1836
rect 3818 1820 3830 1836
tri 3818 1808 3830 1820 ne
rect 4319 1860 4351 1874
rect 4257 1808 4272 1836
rect 4398 1820 4410 1836
tri 4398 1808 4410 1820 ne
rect 4899 1860 4931 1874
rect 4837 1808 4852 1836
rect 4978 1820 4990 1836
tri 4978 1808 4990 1820 ne
rect 5479 1860 5511 1874
rect 5417 1808 5432 1836
rect 5558 1820 5570 1836
tri 5558 1808 5570 1820 ne
rect 6059 1860 6091 1874
rect 5997 1808 6012 1836
rect 6138 1820 6150 1836
tri 6138 1808 6150 1820 ne
rect 6639 1860 6671 1874
rect 6577 1808 6592 1836
rect 6718 1820 6730 1836
tri 6718 1808 6730 1820 ne
rect 259 1590 291 1604
rect 197 1538 212 1566
rect 338 1550 350 1566
tri 338 1538 350 1550 ne
rect 839 1590 871 1604
rect 777 1538 792 1566
rect 918 1550 930 1566
tri 918 1538 930 1550 ne
rect 1419 1590 1451 1604
rect 1357 1538 1372 1566
rect 1498 1550 1510 1566
tri 1498 1538 1510 1550 ne
rect 1999 1590 2031 1604
rect 1937 1538 1952 1566
rect 2078 1550 2090 1566
tri 2078 1538 2090 1550 ne
rect 2579 1590 2611 1604
rect 2517 1538 2532 1566
rect 2658 1550 2670 1566
tri 2658 1538 2670 1550 ne
rect 3159 1590 3191 1604
rect 3097 1538 3112 1566
rect 3238 1550 3250 1566
tri 3238 1538 3250 1550 ne
rect 3739 1590 3771 1604
rect 3677 1538 3692 1566
rect 3818 1550 3830 1566
tri 3818 1538 3830 1550 ne
rect 4319 1590 4351 1604
rect 4257 1538 4272 1566
rect 4398 1550 4410 1566
tri 4398 1538 4410 1550 ne
rect 4899 1590 4931 1604
rect 4837 1538 4852 1566
rect 4978 1550 4990 1566
tri 4978 1538 4990 1550 ne
rect 5479 1590 5511 1604
rect 5417 1538 5432 1566
rect 5558 1550 5570 1566
tri 5558 1538 5570 1550 ne
rect 6059 1590 6091 1604
rect 5997 1538 6012 1566
rect 6138 1550 6150 1566
tri 6138 1538 6150 1550 ne
rect 6639 1590 6671 1604
rect 6577 1538 6592 1566
rect 6718 1550 6730 1566
tri 6718 1538 6730 1550 ne
rect 259 1320 291 1334
rect 197 1268 212 1296
rect 338 1280 350 1296
tri 338 1268 350 1280 ne
rect 839 1320 871 1334
rect 777 1268 792 1296
rect 918 1280 930 1296
tri 918 1268 930 1280 ne
rect 1419 1320 1451 1334
rect 1357 1268 1372 1296
rect 1498 1280 1510 1296
tri 1498 1268 1510 1280 ne
rect 1999 1320 2031 1334
rect 1937 1268 1952 1296
rect 2078 1280 2090 1296
tri 2078 1268 2090 1280 ne
rect 2579 1320 2611 1334
rect 2517 1268 2532 1296
rect 2658 1280 2670 1296
tri 2658 1268 2670 1280 ne
rect 3159 1320 3191 1334
rect 3097 1268 3112 1296
rect 3238 1280 3250 1296
tri 3238 1268 3250 1280 ne
rect 3739 1320 3771 1334
rect 3677 1268 3692 1296
rect 3818 1280 3830 1296
tri 3818 1268 3830 1280 ne
rect 4319 1320 4351 1334
rect 4257 1268 4272 1296
rect 4398 1280 4410 1296
tri 4398 1268 4410 1280 ne
rect 4899 1320 4931 1334
rect 4837 1268 4852 1296
rect 4978 1280 4990 1296
tri 4978 1268 4990 1280 ne
rect 5479 1320 5511 1334
rect 5417 1268 5432 1296
rect 5558 1280 5570 1296
tri 5558 1268 5570 1280 ne
rect 6059 1320 6091 1334
rect 5997 1268 6012 1296
rect 6138 1280 6150 1296
tri 6138 1268 6150 1280 ne
rect 6639 1320 6671 1334
rect 6577 1268 6592 1296
rect 6718 1280 6730 1296
tri 6718 1268 6730 1280 ne
rect 259 1050 291 1064
rect 197 998 212 1026
rect 338 1010 350 1026
tri 338 998 350 1010 ne
rect 839 1050 871 1064
rect 777 998 792 1026
rect 918 1010 930 1026
tri 918 998 930 1010 ne
rect 1419 1050 1451 1064
rect 1357 998 1372 1026
rect 1498 1010 1510 1026
tri 1498 998 1510 1010 ne
rect 1999 1050 2031 1064
rect 1937 998 1952 1026
rect 2078 1010 2090 1026
tri 2078 998 2090 1010 ne
rect 2579 1050 2611 1064
rect 2517 998 2532 1026
rect 2658 1010 2670 1026
tri 2658 998 2670 1010 ne
rect 3159 1050 3191 1064
rect 3097 998 3112 1026
rect 3238 1010 3250 1026
tri 3238 998 3250 1010 ne
rect 3739 1050 3771 1064
rect 3677 998 3692 1026
rect 3818 1010 3830 1026
tri 3818 998 3830 1010 ne
rect 4319 1050 4351 1064
rect 4257 998 4272 1026
rect 4398 1010 4410 1026
tri 4398 998 4410 1010 ne
rect 4899 1049 4931 1063
rect 4837 997 4852 1025
rect 4978 1009 4990 1025
tri 4978 997 4990 1009 ne
rect 5479 1049 5511 1063
rect 5417 997 5432 1025
rect 5558 1009 5570 1025
tri 5558 997 5570 1009 ne
rect 6059 1049 6091 1063
rect 5997 997 6012 1025
rect 6138 1009 6150 1025
tri 6138 997 6150 1009 ne
rect 6639 1049 6671 1063
rect 6577 997 6592 1025
rect 6718 1009 6730 1025
tri 6718 997 6730 1009 ne
rect 259 780 291 794
rect 197 728 212 756
rect 338 740 350 756
tri 338 728 350 740 ne
rect 839 780 871 794
rect 777 728 792 756
rect 918 740 930 756
tri 918 728 930 740 ne
rect 1419 780 1451 794
rect 1357 728 1372 756
rect 1498 740 1510 756
tri 1498 728 1510 740 ne
rect 1999 780 2031 794
rect 1937 728 1952 756
rect 2078 740 2090 756
tri 2078 728 2090 740 ne
rect 2579 780 2611 794
rect 2517 728 2532 756
rect 2658 740 2670 756
tri 2658 728 2670 740 ne
rect 3159 780 3191 794
rect 3097 728 3112 756
rect 3238 740 3250 756
tri 3238 728 3250 740 ne
rect 3739 780 3771 794
rect 3677 728 3692 756
rect 3818 740 3830 756
tri 3818 728 3830 740 ne
rect 4319 780 4351 794
rect 4257 728 4272 756
rect 4398 740 4410 756
tri 4398 728 4410 740 ne
rect 4899 779 4931 793
rect 4837 727 4852 755
rect 4978 739 4990 755
tri 4978 727 4990 739 ne
rect 5479 779 5511 793
rect 5417 727 5432 755
rect 5558 739 5570 755
tri 5558 727 5570 739 ne
rect 6059 779 6091 793
rect 5997 727 6012 755
rect 6138 739 6150 755
tri 6138 727 6150 739 ne
rect 6639 779 6671 793
rect 6577 727 6592 755
rect 6718 739 6730 755
tri 6718 727 6730 739 ne
rect 259 510 291 524
rect 197 458 212 486
rect 338 470 350 486
tri 338 458 350 470 ne
rect 839 510 871 524
rect 777 458 792 486
rect 918 470 930 486
tri 918 458 930 470 ne
rect 1419 510 1451 524
rect 1357 458 1372 486
rect 1498 470 1510 486
tri 1498 458 1510 470 ne
rect 1999 510 2031 524
rect 1937 458 1952 486
rect 2078 470 2090 486
tri 2078 458 2090 470 ne
rect 2579 510 2611 524
rect 2517 458 2532 486
rect 2658 470 2670 486
tri 2658 458 2670 470 ne
rect 3159 510 3191 524
rect 3097 458 3112 486
rect 3238 470 3250 486
tri 3238 458 3250 470 ne
rect 3739 510 3771 524
rect 3677 458 3692 486
rect 3818 470 3830 486
tri 3818 458 3830 470 ne
rect 4319 510 4351 524
rect 4257 458 4272 486
rect 4398 470 4410 486
tri 4398 458 4410 470 ne
rect 4899 509 4931 523
rect 4837 457 4852 485
rect 4978 469 4990 485
tri 4978 457 4990 469 ne
rect 5479 509 5511 523
rect 5417 457 5432 485
rect 5558 469 5570 485
tri 5558 457 5570 469 ne
rect 6059 509 6091 523
rect 5997 457 6012 485
rect 6138 469 6150 485
tri 6138 457 6150 469 ne
rect 6639 509 6671 523
rect 6577 457 6592 485
rect 6718 469 6730 485
tri 6718 457 6730 469 ne
rect 259 240 291 254
rect 197 188 212 216
rect 338 200 350 216
tri 338 188 350 200 ne
rect 839 240 871 254
rect 777 188 792 216
rect 918 200 930 216
tri 918 188 930 200 ne
rect 1419 240 1451 254
rect 1357 188 1372 216
rect 1498 200 1510 216
tri 1498 188 1510 200 ne
rect 1999 240 2031 254
rect 1937 188 1952 216
rect 2078 200 2090 216
tri 2078 188 2090 200 ne
rect 2579 240 2611 254
rect 2517 188 2532 216
rect 2658 200 2670 216
tri 2658 188 2670 200 ne
rect 3159 240 3191 254
rect 3097 188 3112 216
rect 3238 200 3250 216
tri 3238 188 3250 200 ne
rect 3739 240 3771 254
rect 3677 188 3692 216
rect 3818 200 3830 216
tri 3818 188 3830 200 ne
rect 4319 240 4351 254
rect 4257 188 4272 216
rect 4398 200 4410 216
tri 4398 188 4410 200 ne
rect 4899 239 4931 253
rect 4837 187 4852 215
rect 4978 199 4990 215
tri 4978 187 4990 199 ne
rect 5479 239 5511 253
rect 5417 187 5432 215
rect 5558 199 5570 215
tri 5558 187 5570 199 ne
rect 6059 239 6091 253
rect 5997 187 6012 215
rect 6138 199 6150 215
tri 6138 187 6150 199 ne
rect 6639 239 6671 253
rect 6577 187 6592 215
rect 6718 199 6730 215
tri 6718 187 6730 199 ne
rect 259 -30 291 -16
rect 197 -82 212 -54
rect 338 -70 350 -54
tri 338 -82 350 -70 ne
rect 839 -30 871 -16
rect 777 -82 792 -54
rect 918 -70 930 -54
tri 918 -82 930 -70 ne
rect 1419 -30 1451 -16
rect 1357 -82 1372 -54
rect 1498 -70 1510 -54
tri 1498 -82 1510 -70 ne
rect 1999 -30 2031 -16
rect 1937 -82 1952 -54
rect 2078 -70 2090 -54
tri 2078 -82 2090 -70 ne
rect 2579 -30 2611 -16
rect 2517 -82 2532 -54
rect 2658 -70 2670 -54
tri 2658 -82 2670 -70 ne
rect 3159 -30 3191 -16
rect 3097 -82 3112 -54
rect 3238 -70 3250 -54
tri 3238 -82 3250 -70 ne
rect 3739 -30 3771 -16
rect 3677 -82 3692 -54
rect 3818 -70 3830 -54
tri 3818 -82 3830 -70 ne
rect 4319 -30 4351 -16
rect 4257 -82 4272 -54
rect 4398 -70 4410 -54
tri 4398 -82 4410 -70 ne
rect 4899 -31 4931 -17
rect 4837 -83 4852 -55
rect 4978 -71 4990 -55
tri 4978 -83 4990 -71 ne
rect 5479 -31 5511 -17
rect 5417 -83 5432 -55
rect 5558 -71 5570 -55
tri 5558 -83 5570 -71 ne
rect 6059 -31 6091 -17
rect 5997 -83 6012 -55
rect 6138 -71 6150 -55
tri 6138 -83 6150 -71 ne
rect 6639 -31 6671 -17
rect 6577 -83 6592 -55
rect 6718 -71 6730 -55
tri 6718 -83 6730 -71 ne
rect 259 -300 291 -286
rect 197 -352 212 -324
rect 338 -340 350 -324
tri 338 -352 350 -340 ne
rect 839 -300 871 -286
rect 777 -352 792 -324
rect 918 -340 930 -324
tri 918 -352 930 -340 ne
rect 1419 -300 1451 -286
rect 1357 -352 1372 -324
rect 1498 -340 1510 -324
tri 1498 -352 1510 -340 ne
rect 1999 -300 2031 -286
rect 1937 -352 1952 -324
rect 2078 -340 2090 -324
tri 2078 -352 2090 -340 ne
rect 2579 -300 2611 -286
rect 2517 -352 2532 -324
rect 2658 -340 2670 -324
tri 2658 -352 2670 -340 ne
rect 3159 -300 3191 -286
rect 3097 -352 3112 -324
rect 3238 -340 3250 -324
tri 3238 -352 3250 -340 ne
rect 3739 -300 3771 -286
rect 3677 -352 3692 -324
rect 3818 -340 3830 -324
tri 3818 -352 3830 -340 ne
rect 4319 -300 4351 -286
rect 4257 -352 4272 -324
rect 4398 -340 4410 -324
tri 4398 -352 4410 -340 ne
rect 4899 -301 4931 -287
rect 4837 -353 4852 -325
rect 4978 -341 4990 -325
tri 4978 -353 4990 -341 ne
rect 5479 -301 5511 -287
rect 5417 -353 5432 -325
rect 5558 -341 5570 -325
tri 5558 -353 5570 -341 ne
rect 6059 -301 6091 -287
rect 5997 -353 6012 -325
rect 6138 -341 6150 -325
tri 6138 -353 6150 -341 ne
rect 6639 -301 6671 -287
rect 6577 -353 6592 -325
rect 6718 -341 6730 -325
tri 6718 -353 6730 -341 ne
rect 259 -570 291 -556
rect 197 -622 212 -594
rect 338 -610 350 -594
tri 338 -622 350 -610 ne
rect 839 -570 871 -556
rect 777 -622 792 -594
rect 918 -610 930 -594
tri 918 -622 930 -610 ne
rect 1419 -570 1451 -556
rect 1357 -622 1372 -594
rect 1498 -610 1510 -594
tri 1498 -622 1510 -610 ne
rect 1999 -570 2031 -556
rect 1937 -622 1952 -594
rect 2078 -610 2090 -594
tri 2078 -622 2090 -610 ne
rect 2579 -570 2611 -556
rect 2517 -622 2532 -594
rect 2658 -610 2670 -594
tri 2658 -622 2670 -610 ne
rect 3159 -570 3191 -556
rect 3097 -622 3112 -594
rect 3238 -610 3250 -594
tri 3238 -622 3250 -610 ne
rect 3739 -570 3771 -556
rect 3677 -622 3692 -594
rect 3818 -610 3830 -594
tri 3818 -622 3830 -610 ne
rect 4319 -570 4351 -556
rect 4257 -622 4272 -594
rect 4398 -610 4410 -594
tri 4398 -622 4410 -610 ne
rect 4899 -571 4931 -557
rect 4837 -623 4852 -595
rect 4978 -611 4990 -595
tri 4978 -623 4990 -611 ne
rect 5479 -571 5511 -557
rect 5417 -623 5432 -595
rect 5558 -611 5570 -595
tri 5558 -623 5570 -611 ne
rect 6059 -571 6091 -557
rect 5997 -623 6012 -595
rect 6138 -611 6150 -595
tri 6138 -623 6150 -611 ne
rect 6639 -571 6671 -557
rect 6577 -623 6592 -595
rect 6718 -611 6730 -595
tri 6718 -623 6730 -611 ne
rect 259 -840 291 -826
rect 197 -892 212 -864
rect 338 -880 350 -864
tri 338 -892 350 -880 ne
rect 839 -840 871 -826
rect 777 -892 792 -864
rect 918 -880 930 -864
tri 918 -892 930 -880 ne
rect 1419 -840 1451 -826
rect 1357 -892 1372 -864
rect 1498 -880 1510 -864
tri 1498 -892 1510 -880 ne
rect 1999 -840 2031 -826
rect 1937 -892 1952 -864
rect 2078 -880 2090 -864
tri 2078 -892 2090 -880 ne
rect 2579 -840 2611 -826
rect 2517 -892 2532 -864
rect 2658 -880 2670 -864
tri 2658 -892 2670 -880 ne
rect 3159 -840 3191 -826
rect 3097 -892 3112 -864
rect 3238 -880 3250 -864
tri 3238 -892 3250 -880 ne
rect 3739 -840 3771 -826
rect 3677 -892 3692 -864
rect 3818 -880 3830 -864
tri 3818 -892 3830 -880 ne
rect 4319 -840 4351 -826
rect 4257 -892 4272 -864
rect 4398 -880 4410 -864
tri 4398 -892 4410 -880 ne
rect 4899 -841 4931 -827
rect 4837 -893 4852 -865
rect 4978 -881 4990 -865
tri 4978 -893 4990 -881 ne
rect 5479 -841 5511 -827
rect 5417 -893 5432 -865
rect 5558 -881 5570 -865
tri 5558 -893 5570 -881 ne
rect 6059 -841 6091 -827
rect 5997 -893 6012 -865
rect 6138 -881 6150 -865
tri 6138 -893 6150 -881 ne
rect 6639 -841 6671 -827
rect 6577 -893 6592 -865
rect 6718 -881 6730 -865
tri 6718 -893 6730 -881 ne
rect 259 -1110 291 -1096
rect 197 -1162 212 -1134
rect 338 -1150 350 -1134
tri 338 -1162 350 -1150 ne
rect 839 -1110 871 -1096
rect 777 -1162 792 -1134
rect 918 -1150 930 -1134
tri 918 -1162 930 -1150 ne
rect 1419 -1110 1451 -1096
rect 1357 -1162 1372 -1134
rect 1498 -1150 1510 -1134
tri 1498 -1162 1510 -1150 ne
rect 1999 -1110 2031 -1096
rect 1937 -1162 1952 -1134
rect 2078 -1150 2090 -1134
tri 2078 -1162 2090 -1150 ne
rect 2579 -1110 2611 -1096
rect 2517 -1162 2532 -1134
rect 2658 -1150 2670 -1134
tri 2658 -1162 2670 -1150 ne
rect 3159 -1110 3191 -1096
rect 3097 -1162 3112 -1134
rect 3238 -1150 3250 -1134
tri 3238 -1162 3250 -1150 ne
rect 3739 -1110 3771 -1096
rect 3677 -1162 3692 -1134
rect 3818 -1150 3830 -1134
tri 3818 -1162 3830 -1150 ne
rect 4319 -1110 4351 -1096
rect 4257 -1162 4272 -1134
rect 4398 -1150 4410 -1134
tri 4398 -1162 4410 -1150 ne
rect 4899 -1111 4931 -1097
rect 4837 -1163 4852 -1135
rect 4978 -1151 4990 -1135
tri 4978 -1163 4990 -1151 ne
rect 5479 -1111 5511 -1097
rect 5417 -1163 5432 -1135
rect 5558 -1151 5570 -1135
tri 5558 -1163 5570 -1151 ne
rect 6059 -1111 6091 -1097
rect 5997 -1163 6012 -1135
rect 6138 -1151 6150 -1135
tri 6138 -1163 6150 -1151 ne
rect 6639 -1111 6671 -1097
rect 6577 -1163 6592 -1135
rect 6718 -1151 6730 -1135
tri 6718 -1163 6730 -1151 ne
rect 259 -1380 291 -1366
rect 197 -1432 212 -1404
rect 338 -1420 350 -1404
tri 338 -1432 350 -1420 ne
rect 839 -1380 871 -1366
rect 777 -1432 792 -1404
rect 918 -1420 930 -1404
tri 918 -1432 930 -1420 ne
rect 1419 -1380 1451 -1366
rect 1357 -1432 1372 -1404
rect 1498 -1420 1510 -1404
tri 1498 -1432 1510 -1420 ne
rect 1999 -1380 2031 -1366
rect 1937 -1432 1952 -1404
rect 2078 -1420 2090 -1404
tri 2078 -1432 2090 -1420 ne
rect 2579 -1380 2611 -1366
rect 2517 -1432 2532 -1404
rect 2658 -1420 2670 -1404
tri 2658 -1432 2670 -1420 ne
rect 3159 -1380 3191 -1366
rect 3097 -1432 3112 -1404
rect 3238 -1420 3250 -1404
tri 3238 -1432 3250 -1420 ne
rect 3739 -1380 3771 -1366
rect 3677 -1432 3692 -1404
rect 3818 -1420 3830 -1404
tri 3818 -1432 3830 -1420 ne
rect 4319 -1380 4351 -1366
rect 4257 -1432 4272 -1404
rect 4398 -1420 4410 -1404
tri 4398 -1432 4410 -1420 ne
rect 4899 -1381 4931 -1367
rect 4837 -1433 4852 -1405
rect 4978 -1421 4990 -1405
tri 4978 -1433 4990 -1421 ne
rect 5479 -1381 5511 -1367
rect 5417 -1433 5432 -1405
rect 5558 -1421 5570 -1405
tri 5558 -1433 5570 -1421 ne
rect 6059 -1381 6091 -1367
rect 5997 -1433 6012 -1405
rect 6138 -1421 6150 -1405
tri 6138 -1433 6150 -1421 ne
rect 6639 -1381 6671 -1367
rect 6577 -1433 6592 -1405
rect 6718 -1421 6730 -1405
tri 6718 -1433 6730 -1421 ne
rect 259 -1650 291 -1636
rect 197 -1702 212 -1674
rect 338 -1690 350 -1674
tri 338 -1702 350 -1690 ne
rect 839 -1650 871 -1636
rect 777 -1702 792 -1674
rect 918 -1690 930 -1674
tri 918 -1702 930 -1690 ne
rect 1419 -1650 1451 -1636
rect 1357 -1702 1372 -1674
rect 1498 -1690 1510 -1674
tri 1498 -1702 1510 -1690 ne
rect 1999 -1650 2031 -1636
rect 1937 -1702 1952 -1674
rect 2078 -1690 2090 -1674
tri 2078 -1702 2090 -1690 ne
rect 2579 -1650 2611 -1636
rect 2517 -1702 2532 -1674
rect 2658 -1690 2670 -1674
tri 2658 -1702 2670 -1690 ne
rect 3159 -1650 3191 -1636
rect 3097 -1702 3112 -1674
rect 3238 -1690 3250 -1674
tri 3238 -1702 3250 -1690 ne
rect 3739 -1650 3771 -1636
rect 3677 -1702 3692 -1674
rect 3818 -1690 3830 -1674
tri 3818 -1702 3830 -1690 ne
rect 4319 -1650 4351 -1636
rect 4257 -1702 4272 -1674
rect 4398 -1690 4410 -1674
tri 4398 -1702 4410 -1690 ne
rect 4899 -1651 4931 -1637
rect 4837 -1703 4852 -1675
rect 4978 -1691 4990 -1675
tri 4978 -1703 4990 -1691 ne
rect 5479 -1651 5511 -1637
rect 5417 -1703 5432 -1675
rect 5558 -1691 5570 -1675
tri 5558 -1703 5570 -1691 ne
rect 6059 -1651 6091 -1637
rect 5997 -1703 6012 -1675
rect 6138 -1691 6150 -1675
tri 6138 -1703 6150 -1691 ne
rect 6639 -1651 6671 -1637
rect 6577 -1703 6592 -1675
rect 6718 -1691 6730 -1675
tri 6718 -1703 6730 -1691 ne
rect 259 -1920 291 -1906
rect 197 -1972 212 -1944
rect 338 -1960 350 -1944
tri 338 -1972 350 -1960 ne
rect 839 -1920 871 -1906
rect 777 -1972 792 -1944
rect 918 -1960 930 -1944
tri 918 -1972 930 -1960 ne
rect 1419 -1920 1451 -1906
rect 1357 -1972 1372 -1944
rect 1498 -1960 1510 -1944
tri 1498 -1972 1510 -1960 ne
rect 1999 -1920 2031 -1906
rect 1937 -1972 1952 -1944
rect 2078 -1960 2090 -1944
tri 2078 -1972 2090 -1960 ne
rect 2579 -1920 2611 -1906
rect 2517 -1972 2532 -1944
rect 2658 -1960 2670 -1944
tri 2658 -1972 2670 -1960 ne
rect 3159 -1920 3191 -1906
rect 3097 -1972 3112 -1944
rect 3238 -1960 3250 -1944
tri 3238 -1972 3250 -1960 ne
rect 3739 -1920 3771 -1906
rect 3677 -1972 3692 -1944
rect 3818 -1960 3830 -1944
tri 3818 -1972 3830 -1960 ne
rect 4319 -1920 4351 -1906
rect 4257 -1972 4272 -1944
rect 4398 -1960 4410 -1944
tri 4398 -1972 4410 -1960 ne
rect 4899 -1921 4931 -1907
rect 4837 -1973 4852 -1945
rect 4978 -1961 4990 -1945
tri 4978 -1973 4990 -1961 ne
rect 5479 -1921 5511 -1907
rect 5417 -1973 5432 -1945
rect 5558 -1961 5570 -1945
tri 5558 -1973 5570 -1961 ne
rect 6059 -1921 6091 -1907
rect 5997 -1973 6012 -1945
rect 6138 -1961 6150 -1945
tri 6138 -1973 6150 -1961 ne
rect 6639 -1921 6671 -1907
rect 6577 -1973 6592 -1945
rect 6718 -1961 6730 -1945
tri 6718 -1973 6730 -1961 ne
<< psubdiffcont >>
rect 261 1918 289 1920
rect 841 1918 869 1920
rect 1421 1918 1449 1920
rect 2001 1918 2029 1920
rect 2581 1918 2609 1920
rect 3161 1918 3189 1920
rect 3741 1918 3769 1920
rect 4321 1918 4349 1920
rect 4901 1918 4929 1920
rect 5481 1918 5509 1920
rect 6061 1918 6089 1920
rect 6641 1918 6669 1920
rect 261 1648 289 1650
rect 841 1648 869 1650
rect 1421 1648 1449 1650
rect 2001 1648 2029 1650
rect 2581 1648 2609 1650
rect 3161 1648 3189 1650
rect 3741 1648 3769 1650
rect 4321 1648 4349 1650
rect 4901 1648 4929 1650
rect 5481 1648 5509 1650
rect 6061 1648 6089 1650
rect 6641 1648 6669 1650
rect 261 1378 289 1380
rect 841 1378 869 1380
rect 1421 1378 1449 1380
rect 2001 1378 2029 1380
rect 2581 1378 2609 1380
rect 3161 1378 3189 1380
rect 3741 1378 3769 1380
rect 4321 1378 4349 1380
rect 4901 1378 4929 1380
rect 5481 1378 5509 1380
rect 6061 1378 6089 1380
rect 6641 1378 6669 1380
rect 261 1108 289 1110
rect 841 1108 869 1110
rect 1421 1108 1449 1110
rect 2001 1108 2029 1110
rect 2581 1108 2609 1110
rect 3161 1108 3189 1110
rect 3741 1108 3769 1110
rect 4321 1108 4349 1110
rect 4901 1108 4929 1110
rect 5481 1108 5509 1110
rect 6061 1108 6089 1110
rect 6641 1108 6669 1110
rect 261 838 289 840
rect 841 838 869 840
rect 1421 838 1449 840
rect 2001 838 2029 840
rect 2581 838 2609 840
rect 3161 838 3189 840
rect 3741 838 3769 840
rect 4321 838 4349 840
rect 4901 837 4929 839
rect 5481 837 5509 839
rect 6061 837 6089 839
rect 6641 837 6669 839
rect 261 568 289 570
rect 841 568 869 570
rect 1421 568 1449 570
rect 2001 568 2029 570
rect 2581 568 2609 570
rect 3161 568 3189 570
rect 3741 568 3769 570
rect 4321 568 4349 570
rect 4901 567 4929 569
rect 5481 567 5509 569
rect 6061 567 6089 569
rect 6641 567 6669 569
rect 261 298 289 300
rect 841 298 869 300
rect 1421 298 1449 300
rect 2001 298 2029 300
rect 2581 298 2609 300
rect 3161 298 3189 300
rect 3741 298 3769 300
rect 4321 298 4349 300
rect 4901 297 4929 299
rect 5481 297 5509 299
rect 6061 297 6089 299
rect 6641 297 6669 299
rect 261 28 289 30
rect 841 28 869 30
rect 1421 28 1449 30
rect 2001 28 2029 30
rect 2581 28 2609 30
rect 3161 28 3189 30
rect 3741 28 3769 30
rect 4321 28 4349 30
rect 4901 27 4929 29
rect 5481 27 5509 29
rect 6061 27 6089 29
rect 6641 27 6669 29
rect 261 -242 289 -240
rect 841 -242 869 -240
rect 1421 -242 1449 -240
rect 2001 -242 2029 -240
rect 2581 -242 2609 -240
rect 3161 -242 3189 -240
rect 3741 -242 3769 -240
rect 4321 -242 4349 -240
rect 4901 -243 4929 -241
rect 5481 -243 5509 -241
rect 6061 -243 6089 -241
rect 6641 -243 6669 -241
rect 261 -512 289 -510
rect 841 -512 869 -510
rect 1421 -512 1449 -510
rect 2001 -512 2029 -510
rect 2581 -512 2609 -510
rect 3161 -512 3189 -510
rect 3741 -512 3769 -510
rect 4321 -512 4349 -510
rect 4901 -513 4929 -511
rect 5481 -513 5509 -511
rect 6061 -513 6089 -511
rect 6641 -513 6669 -511
rect 261 -782 289 -780
rect 841 -782 869 -780
rect 1421 -782 1449 -780
rect 2001 -782 2029 -780
rect 2581 -782 2609 -780
rect 3161 -782 3189 -780
rect 3741 -782 3769 -780
rect 4321 -782 4349 -780
rect 4901 -783 4929 -781
rect 5481 -783 5509 -781
rect 6061 -783 6089 -781
rect 6641 -783 6669 -781
rect 261 -1052 289 -1050
rect 841 -1052 869 -1050
rect 1421 -1052 1449 -1050
rect 2001 -1052 2029 -1050
rect 2581 -1052 2609 -1050
rect 3161 -1052 3189 -1050
rect 3741 -1052 3769 -1050
rect 4321 -1052 4349 -1050
rect 4901 -1053 4929 -1051
rect 5481 -1053 5509 -1051
rect 6061 -1053 6089 -1051
rect 6641 -1053 6669 -1051
rect 261 -1322 289 -1320
rect 841 -1322 869 -1320
rect 1421 -1322 1449 -1320
rect 2001 -1322 2029 -1320
rect 2581 -1322 2609 -1320
rect 3161 -1322 3189 -1320
rect 3741 -1322 3769 -1320
rect 4321 -1322 4349 -1320
rect 4901 -1323 4929 -1321
rect 5481 -1323 5509 -1321
rect 6061 -1323 6089 -1321
rect 6641 -1323 6669 -1321
rect 261 -1592 289 -1590
rect 841 -1592 869 -1590
rect 1421 -1592 1449 -1590
rect 2001 -1592 2029 -1590
rect 2581 -1592 2609 -1590
rect 3161 -1592 3189 -1590
rect 3741 -1592 3769 -1590
rect 4321 -1592 4349 -1590
rect 4901 -1593 4929 -1591
rect 5481 -1593 5509 -1591
rect 6061 -1593 6089 -1591
rect 6641 -1593 6669 -1591
rect 261 -1862 289 -1860
rect 841 -1862 869 -1860
rect 1421 -1862 1449 -1860
rect 2001 -1862 2029 -1860
rect 2581 -1862 2609 -1860
rect 3161 -1862 3189 -1860
rect 3741 -1862 3769 -1860
rect 4321 -1862 4349 -1860
rect 4901 -1863 4929 -1861
rect 5481 -1863 5509 -1861
rect 6061 -1863 6089 -1861
rect 6641 -1863 6669 -1861
rect 261 -2132 289 -2130
rect 841 -2132 869 -2130
rect 1421 -2132 1449 -2130
rect 2001 -2132 2029 -2130
rect 2581 -2132 2609 -2130
rect 3161 -2132 3189 -2130
rect 3741 -2132 3769 -2130
rect 4321 -2132 4349 -2130
rect 4901 -2133 4929 -2131
rect 5481 -2133 5509 -2131
rect 6061 -2133 6089 -2131
rect 6641 -2133 6669 -2131
<< nsubdiffcont >>
rect 261 2128 289 2130
rect 841 2128 869 2130
rect 1421 2128 1449 2130
rect 2001 2128 2029 2130
rect 2581 2128 2609 2130
rect 3161 2128 3189 2130
rect 3741 2128 3769 2130
rect 4321 2128 4349 2130
rect 4901 2128 4929 2130
rect 5481 2128 5509 2130
rect 6061 2128 6089 2130
rect 6641 2128 6669 2130
rect 261 1858 289 1860
rect 841 1858 869 1860
rect 1421 1858 1449 1860
rect 2001 1858 2029 1860
rect 2581 1858 2609 1860
rect 3161 1858 3189 1860
rect 3741 1858 3769 1860
rect 4321 1858 4349 1860
rect 4901 1858 4929 1860
rect 5481 1858 5509 1860
rect 6061 1858 6089 1860
rect 6641 1858 6669 1860
rect 261 1588 289 1590
rect 841 1588 869 1590
rect 1421 1588 1449 1590
rect 2001 1588 2029 1590
rect 2581 1588 2609 1590
rect 3161 1588 3189 1590
rect 3741 1588 3769 1590
rect 4321 1588 4349 1590
rect 4901 1588 4929 1590
rect 5481 1588 5509 1590
rect 6061 1588 6089 1590
rect 6641 1588 6669 1590
rect 261 1318 289 1320
rect 841 1318 869 1320
rect 1421 1318 1449 1320
rect 2001 1318 2029 1320
rect 2581 1318 2609 1320
rect 3161 1318 3189 1320
rect 3741 1318 3769 1320
rect 4321 1318 4349 1320
rect 4901 1318 4929 1320
rect 5481 1318 5509 1320
rect 6061 1318 6089 1320
rect 6641 1318 6669 1320
rect 261 1048 289 1050
rect 841 1048 869 1050
rect 1421 1048 1449 1050
rect 2001 1048 2029 1050
rect 2581 1048 2609 1050
rect 3161 1048 3189 1050
rect 3741 1048 3769 1050
rect 4321 1048 4349 1050
rect 4901 1047 4929 1049
rect 5481 1047 5509 1049
rect 6061 1047 6089 1049
rect 6641 1047 6669 1049
rect 261 778 289 780
rect 841 778 869 780
rect 1421 778 1449 780
rect 2001 778 2029 780
rect 2581 778 2609 780
rect 3161 778 3189 780
rect 3741 778 3769 780
rect 4321 778 4349 780
rect 4901 777 4929 779
rect 5481 777 5509 779
rect 6061 777 6089 779
rect 6641 777 6669 779
rect 261 508 289 510
rect 841 508 869 510
rect 1421 508 1449 510
rect 2001 508 2029 510
rect 2581 508 2609 510
rect 3161 508 3189 510
rect 3741 508 3769 510
rect 4321 508 4349 510
rect 4901 507 4929 509
rect 5481 507 5509 509
rect 6061 507 6089 509
rect 6641 507 6669 509
rect 261 238 289 240
rect 841 238 869 240
rect 1421 238 1449 240
rect 2001 238 2029 240
rect 2581 238 2609 240
rect 3161 238 3189 240
rect 3741 238 3769 240
rect 4321 238 4349 240
rect 4901 237 4929 239
rect 5481 237 5509 239
rect 6061 237 6089 239
rect 6641 237 6669 239
rect 261 -32 289 -30
rect 841 -32 869 -30
rect 1421 -32 1449 -30
rect 2001 -32 2029 -30
rect 2581 -32 2609 -30
rect 3161 -32 3189 -30
rect 3741 -32 3769 -30
rect 4321 -32 4349 -30
rect 4901 -33 4929 -31
rect 5481 -33 5509 -31
rect 6061 -33 6089 -31
rect 6641 -33 6669 -31
rect 261 -302 289 -300
rect 841 -302 869 -300
rect 1421 -302 1449 -300
rect 2001 -302 2029 -300
rect 2581 -302 2609 -300
rect 3161 -302 3189 -300
rect 3741 -302 3769 -300
rect 4321 -302 4349 -300
rect 4901 -303 4929 -301
rect 5481 -303 5509 -301
rect 6061 -303 6089 -301
rect 6641 -303 6669 -301
rect 261 -572 289 -570
rect 841 -572 869 -570
rect 1421 -572 1449 -570
rect 2001 -572 2029 -570
rect 2581 -572 2609 -570
rect 3161 -572 3189 -570
rect 3741 -572 3769 -570
rect 4321 -572 4349 -570
rect 4901 -573 4929 -571
rect 5481 -573 5509 -571
rect 6061 -573 6089 -571
rect 6641 -573 6669 -571
rect 261 -842 289 -840
rect 841 -842 869 -840
rect 1421 -842 1449 -840
rect 2001 -842 2029 -840
rect 2581 -842 2609 -840
rect 3161 -842 3189 -840
rect 3741 -842 3769 -840
rect 4321 -842 4349 -840
rect 4901 -843 4929 -841
rect 5481 -843 5509 -841
rect 6061 -843 6089 -841
rect 6641 -843 6669 -841
rect 261 -1112 289 -1110
rect 841 -1112 869 -1110
rect 1421 -1112 1449 -1110
rect 2001 -1112 2029 -1110
rect 2581 -1112 2609 -1110
rect 3161 -1112 3189 -1110
rect 3741 -1112 3769 -1110
rect 4321 -1112 4349 -1110
rect 4901 -1113 4929 -1111
rect 5481 -1113 5509 -1111
rect 6061 -1113 6089 -1111
rect 6641 -1113 6669 -1111
rect 261 -1382 289 -1380
rect 841 -1382 869 -1380
rect 1421 -1382 1449 -1380
rect 2001 -1382 2029 -1380
rect 2581 -1382 2609 -1380
rect 3161 -1382 3189 -1380
rect 3741 -1382 3769 -1380
rect 4321 -1382 4349 -1380
rect 4901 -1383 4929 -1381
rect 5481 -1383 5509 -1381
rect 6061 -1383 6089 -1381
rect 6641 -1383 6669 -1381
rect 261 -1652 289 -1650
rect 841 -1652 869 -1650
rect 1421 -1652 1449 -1650
rect 2001 -1652 2029 -1650
rect 2581 -1652 2609 -1650
rect 3161 -1652 3189 -1650
rect 3741 -1652 3769 -1650
rect 4321 -1652 4349 -1650
rect 4901 -1653 4929 -1651
rect 5481 -1653 5509 -1651
rect 6061 -1653 6089 -1651
rect 6641 -1653 6669 -1651
rect 261 -1922 289 -1920
rect 841 -1922 869 -1920
rect 1421 -1922 1449 -1920
rect 2001 -1922 2029 -1920
rect 2581 -1922 2609 -1920
rect 3161 -1922 3189 -1920
rect 3741 -1922 3769 -1920
rect 4321 -1922 4349 -1920
rect 4901 -1923 4929 -1921
rect 5481 -1923 5509 -1921
rect 6061 -1923 6089 -1921
rect 6641 -1923 6669 -1921
<< poly >>
rect -1 2144 6931 2174
rect 106 2116 136 2144
rect 221 2106 251 2128
rect 299 2106 329 2128
rect 414 2116 444 2144
rect 106 2066 136 2088
rect 686 2116 716 2144
rect 801 2106 831 2128
rect 879 2106 909 2128
rect 994 2116 1024 2144
rect 221 2045 251 2078
rect 42 1984 72 2006
rect 128 1984 143 2018
rect 221 1984 251 2011
rect 299 2045 329 2078
rect 414 2066 444 2088
rect 686 2066 716 2088
rect 1266 2116 1296 2144
rect 1381 2106 1411 2128
rect 1459 2106 1489 2128
rect 1574 2116 1604 2144
rect 801 2045 831 2078
rect 299 1984 329 2011
rect 407 1984 422 2018
rect 478 1984 508 2006
rect 622 1984 652 2006
rect 708 1984 723 2018
rect 801 1984 831 2011
rect 879 2045 909 2078
rect 994 2066 1024 2088
rect 1266 2066 1296 2088
rect 1846 2116 1876 2144
rect 1961 2106 1991 2128
rect 2039 2106 2069 2128
rect 2154 2116 2184 2144
rect 1381 2045 1411 2078
rect 879 1984 909 2011
rect 987 1984 1002 2018
rect 1058 1984 1088 2006
rect 1202 1984 1232 2006
rect 1288 1984 1303 2018
rect 1381 1984 1411 2011
rect 1459 2045 1489 2078
rect 1574 2066 1604 2088
rect 1846 2066 1876 2088
rect 2426 2116 2456 2144
rect 2541 2106 2571 2128
rect 2619 2106 2649 2128
rect 2734 2116 2764 2144
rect 1961 2045 1991 2078
rect 1459 1984 1489 2011
rect 1567 1984 1582 2018
rect 1638 1984 1668 2006
rect 1782 1984 1812 2006
rect 1868 1984 1883 2018
rect 1961 1984 1991 2011
rect 2039 2045 2069 2078
rect 2154 2066 2184 2088
rect 2426 2066 2456 2088
rect 3006 2116 3036 2144
rect 3121 2106 3151 2128
rect 3199 2106 3229 2128
rect 3314 2116 3344 2144
rect 2541 2045 2571 2078
rect 2039 1984 2069 2011
rect 2147 1984 2162 2018
rect 2218 1984 2248 2006
rect 2362 1984 2392 2006
rect 2448 1984 2463 2018
rect 2541 1984 2571 2011
rect 2619 2045 2649 2078
rect 2734 2066 2764 2088
rect 3006 2066 3036 2088
rect 3586 2116 3616 2144
rect 3701 2106 3731 2128
rect 3779 2106 3809 2128
rect 3894 2116 3924 2144
rect 3121 2045 3151 2078
rect 2619 1984 2649 2011
rect 2727 1984 2742 2018
rect 2798 1984 2828 2006
rect 2942 1984 2972 2006
rect 3028 1984 3043 2018
rect 3121 1984 3151 2011
rect 3199 2045 3229 2078
rect 3314 2066 3344 2088
rect 3586 2066 3616 2088
rect 4166 2116 4196 2144
rect 4281 2106 4311 2128
rect 4359 2106 4389 2128
rect 4474 2116 4504 2144
rect 3701 2045 3731 2078
rect 3199 1984 3229 2011
rect 3307 1984 3322 2018
rect 3378 1984 3408 2006
rect 3522 1984 3552 2006
rect 3608 1984 3623 2018
rect 3701 1984 3731 2011
rect 3779 2045 3809 2078
rect 3894 2066 3924 2088
rect 4166 2066 4196 2088
rect 4746 2116 4776 2144
rect 4861 2106 4891 2128
rect 4939 2106 4969 2128
rect 5054 2116 5084 2144
rect 4281 2045 4311 2078
rect 3779 1984 3809 2011
rect 3887 1984 3902 2018
rect 3958 1984 3988 2006
rect 4102 1984 4132 2006
rect 4188 1984 4203 2018
rect 4281 1984 4311 2011
rect 4359 2045 4389 2078
rect 4474 2066 4504 2088
rect 4746 2066 4776 2088
rect 5326 2116 5356 2144
rect 5441 2106 5471 2128
rect 5519 2106 5549 2128
rect 5634 2116 5664 2144
rect 4861 2045 4891 2078
rect 4359 1984 4389 2011
rect 4467 1984 4482 2018
rect 4538 1984 4568 2006
rect 4682 1984 4712 2006
rect 4768 1984 4783 2018
rect 4861 1984 4891 2011
rect 4939 2045 4969 2078
rect 5054 2066 5084 2088
rect 5326 2066 5356 2088
rect 5906 2116 5936 2144
rect 6021 2106 6051 2128
rect 6099 2106 6129 2128
rect 6214 2116 6244 2144
rect 5441 2045 5471 2078
rect 4939 1984 4969 2011
rect 5047 1984 5062 2018
rect 5118 1984 5148 2006
rect 5262 1984 5292 2006
rect 5348 1984 5363 2018
rect 5441 1984 5471 2011
rect 5519 2045 5549 2078
rect 5634 2066 5664 2088
rect 5906 2066 5936 2088
rect 6486 2116 6516 2144
rect 6601 2106 6631 2128
rect 6679 2106 6709 2128
rect 6794 2116 6824 2144
rect 6021 2045 6051 2078
rect 5519 1984 5549 2011
rect 5627 1984 5642 2018
rect 5698 1984 5728 2006
rect 5842 1984 5872 2006
rect 5928 1984 5943 2018
rect 6021 1984 6051 2011
rect 6099 2045 6129 2078
rect 6214 2066 6244 2088
rect 6486 2066 6516 2088
rect 6601 2045 6631 2078
rect 6099 1984 6129 2011
rect 6207 1984 6222 2018
rect 6278 1984 6308 2006
rect 6422 1984 6452 2006
rect 6508 1984 6523 2018
rect 6601 1984 6631 2011
rect 6679 2045 6709 2078
rect 6794 2066 6824 2088
rect 6679 1984 6709 2011
rect 6787 1984 6802 2018
rect 6858 1984 6888 2006
rect 128 1970 158 1984
rect 392 1970 422 1984
rect 708 1970 738 1984
rect 972 1970 1002 1984
rect 1288 1970 1318 1984
rect 1552 1970 1582 1984
rect 1868 1970 1898 1984
rect 2132 1970 2162 1984
rect 2448 1970 2478 1984
rect 2712 1970 2742 1984
rect 3028 1970 3058 1984
rect 3292 1970 3322 1984
rect 3608 1970 3638 1984
rect 3872 1970 3902 1984
rect 4188 1970 4218 1984
rect 4452 1970 4482 1984
rect 4768 1970 4798 1984
rect 5032 1970 5062 1984
rect 5348 1970 5378 1984
rect 5612 1970 5642 1984
rect 5928 1970 5958 1984
rect 6192 1970 6222 1984
rect 6508 1970 6538 1984
rect 6772 1970 6802 1984
rect 42 1920 72 1942
rect 128 1920 158 1942
rect 221 1920 251 1942
rect 299 1920 329 1942
rect 392 1920 422 1942
rect 478 1920 508 1942
rect 622 1920 652 1942
rect 708 1920 738 1942
rect 801 1920 831 1942
rect 879 1920 909 1942
rect 972 1920 1002 1942
rect 1058 1920 1088 1942
rect 1202 1920 1232 1942
rect 1288 1920 1318 1942
rect 1381 1920 1411 1942
rect 1459 1920 1489 1942
rect 1552 1920 1582 1942
rect 1638 1920 1668 1942
rect 1782 1920 1812 1942
rect 1868 1920 1898 1942
rect 1961 1920 1991 1942
rect 2039 1920 2069 1942
rect 2132 1920 2162 1942
rect 2218 1920 2248 1942
rect 2362 1920 2392 1942
rect 2448 1920 2478 1942
rect 2541 1920 2571 1942
rect 2619 1920 2649 1942
rect 2712 1920 2742 1942
rect 2798 1920 2828 1942
rect 2942 1920 2972 1942
rect 3028 1920 3058 1942
rect 3121 1920 3151 1942
rect 3199 1920 3229 1942
rect 3292 1920 3322 1942
rect 3378 1920 3408 1942
rect 3522 1920 3552 1942
rect 3608 1920 3638 1942
rect 3701 1920 3731 1942
rect 3779 1920 3809 1942
rect 3872 1920 3902 1942
rect 3958 1920 3988 1942
rect 4102 1920 4132 1942
rect 4188 1920 4218 1942
rect 4281 1920 4311 1942
rect 4359 1920 4389 1942
rect 4452 1920 4482 1942
rect 4538 1920 4568 1942
rect 4682 1920 4712 1942
rect 4768 1920 4798 1942
rect 4861 1920 4891 1942
rect 4939 1920 4969 1942
rect 5032 1920 5062 1942
rect 5118 1920 5148 1942
rect 5262 1920 5292 1942
rect 5348 1920 5378 1942
rect 5441 1920 5471 1942
rect 5519 1920 5549 1942
rect 5612 1920 5642 1942
rect 5698 1920 5728 1942
rect 5842 1920 5872 1942
rect 5928 1920 5958 1942
rect 6021 1920 6051 1942
rect 6099 1920 6129 1942
rect 6192 1920 6222 1942
rect 6278 1920 6308 1942
rect 6422 1920 6452 1942
rect 6508 1920 6538 1942
rect 6601 1920 6631 1942
rect 6679 1920 6709 1942
rect 6772 1920 6802 1942
rect 6858 1920 6888 1942
rect -1 1874 6931 1904
rect 106 1846 136 1874
rect 221 1836 251 1858
rect 299 1836 329 1858
rect 414 1846 444 1874
rect 106 1796 136 1818
rect 686 1846 716 1874
rect 801 1836 831 1858
rect 879 1836 909 1858
rect 994 1846 1024 1874
rect 221 1775 251 1808
rect 42 1714 72 1736
rect 128 1714 143 1748
rect 221 1714 251 1741
rect 299 1775 329 1808
rect 414 1796 444 1818
rect 686 1796 716 1818
rect 1266 1846 1296 1874
rect 1381 1836 1411 1858
rect 1459 1836 1489 1858
rect 1574 1846 1604 1874
rect 801 1775 831 1808
rect 299 1714 329 1741
rect 407 1714 422 1748
rect 478 1714 508 1736
rect 622 1714 652 1736
rect 708 1714 723 1748
rect 801 1714 831 1741
rect 879 1775 909 1808
rect 994 1796 1024 1818
rect 1266 1796 1296 1818
rect 1846 1846 1876 1874
rect 1961 1836 1991 1858
rect 2039 1836 2069 1858
rect 2154 1846 2184 1874
rect 1381 1775 1411 1808
rect 879 1714 909 1741
rect 987 1714 1002 1748
rect 1058 1714 1088 1736
rect 1202 1714 1232 1736
rect 1288 1714 1303 1748
rect 1381 1714 1411 1741
rect 1459 1775 1489 1808
rect 1574 1796 1604 1818
rect 1846 1796 1876 1818
rect 2426 1846 2456 1874
rect 2541 1836 2571 1858
rect 2619 1836 2649 1858
rect 2734 1846 2764 1874
rect 1961 1775 1991 1808
rect 1459 1714 1489 1741
rect 1567 1714 1582 1748
rect 1638 1714 1668 1736
rect 1782 1714 1812 1736
rect 1868 1714 1883 1748
rect 1961 1714 1991 1741
rect 2039 1775 2069 1808
rect 2154 1796 2184 1818
rect 2426 1796 2456 1818
rect 3006 1846 3036 1874
rect 3121 1836 3151 1858
rect 3199 1836 3229 1858
rect 3314 1846 3344 1874
rect 2541 1775 2571 1808
rect 2039 1714 2069 1741
rect 2147 1714 2162 1748
rect 2218 1714 2248 1736
rect 2362 1714 2392 1736
rect 2448 1714 2463 1748
rect 2541 1714 2571 1741
rect 2619 1775 2649 1808
rect 2734 1796 2764 1818
rect 3006 1796 3036 1818
rect 3586 1846 3616 1874
rect 3701 1836 3731 1858
rect 3779 1836 3809 1858
rect 3894 1846 3924 1874
rect 3121 1775 3151 1808
rect 2619 1714 2649 1741
rect 2727 1714 2742 1748
rect 2798 1714 2828 1736
rect 2942 1714 2972 1736
rect 3028 1714 3043 1748
rect 3121 1714 3151 1741
rect 3199 1775 3229 1808
rect 3314 1796 3344 1818
rect 3586 1796 3616 1818
rect 4166 1846 4196 1874
rect 4281 1836 4311 1858
rect 4359 1836 4389 1858
rect 4474 1846 4504 1874
rect 3701 1775 3731 1808
rect 3199 1714 3229 1741
rect 3307 1714 3322 1748
rect 3378 1714 3408 1736
rect 3522 1714 3552 1736
rect 3608 1714 3623 1748
rect 3701 1714 3731 1741
rect 3779 1775 3809 1808
rect 3894 1796 3924 1818
rect 4166 1796 4196 1818
rect 4746 1846 4776 1874
rect 4861 1836 4891 1858
rect 4939 1836 4969 1858
rect 5054 1846 5084 1874
rect 4281 1775 4311 1808
rect 3779 1714 3809 1741
rect 3887 1714 3902 1748
rect 3958 1714 3988 1736
rect 4102 1714 4132 1736
rect 4188 1714 4203 1748
rect 4281 1714 4311 1741
rect 4359 1775 4389 1808
rect 4474 1796 4504 1818
rect 4746 1796 4776 1818
rect 5326 1846 5356 1874
rect 5441 1836 5471 1858
rect 5519 1836 5549 1858
rect 5634 1846 5664 1874
rect 4861 1775 4891 1808
rect 4359 1714 4389 1741
rect 4467 1714 4482 1748
rect 4538 1714 4568 1736
rect 4682 1714 4712 1736
rect 4768 1714 4783 1748
rect 4861 1714 4891 1741
rect 4939 1775 4969 1808
rect 5054 1796 5084 1818
rect 5326 1796 5356 1818
rect 5906 1846 5936 1874
rect 6021 1836 6051 1858
rect 6099 1836 6129 1858
rect 6214 1846 6244 1874
rect 5441 1775 5471 1808
rect 4939 1714 4969 1741
rect 5047 1714 5062 1748
rect 5118 1714 5148 1736
rect 5262 1714 5292 1736
rect 5348 1714 5363 1748
rect 5441 1714 5471 1741
rect 5519 1775 5549 1808
rect 5634 1796 5664 1818
rect 5906 1796 5936 1818
rect 6486 1846 6516 1874
rect 6601 1836 6631 1858
rect 6679 1836 6709 1858
rect 6794 1846 6824 1874
rect 6021 1775 6051 1808
rect 5519 1714 5549 1741
rect 5627 1714 5642 1748
rect 5698 1714 5728 1736
rect 5842 1714 5872 1736
rect 5928 1714 5943 1748
rect 6021 1714 6051 1741
rect 6099 1775 6129 1808
rect 6214 1796 6244 1818
rect 6486 1796 6516 1818
rect 6601 1775 6631 1808
rect 6099 1714 6129 1741
rect 6207 1714 6222 1748
rect 6278 1714 6308 1736
rect 6422 1714 6452 1736
rect 6508 1714 6523 1748
rect 6601 1714 6631 1741
rect 6679 1775 6709 1808
rect 6794 1796 6824 1818
rect 6679 1714 6709 1741
rect 6787 1714 6802 1748
rect 6858 1714 6888 1736
rect 128 1700 158 1714
rect 392 1700 422 1714
rect 708 1700 738 1714
rect 972 1700 1002 1714
rect 1288 1700 1318 1714
rect 1552 1700 1582 1714
rect 1868 1700 1898 1714
rect 2132 1700 2162 1714
rect 2448 1700 2478 1714
rect 2712 1700 2742 1714
rect 3028 1700 3058 1714
rect 3292 1700 3322 1714
rect 3608 1700 3638 1714
rect 3872 1700 3902 1714
rect 4188 1700 4218 1714
rect 4452 1700 4482 1714
rect 4768 1700 4798 1714
rect 5032 1700 5062 1714
rect 5348 1700 5378 1714
rect 5612 1700 5642 1714
rect 5928 1700 5958 1714
rect 6192 1700 6222 1714
rect 6508 1700 6538 1714
rect 6772 1700 6802 1714
rect 42 1650 72 1672
rect 128 1650 158 1672
rect 221 1650 251 1672
rect 299 1650 329 1672
rect 392 1650 422 1672
rect 478 1650 508 1672
rect 622 1650 652 1672
rect 708 1650 738 1672
rect 801 1650 831 1672
rect 879 1650 909 1672
rect 972 1650 1002 1672
rect 1058 1650 1088 1672
rect 1202 1650 1232 1672
rect 1288 1650 1318 1672
rect 1381 1650 1411 1672
rect 1459 1650 1489 1672
rect 1552 1650 1582 1672
rect 1638 1650 1668 1672
rect 1782 1650 1812 1672
rect 1868 1650 1898 1672
rect 1961 1650 1991 1672
rect 2039 1650 2069 1672
rect 2132 1650 2162 1672
rect 2218 1650 2248 1672
rect 2362 1650 2392 1672
rect 2448 1650 2478 1672
rect 2541 1650 2571 1672
rect 2619 1650 2649 1672
rect 2712 1650 2742 1672
rect 2798 1650 2828 1672
rect 2942 1650 2972 1672
rect 3028 1650 3058 1672
rect 3121 1650 3151 1672
rect 3199 1650 3229 1672
rect 3292 1650 3322 1672
rect 3378 1650 3408 1672
rect 3522 1650 3552 1672
rect 3608 1650 3638 1672
rect 3701 1650 3731 1672
rect 3779 1650 3809 1672
rect 3872 1650 3902 1672
rect 3958 1650 3988 1672
rect 4102 1650 4132 1672
rect 4188 1650 4218 1672
rect 4281 1650 4311 1672
rect 4359 1650 4389 1672
rect 4452 1650 4482 1672
rect 4538 1650 4568 1672
rect 4682 1650 4712 1672
rect 4768 1650 4798 1672
rect 4861 1650 4891 1672
rect 4939 1650 4969 1672
rect 5032 1650 5062 1672
rect 5118 1650 5148 1672
rect 5262 1650 5292 1672
rect 5348 1650 5378 1672
rect 5441 1650 5471 1672
rect 5519 1650 5549 1672
rect 5612 1650 5642 1672
rect 5698 1650 5728 1672
rect 5842 1650 5872 1672
rect 5928 1650 5958 1672
rect 6021 1650 6051 1672
rect 6099 1650 6129 1672
rect 6192 1650 6222 1672
rect 6278 1650 6308 1672
rect 6422 1650 6452 1672
rect 6508 1650 6538 1672
rect 6601 1650 6631 1672
rect 6679 1650 6709 1672
rect 6772 1650 6802 1672
rect 6858 1650 6888 1672
rect -1 1604 6931 1634
rect 106 1576 136 1604
rect 221 1566 251 1588
rect 299 1566 329 1588
rect 414 1576 444 1604
rect 106 1526 136 1548
rect 686 1576 716 1604
rect 801 1566 831 1588
rect 879 1566 909 1588
rect 994 1576 1024 1604
rect 221 1505 251 1538
rect 42 1444 72 1466
rect 128 1444 143 1478
rect 221 1444 251 1471
rect 299 1505 329 1538
rect 414 1526 444 1548
rect 686 1526 716 1548
rect 1266 1576 1296 1604
rect 1381 1566 1411 1588
rect 1459 1566 1489 1588
rect 1574 1576 1604 1604
rect 801 1505 831 1538
rect 299 1444 329 1471
rect 407 1444 422 1478
rect 478 1444 508 1466
rect 622 1444 652 1466
rect 708 1444 723 1478
rect 801 1444 831 1471
rect 879 1505 909 1538
rect 994 1526 1024 1548
rect 1266 1526 1296 1548
rect 1846 1576 1876 1604
rect 1961 1566 1991 1588
rect 2039 1566 2069 1588
rect 2154 1576 2184 1604
rect 1381 1505 1411 1538
rect 879 1444 909 1471
rect 987 1444 1002 1478
rect 1058 1444 1088 1466
rect 1202 1444 1232 1466
rect 1288 1444 1303 1478
rect 1381 1444 1411 1471
rect 1459 1505 1489 1538
rect 1574 1526 1604 1548
rect 1846 1526 1876 1548
rect 2426 1576 2456 1604
rect 2541 1566 2571 1588
rect 2619 1566 2649 1588
rect 2734 1576 2764 1604
rect 1961 1505 1991 1538
rect 1459 1444 1489 1471
rect 1567 1444 1582 1478
rect 1638 1444 1668 1466
rect 1782 1444 1812 1466
rect 1868 1444 1883 1478
rect 1961 1444 1991 1471
rect 2039 1505 2069 1538
rect 2154 1526 2184 1548
rect 2426 1526 2456 1548
rect 3006 1576 3036 1604
rect 3121 1566 3151 1588
rect 3199 1566 3229 1588
rect 3314 1576 3344 1604
rect 2541 1505 2571 1538
rect 2039 1444 2069 1471
rect 2147 1444 2162 1478
rect 2218 1444 2248 1466
rect 2362 1444 2392 1466
rect 2448 1444 2463 1478
rect 2541 1444 2571 1471
rect 2619 1505 2649 1538
rect 2734 1526 2764 1548
rect 3006 1526 3036 1548
rect 3586 1576 3616 1604
rect 3701 1566 3731 1588
rect 3779 1566 3809 1588
rect 3894 1576 3924 1604
rect 3121 1505 3151 1538
rect 2619 1444 2649 1471
rect 2727 1444 2742 1478
rect 2798 1444 2828 1466
rect 2942 1444 2972 1466
rect 3028 1444 3043 1478
rect 3121 1444 3151 1471
rect 3199 1505 3229 1538
rect 3314 1526 3344 1548
rect 3586 1526 3616 1548
rect 4166 1576 4196 1604
rect 4281 1566 4311 1588
rect 4359 1566 4389 1588
rect 4474 1576 4504 1604
rect 3701 1505 3731 1538
rect 3199 1444 3229 1471
rect 3307 1444 3322 1478
rect 3378 1444 3408 1466
rect 3522 1444 3552 1466
rect 3608 1444 3623 1478
rect 3701 1444 3731 1471
rect 3779 1505 3809 1538
rect 3894 1526 3924 1548
rect 4166 1526 4196 1548
rect 4746 1576 4776 1604
rect 4861 1566 4891 1588
rect 4939 1566 4969 1588
rect 5054 1576 5084 1604
rect 4281 1505 4311 1538
rect 3779 1444 3809 1471
rect 3887 1444 3902 1478
rect 3958 1444 3988 1466
rect 4102 1444 4132 1466
rect 4188 1444 4203 1478
rect 4281 1444 4311 1471
rect 4359 1505 4389 1538
rect 4474 1526 4504 1548
rect 4746 1526 4776 1548
rect 5326 1576 5356 1604
rect 5441 1566 5471 1588
rect 5519 1566 5549 1588
rect 5634 1576 5664 1604
rect 4861 1505 4891 1538
rect 4359 1444 4389 1471
rect 4467 1444 4482 1478
rect 4538 1444 4568 1466
rect 4682 1444 4712 1466
rect 4768 1444 4783 1478
rect 4861 1444 4891 1471
rect 4939 1505 4969 1538
rect 5054 1526 5084 1548
rect 5326 1526 5356 1548
rect 5906 1576 5936 1604
rect 6021 1566 6051 1588
rect 6099 1566 6129 1588
rect 6214 1576 6244 1604
rect 5441 1505 5471 1538
rect 4939 1444 4969 1471
rect 5047 1444 5062 1478
rect 5118 1444 5148 1466
rect 5262 1444 5292 1466
rect 5348 1444 5363 1478
rect 5441 1444 5471 1471
rect 5519 1505 5549 1538
rect 5634 1526 5664 1548
rect 5906 1526 5936 1548
rect 6486 1576 6516 1604
rect 6601 1566 6631 1588
rect 6679 1566 6709 1588
rect 6794 1576 6824 1604
rect 6021 1505 6051 1538
rect 5519 1444 5549 1471
rect 5627 1444 5642 1478
rect 5698 1444 5728 1466
rect 5842 1444 5872 1466
rect 5928 1444 5943 1478
rect 6021 1444 6051 1471
rect 6099 1505 6129 1538
rect 6214 1526 6244 1548
rect 6486 1526 6516 1548
rect 6601 1505 6631 1538
rect 6099 1444 6129 1471
rect 6207 1444 6222 1478
rect 6278 1444 6308 1466
rect 6422 1444 6452 1466
rect 6508 1444 6523 1478
rect 6601 1444 6631 1471
rect 6679 1505 6709 1538
rect 6794 1526 6824 1548
rect 6679 1444 6709 1471
rect 6787 1444 6802 1478
rect 6858 1444 6888 1466
rect 128 1430 158 1444
rect 392 1430 422 1444
rect 708 1430 738 1444
rect 972 1430 1002 1444
rect 1288 1430 1318 1444
rect 1552 1430 1582 1444
rect 1868 1430 1898 1444
rect 2132 1430 2162 1444
rect 2448 1430 2478 1444
rect 2712 1430 2742 1444
rect 3028 1430 3058 1444
rect 3292 1430 3322 1444
rect 3608 1430 3638 1444
rect 3872 1430 3902 1444
rect 4188 1430 4218 1444
rect 4452 1430 4482 1444
rect 4768 1430 4798 1444
rect 5032 1430 5062 1444
rect 5348 1430 5378 1444
rect 5612 1430 5642 1444
rect 5928 1430 5958 1444
rect 6192 1430 6222 1444
rect 6508 1430 6538 1444
rect 6772 1430 6802 1444
rect 42 1380 72 1402
rect 128 1380 158 1402
rect 221 1380 251 1402
rect 299 1380 329 1402
rect 392 1380 422 1402
rect 478 1380 508 1402
rect 622 1380 652 1402
rect 708 1380 738 1402
rect 801 1380 831 1402
rect 879 1380 909 1402
rect 972 1380 1002 1402
rect 1058 1380 1088 1402
rect 1202 1380 1232 1402
rect 1288 1380 1318 1402
rect 1381 1380 1411 1402
rect 1459 1380 1489 1402
rect 1552 1380 1582 1402
rect 1638 1380 1668 1402
rect 1782 1380 1812 1402
rect 1868 1380 1898 1402
rect 1961 1380 1991 1402
rect 2039 1380 2069 1402
rect 2132 1380 2162 1402
rect 2218 1380 2248 1402
rect 2362 1380 2392 1402
rect 2448 1380 2478 1402
rect 2541 1380 2571 1402
rect 2619 1380 2649 1402
rect 2712 1380 2742 1402
rect 2798 1380 2828 1402
rect 2942 1380 2972 1402
rect 3028 1380 3058 1402
rect 3121 1380 3151 1402
rect 3199 1380 3229 1402
rect 3292 1380 3322 1402
rect 3378 1380 3408 1402
rect 3522 1380 3552 1402
rect 3608 1380 3638 1402
rect 3701 1380 3731 1402
rect 3779 1380 3809 1402
rect 3872 1380 3902 1402
rect 3958 1380 3988 1402
rect 4102 1380 4132 1402
rect 4188 1380 4218 1402
rect 4281 1380 4311 1402
rect 4359 1380 4389 1402
rect 4452 1380 4482 1402
rect 4538 1380 4568 1402
rect 4682 1380 4712 1402
rect 4768 1380 4798 1402
rect 4861 1380 4891 1402
rect 4939 1380 4969 1402
rect 5032 1380 5062 1402
rect 5118 1380 5148 1402
rect 5262 1380 5292 1402
rect 5348 1380 5378 1402
rect 5441 1380 5471 1402
rect 5519 1380 5549 1402
rect 5612 1380 5642 1402
rect 5698 1380 5728 1402
rect 5842 1380 5872 1402
rect 5928 1380 5958 1402
rect 6021 1380 6051 1402
rect 6099 1380 6129 1402
rect 6192 1380 6222 1402
rect 6278 1380 6308 1402
rect 6422 1380 6452 1402
rect 6508 1380 6538 1402
rect 6601 1380 6631 1402
rect 6679 1380 6709 1402
rect 6772 1380 6802 1402
rect 6858 1380 6888 1402
rect -1 1334 6931 1364
rect 106 1306 136 1334
rect 221 1296 251 1318
rect 299 1296 329 1318
rect 414 1306 444 1334
rect 106 1256 136 1278
rect 686 1306 716 1334
rect 801 1296 831 1318
rect 879 1296 909 1318
rect 994 1306 1024 1334
rect 221 1235 251 1268
rect 42 1174 72 1196
rect 128 1174 143 1208
rect 221 1174 251 1201
rect 299 1235 329 1268
rect 414 1256 444 1278
rect 686 1256 716 1278
rect 1266 1306 1296 1334
rect 1381 1296 1411 1318
rect 1459 1296 1489 1318
rect 1574 1306 1604 1334
rect 801 1235 831 1268
rect 299 1174 329 1201
rect 407 1174 422 1208
rect 478 1174 508 1196
rect 622 1174 652 1196
rect 708 1174 723 1208
rect 801 1174 831 1201
rect 879 1235 909 1268
rect 994 1256 1024 1278
rect 1266 1256 1296 1278
rect 1846 1306 1876 1334
rect 1961 1296 1991 1318
rect 2039 1296 2069 1318
rect 2154 1306 2184 1334
rect 1381 1235 1411 1268
rect 879 1174 909 1201
rect 987 1174 1002 1208
rect 1058 1174 1088 1196
rect 1202 1174 1232 1196
rect 1288 1174 1303 1208
rect 1381 1174 1411 1201
rect 1459 1235 1489 1268
rect 1574 1256 1604 1278
rect 1846 1256 1876 1278
rect 2426 1306 2456 1334
rect 2541 1296 2571 1318
rect 2619 1296 2649 1318
rect 2734 1306 2764 1334
rect 1961 1235 1991 1268
rect 1459 1174 1489 1201
rect 1567 1174 1582 1208
rect 1638 1174 1668 1196
rect 1782 1174 1812 1196
rect 1868 1174 1883 1208
rect 1961 1174 1991 1201
rect 2039 1235 2069 1268
rect 2154 1256 2184 1278
rect 2426 1256 2456 1278
rect 3006 1306 3036 1334
rect 3121 1296 3151 1318
rect 3199 1296 3229 1318
rect 3314 1306 3344 1334
rect 2541 1235 2571 1268
rect 2039 1174 2069 1201
rect 2147 1174 2162 1208
rect 2218 1174 2248 1196
rect 2362 1174 2392 1196
rect 2448 1174 2463 1208
rect 2541 1174 2571 1201
rect 2619 1235 2649 1268
rect 2734 1256 2764 1278
rect 3006 1256 3036 1278
rect 3586 1306 3616 1334
rect 3701 1296 3731 1318
rect 3779 1296 3809 1318
rect 3894 1306 3924 1334
rect 3121 1235 3151 1268
rect 2619 1174 2649 1201
rect 2727 1174 2742 1208
rect 2798 1174 2828 1196
rect 2942 1174 2972 1196
rect 3028 1174 3043 1208
rect 3121 1174 3151 1201
rect 3199 1235 3229 1268
rect 3314 1256 3344 1278
rect 3586 1256 3616 1278
rect 4166 1306 4196 1334
rect 4281 1296 4311 1318
rect 4359 1296 4389 1318
rect 4474 1306 4504 1334
rect 3701 1235 3731 1268
rect 3199 1174 3229 1201
rect 3307 1174 3322 1208
rect 3378 1174 3408 1196
rect 3522 1174 3552 1196
rect 3608 1174 3623 1208
rect 3701 1174 3731 1201
rect 3779 1235 3809 1268
rect 3894 1256 3924 1278
rect 4166 1256 4196 1278
rect 4746 1306 4776 1334
rect 4861 1296 4891 1318
rect 4939 1296 4969 1318
rect 5054 1306 5084 1334
rect 4281 1235 4311 1268
rect 3779 1174 3809 1201
rect 3887 1174 3902 1208
rect 3958 1174 3988 1196
rect 4102 1174 4132 1196
rect 4188 1174 4203 1208
rect 4281 1174 4311 1201
rect 4359 1235 4389 1268
rect 4474 1256 4504 1278
rect 4746 1256 4776 1278
rect 5326 1306 5356 1334
rect 5441 1296 5471 1318
rect 5519 1296 5549 1318
rect 5634 1306 5664 1334
rect 4861 1235 4891 1268
rect 4359 1174 4389 1201
rect 4467 1174 4482 1208
rect 4538 1174 4568 1196
rect 4682 1174 4712 1196
rect 4768 1174 4783 1208
rect 4861 1174 4891 1201
rect 4939 1235 4969 1268
rect 5054 1256 5084 1278
rect 5326 1256 5356 1278
rect 5906 1306 5936 1334
rect 6021 1296 6051 1318
rect 6099 1296 6129 1318
rect 6214 1306 6244 1334
rect 5441 1235 5471 1268
rect 4939 1174 4969 1201
rect 5047 1174 5062 1208
rect 5118 1174 5148 1196
rect 5262 1174 5292 1196
rect 5348 1174 5363 1208
rect 5441 1174 5471 1201
rect 5519 1235 5549 1268
rect 5634 1256 5664 1278
rect 5906 1256 5936 1278
rect 6486 1306 6516 1334
rect 6601 1296 6631 1318
rect 6679 1296 6709 1318
rect 6794 1306 6824 1334
rect 6021 1235 6051 1268
rect 5519 1174 5549 1201
rect 5627 1174 5642 1208
rect 5698 1174 5728 1196
rect 5842 1174 5872 1196
rect 5928 1174 5943 1208
rect 6021 1174 6051 1201
rect 6099 1235 6129 1268
rect 6214 1256 6244 1278
rect 6486 1256 6516 1278
rect 6601 1235 6631 1268
rect 6099 1174 6129 1201
rect 6207 1174 6222 1208
rect 6278 1174 6308 1196
rect 6422 1174 6452 1196
rect 6508 1174 6523 1208
rect 6601 1174 6631 1201
rect 6679 1235 6709 1268
rect 6794 1256 6824 1278
rect 6679 1174 6709 1201
rect 6787 1174 6802 1208
rect 6858 1174 6888 1196
rect 128 1160 158 1174
rect 392 1160 422 1174
rect 708 1160 738 1174
rect 972 1160 1002 1174
rect 1288 1160 1318 1174
rect 1552 1160 1582 1174
rect 1868 1160 1898 1174
rect 2132 1160 2162 1174
rect 2448 1160 2478 1174
rect 2712 1160 2742 1174
rect 3028 1160 3058 1174
rect 3292 1160 3322 1174
rect 3608 1160 3638 1174
rect 3872 1160 3902 1174
rect 4188 1160 4218 1174
rect 4452 1160 4482 1174
rect 4768 1160 4798 1174
rect 5032 1160 5062 1174
rect 5348 1160 5378 1174
rect 5612 1160 5642 1174
rect 5928 1160 5958 1174
rect 6192 1160 6222 1174
rect 6508 1160 6538 1174
rect 6772 1160 6802 1174
rect 42 1110 72 1132
rect 128 1110 158 1132
rect 221 1110 251 1132
rect 299 1110 329 1132
rect 392 1110 422 1132
rect 478 1110 508 1132
rect 622 1110 652 1132
rect 708 1110 738 1132
rect 801 1110 831 1132
rect 879 1110 909 1132
rect 972 1110 1002 1132
rect 1058 1110 1088 1132
rect 1202 1110 1232 1132
rect 1288 1110 1318 1132
rect 1381 1110 1411 1132
rect 1459 1110 1489 1132
rect 1552 1110 1582 1132
rect 1638 1110 1668 1132
rect 1782 1110 1812 1132
rect 1868 1110 1898 1132
rect 1961 1110 1991 1132
rect 2039 1110 2069 1132
rect 2132 1110 2162 1132
rect 2218 1110 2248 1132
rect 2362 1110 2392 1132
rect 2448 1110 2478 1132
rect 2541 1110 2571 1132
rect 2619 1110 2649 1132
rect 2712 1110 2742 1132
rect 2798 1110 2828 1132
rect 2942 1110 2972 1132
rect 3028 1110 3058 1132
rect 3121 1110 3151 1132
rect 3199 1110 3229 1132
rect 3292 1110 3322 1132
rect 3378 1110 3408 1132
rect 3522 1110 3552 1132
rect 3608 1110 3638 1132
rect 3701 1110 3731 1132
rect 3779 1110 3809 1132
rect 3872 1110 3902 1132
rect 3958 1110 3988 1132
rect 4102 1110 4132 1132
rect 4188 1110 4218 1132
rect 4281 1110 4311 1132
rect 4359 1110 4389 1132
rect 4452 1110 4482 1132
rect 4538 1110 4568 1132
rect 4682 1110 4712 1132
rect 4768 1110 4798 1132
rect 4861 1110 4891 1132
rect 4939 1110 4969 1132
rect 5032 1110 5062 1132
rect 5118 1110 5148 1132
rect 5262 1110 5292 1132
rect 5348 1110 5378 1132
rect 5441 1110 5471 1132
rect 5519 1110 5549 1132
rect 5612 1110 5642 1132
rect 5698 1110 5728 1132
rect 5842 1110 5872 1132
rect 5928 1110 5958 1132
rect 6021 1110 6051 1132
rect 6099 1110 6129 1132
rect 6192 1110 6222 1132
rect 6278 1110 6308 1132
rect 6422 1110 6452 1132
rect 6508 1110 6538 1132
rect 6601 1110 6631 1132
rect 6679 1110 6709 1132
rect 6772 1110 6802 1132
rect 6858 1110 6888 1132
rect -1 1093 4611 1094
rect -1 1064 6931 1093
rect 106 1036 136 1064
rect 221 1026 251 1048
rect 299 1026 329 1048
rect 414 1036 444 1064
rect 106 986 136 1008
rect 686 1036 716 1064
rect 801 1026 831 1048
rect 879 1026 909 1048
rect 994 1036 1024 1064
rect 221 965 251 998
rect 42 904 72 926
rect 128 904 143 938
rect 221 904 251 931
rect 299 965 329 998
rect 414 986 444 1008
rect 686 986 716 1008
rect 1266 1036 1296 1064
rect 1381 1026 1411 1048
rect 1459 1026 1489 1048
rect 1574 1036 1604 1064
rect 801 965 831 998
rect 299 904 329 931
rect 407 904 422 938
rect 478 904 508 926
rect 622 904 652 926
rect 708 904 723 938
rect 801 904 831 931
rect 879 965 909 998
rect 994 986 1024 1008
rect 1266 986 1296 1008
rect 1846 1036 1876 1064
rect 1961 1026 1991 1048
rect 2039 1026 2069 1048
rect 2154 1036 2184 1064
rect 1381 965 1411 998
rect 879 904 909 931
rect 987 904 1002 938
rect 1058 904 1088 926
rect 1202 904 1232 926
rect 1288 904 1303 938
rect 1381 904 1411 931
rect 1459 965 1489 998
rect 1574 986 1604 1008
rect 1846 986 1876 1008
rect 2426 1036 2456 1064
rect 2541 1026 2571 1048
rect 2619 1026 2649 1048
rect 2734 1036 2764 1064
rect 1961 965 1991 998
rect 1459 904 1489 931
rect 1567 904 1582 938
rect 1638 904 1668 926
rect 1782 904 1812 926
rect 1868 904 1883 938
rect 1961 904 1991 931
rect 2039 965 2069 998
rect 2154 986 2184 1008
rect 2426 986 2456 1008
rect 3006 1036 3036 1064
rect 3121 1026 3151 1048
rect 3199 1026 3229 1048
rect 3314 1036 3344 1064
rect 2541 965 2571 998
rect 2039 904 2069 931
rect 2147 904 2162 938
rect 2218 904 2248 926
rect 2362 904 2392 926
rect 2448 904 2463 938
rect 2541 904 2571 931
rect 2619 965 2649 998
rect 2734 986 2764 1008
rect 3006 986 3036 1008
rect 3586 1036 3616 1064
rect 3701 1026 3731 1048
rect 3779 1026 3809 1048
rect 3894 1036 3924 1064
rect 3121 965 3151 998
rect 2619 904 2649 931
rect 2727 904 2742 938
rect 2798 904 2828 926
rect 2942 904 2972 926
rect 3028 904 3043 938
rect 3121 904 3151 931
rect 3199 965 3229 998
rect 3314 986 3344 1008
rect 3586 986 3616 1008
rect 4166 1036 4196 1064
rect 4281 1026 4311 1048
rect 4359 1026 4389 1048
rect 4474 1036 4504 1064
rect 4591 1063 6931 1064
rect 3701 965 3731 998
rect 3199 904 3229 931
rect 3307 904 3322 938
rect 3378 904 3408 926
rect 3522 904 3552 926
rect 3608 904 3623 938
rect 3701 904 3731 931
rect 3779 965 3809 998
rect 3894 986 3924 1008
rect 4166 986 4196 1008
rect 4746 1035 4776 1063
rect 4281 965 4311 998
rect 3779 904 3809 931
rect 3887 904 3902 938
rect 3958 904 3988 926
rect 4102 904 4132 926
rect 4188 904 4203 938
rect 4281 904 4311 931
rect 4359 965 4389 998
rect 4474 986 4504 1008
rect 4861 1025 4891 1047
rect 4939 1025 4969 1047
rect 5054 1035 5084 1063
rect 4746 985 4776 1007
rect 5326 1035 5356 1063
rect 5441 1025 5471 1047
rect 5519 1025 5549 1047
rect 5634 1035 5664 1063
rect 4861 964 4891 997
rect 4359 904 4389 931
rect 4467 904 4482 938
rect 4538 904 4568 926
rect 128 890 158 904
rect 392 890 422 904
rect 708 890 738 904
rect 972 890 1002 904
rect 1288 890 1318 904
rect 1552 890 1582 904
rect 1868 890 1898 904
rect 2132 890 2162 904
rect 2448 890 2478 904
rect 2712 890 2742 904
rect 3028 890 3058 904
rect 3292 890 3322 904
rect 3608 890 3638 904
rect 3872 890 3902 904
rect 4188 890 4218 904
rect 4452 890 4482 904
rect 4682 903 4712 925
rect 4768 903 4783 937
rect 4861 903 4891 930
rect 4939 964 4969 997
rect 5054 985 5084 1007
rect 5326 985 5356 1007
rect 5906 1035 5936 1063
rect 6021 1025 6051 1047
rect 6099 1025 6129 1047
rect 6214 1035 6244 1063
rect 5441 964 5471 997
rect 4939 903 4969 930
rect 5047 903 5062 937
rect 5118 903 5148 925
rect 5262 903 5292 925
rect 5348 903 5363 937
rect 5441 903 5471 930
rect 5519 964 5549 997
rect 5634 985 5664 1007
rect 5906 985 5936 1007
rect 6486 1035 6516 1063
rect 6601 1025 6631 1047
rect 6679 1025 6709 1047
rect 6794 1035 6824 1063
rect 6021 964 6051 997
rect 5519 903 5549 930
rect 5627 903 5642 937
rect 5698 903 5728 925
rect 5842 903 5872 925
rect 5928 903 5943 937
rect 6021 903 6051 930
rect 6099 964 6129 997
rect 6214 985 6244 1007
rect 6486 985 6516 1007
rect 6601 964 6631 997
rect 6099 903 6129 930
rect 6207 903 6222 937
rect 6278 903 6308 925
rect 6422 903 6452 925
rect 6508 903 6523 937
rect 6601 903 6631 930
rect 6679 964 6709 997
rect 6794 985 6824 1007
rect 6679 903 6709 930
rect 6787 903 6802 937
rect 6858 903 6888 925
rect 42 840 72 862
rect 128 840 158 862
rect 221 840 251 862
rect 299 840 329 862
rect 392 840 422 862
rect 478 840 508 862
rect 622 840 652 862
rect 708 840 738 862
rect 801 840 831 862
rect 879 840 909 862
rect 972 840 1002 862
rect 1058 840 1088 862
rect 1202 840 1232 862
rect 1288 840 1318 862
rect 1381 840 1411 862
rect 1459 840 1489 862
rect 1552 840 1582 862
rect 1638 840 1668 862
rect 1782 840 1812 862
rect 1868 840 1898 862
rect 1961 840 1991 862
rect 2039 840 2069 862
rect 2132 840 2162 862
rect 2218 840 2248 862
rect 2362 840 2392 862
rect 2448 840 2478 862
rect 2541 840 2571 862
rect 2619 840 2649 862
rect 2712 840 2742 862
rect 2798 840 2828 862
rect 2942 840 2972 862
rect 3028 840 3058 862
rect 3121 840 3151 862
rect 3199 840 3229 862
rect 3292 840 3322 862
rect 3378 840 3408 862
rect 3522 840 3552 862
rect 3608 840 3638 862
rect 3701 840 3731 862
rect 3779 840 3809 862
rect 3872 840 3902 862
rect 3958 840 3988 862
rect 4102 840 4132 862
rect 4188 840 4218 862
rect 4281 840 4311 862
rect 4359 840 4389 862
rect 4452 840 4482 862
rect 4538 840 4568 862
rect 4768 889 4798 903
rect 5032 889 5062 903
rect 5348 889 5378 903
rect 5612 889 5642 903
rect 5928 889 5958 903
rect 6192 889 6222 903
rect 6508 889 6538 903
rect 6772 889 6802 903
rect 4682 839 4712 861
rect 4768 839 4798 861
rect 4861 839 4891 861
rect 4939 839 4969 861
rect 5032 839 5062 861
rect 5118 839 5148 861
rect 5262 839 5292 861
rect 5348 839 5378 861
rect -1 823 4611 824
rect 5441 839 5471 861
rect 5519 839 5549 861
rect 5612 839 5642 861
rect 5698 839 5728 861
rect 5842 839 5872 861
rect 5928 839 5958 861
rect 6021 839 6051 861
rect 6099 839 6129 861
rect 6192 839 6222 861
rect 6278 839 6308 861
rect 6422 839 6452 861
rect 6508 839 6538 861
rect 6601 839 6631 861
rect 6679 839 6709 861
rect 6772 839 6802 861
rect 6858 839 6888 861
rect -1 794 6931 823
rect 106 766 136 794
rect 221 756 251 778
rect 299 756 329 778
rect 414 766 444 794
rect 106 716 136 738
rect 686 766 716 794
rect 801 756 831 778
rect 879 756 909 778
rect 994 766 1024 794
rect 221 695 251 728
rect 42 634 72 656
rect 128 634 143 668
rect 221 634 251 661
rect 299 695 329 728
rect 414 716 444 738
rect 686 716 716 738
rect 1266 766 1296 794
rect 1381 756 1411 778
rect 1459 756 1489 778
rect 1574 766 1604 794
rect 801 695 831 728
rect 299 634 329 661
rect 407 634 422 668
rect 478 634 508 656
rect 622 634 652 656
rect 708 634 723 668
rect 801 634 831 661
rect 879 695 909 728
rect 994 716 1024 738
rect 1266 716 1296 738
rect 1846 766 1876 794
rect 1961 756 1991 778
rect 2039 756 2069 778
rect 2154 766 2184 794
rect 1381 695 1411 728
rect 879 634 909 661
rect 987 634 1002 668
rect 1058 634 1088 656
rect 1202 634 1232 656
rect 1288 634 1303 668
rect 1381 634 1411 661
rect 1459 695 1489 728
rect 1574 716 1604 738
rect 1846 716 1876 738
rect 2426 766 2456 794
rect 2541 756 2571 778
rect 2619 756 2649 778
rect 2734 766 2764 794
rect 1961 695 1991 728
rect 1459 634 1489 661
rect 1567 634 1582 668
rect 1638 634 1668 656
rect 1782 634 1812 656
rect 1868 634 1883 668
rect 1961 634 1991 661
rect 2039 695 2069 728
rect 2154 716 2184 738
rect 2426 716 2456 738
rect 3006 766 3036 794
rect 3121 756 3151 778
rect 3199 756 3229 778
rect 3314 766 3344 794
rect 2541 695 2571 728
rect 2039 634 2069 661
rect 2147 634 2162 668
rect 2218 634 2248 656
rect 2362 634 2392 656
rect 2448 634 2463 668
rect 2541 634 2571 661
rect 2619 695 2649 728
rect 2734 716 2764 738
rect 3006 716 3036 738
rect 3586 766 3616 794
rect 3701 756 3731 778
rect 3779 756 3809 778
rect 3894 766 3924 794
rect 3121 695 3151 728
rect 2619 634 2649 661
rect 2727 634 2742 668
rect 2798 634 2828 656
rect 2942 634 2972 656
rect 3028 634 3043 668
rect 3121 634 3151 661
rect 3199 695 3229 728
rect 3314 716 3344 738
rect 3586 716 3616 738
rect 4166 766 4196 794
rect 4281 756 4311 778
rect 4359 756 4389 778
rect 4474 766 4504 794
rect 4591 793 6931 794
rect 3701 695 3731 728
rect 3199 634 3229 661
rect 3307 634 3322 668
rect 3378 634 3408 656
rect 3522 634 3552 656
rect 3608 634 3623 668
rect 3701 634 3731 661
rect 3779 695 3809 728
rect 3894 716 3924 738
rect 4166 716 4196 738
rect 4746 765 4776 793
rect 4281 695 4311 728
rect 3779 634 3809 661
rect 3887 634 3902 668
rect 3958 634 3988 656
rect 4102 634 4132 656
rect 4188 634 4203 668
rect 4281 634 4311 661
rect 4359 695 4389 728
rect 4474 716 4504 738
rect 4861 755 4891 777
rect 4939 755 4969 777
rect 5054 765 5084 793
rect 4746 715 4776 737
rect 5326 765 5356 793
rect 5441 755 5471 777
rect 5519 755 5549 777
rect 5634 765 5664 793
rect 4861 694 4891 727
rect 4359 634 4389 661
rect 4467 634 4482 668
rect 4538 634 4568 656
rect 128 620 158 634
rect 392 620 422 634
rect 708 620 738 634
rect 972 620 1002 634
rect 1288 620 1318 634
rect 1552 620 1582 634
rect 1868 620 1898 634
rect 2132 620 2162 634
rect 2448 620 2478 634
rect 2712 620 2742 634
rect 3028 620 3058 634
rect 3292 620 3322 634
rect 3608 620 3638 634
rect 3872 620 3902 634
rect 4188 620 4218 634
rect 4452 620 4482 634
rect 4682 633 4712 655
rect 4768 633 4783 667
rect 4861 633 4891 660
rect 4939 694 4969 727
rect 5054 715 5084 737
rect 5326 715 5356 737
rect 5906 765 5936 793
rect 6021 755 6051 777
rect 6099 755 6129 777
rect 6214 765 6244 793
rect 5441 694 5471 727
rect 4939 633 4969 660
rect 5047 633 5062 667
rect 5118 633 5148 655
rect 5262 633 5292 655
rect 5348 633 5363 667
rect 5441 633 5471 660
rect 5519 694 5549 727
rect 5634 715 5664 737
rect 5906 715 5936 737
rect 6486 765 6516 793
rect 6601 755 6631 777
rect 6679 755 6709 777
rect 6794 765 6824 793
rect 6021 694 6051 727
rect 5519 633 5549 660
rect 5627 633 5642 667
rect 5698 633 5728 655
rect 5842 633 5872 655
rect 5928 633 5943 667
rect 6021 633 6051 660
rect 6099 694 6129 727
rect 6214 715 6244 737
rect 6486 715 6516 737
rect 6601 694 6631 727
rect 6099 633 6129 660
rect 6207 633 6222 667
rect 6278 633 6308 655
rect 6422 633 6452 655
rect 6508 633 6523 667
rect 6601 633 6631 660
rect 6679 694 6709 727
rect 6794 715 6824 737
rect 6679 633 6709 660
rect 6787 633 6802 667
rect 6858 633 6888 655
rect 42 570 72 592
rect 128 570 158 592
rect 221 570 251 592
rect 299 570 329 592
rect 392 570 422 592
rect 478 570 508 592
rect 622 570 652 592
rect 708 570 738 592
rect 801 570 831 592
rect 879 570 909 592
rect 972 570 1002 592
rect 1058 570 1088 592
rect 1202 570 1232 592
rect 1288 570 1318 592
rect 1381 570 1411 592
rect 1459 570 1489 592
rect 1552 570 1582 592
rect 1638 570 1668 592
rect 1782 570 1812 592
rect 1868 570 1898 592
rect 1961 570 1991 592
rect 2039 570 2069 592
rect 2132 570 2162 592
rect 2218 570 2248 592
rect 2362 570 2392 592
rect 2448 570 2478 592
rect 2541 570 2571 592
rect 2619 570 2649 592
rect 2712 570 2742 592
rect 2798 570 2828 592
rect 2942 570 2972 592
rect 3028 570 3058 592
rect 3121 570 3151 592
rect 3199 570 3229 592
rect 3292 570 3322 592
rect 3378 570 3408 592
rect 3522 570 3552 592
rect 3608 570 3638 592
rect 3701 570 3731 592
rect 3779 570 3809 592
rect 3872 570 3902 592
rect 3958 570 3988 592
rect 4102 570 4132 592
rect 4188 570 4218 592
rect 4281 570 4311 592
rect 4359 570 4389 592
rect 4452 570 4482 592
rect 4538 570 4568 592
rect 4768 619 4798 633
rect 5032 619 5062 633
rect 5348 619 5378 633
rect 5612 619 5642 633
rect 5928 619 5958 633
rect 6192 619 6222 633
rect 6508 619 6538 633
rect 6772 619 6802 633
rect 4682 569 4712 591
rect 4768 569 4798 591
rect 4861 569 4891 591
rect 4939 569 4969 591
rect 5032 569 5062 591
rect 5118 569 5148 591
rect 5262 569 5292 591
rect 5348 569 5378 591
rect -1 553 4611 554
rect 5441 569 5471 591
rect 5519 569 5549 591
rect 5612 569 5642 591
rect 5698 569 5728 591
rect 5842 569 5872 591
rect 5928 569 5958 591
rect 6021 569 6051 591
rect 6099 569 6129 591
rect 6192 569 6222 591
rect 6278 569 6308 591
rect 6422 569 6452 591
rect 6508 569 6538 591
rect 6601 569 6631 591
rect 6679 569 6709 591
rect 6772 569 6802 591
rect 6858 569 6888 591
rect -1 524 6931 553
rect 106 496 136 524
rect 221 486 251 508
rect 299 486 329 508
rect 414 496 444 524
rect 106 446 136 468
rect 686 496 716 524
rect 801 486 831 508
rect 879 486 909 508
rect 994 496 1024 524
rect 221 425 251 458
rect 42 364 72 386
rect 128 364 143 398
rect 221 364 251 391
rect 299 425 329 458
rect 414 446 444 468
rect 686 446 716 468
rect 1266 496 1296 524
rect 1381 486 1411 508
rect 1459 486 1489 508
rect 1574 496 1604 524
rect 801 425 831 458
rect 299 364 329 391
rect 407 364 422 398
rect 478 364 508 386
rect 622 364 652 386
rect 708 364 723 398
rect 801 364 831 391
rect 879 425 909 458
rect 994 446 1024 468
rect 1266 446 1296 468
rect 1846 496 1876 524
rect 1961 486 1991 508
rect 2039 486 2069 508
rect 2154 496 2184 524
rect 1381 425 1411 458
rect 879 364 909 391
rect 987 364 1002 398
rect 1058 364 1088 386
rect 1202 364 1232 386
rect 1288 364 1303 398
rect 1381 364 1411 391
rect 1459 425 1489 458
rect 1574 446 1604 468
rect 1846 446 1876 468
rect 2426 496 2456 524
rect 2541 486 2571 508
rect 2619 486 2649 508
rect 2734 496 2764 524
rect 1961 425 1991 458
rect 1459 364 1489 391
rect 1567 364 1582 398
rect 1638 364 1668 386
rect 1782 364 1812 386
rect 1868 364 1883 398
rect 1961 364 1991 391
rect 2039 425 2069 458
rect 2154 446 2184 468
rect 2426 446 2456 468
rect 3006 496 3036 524
rect 3121 486 3151 508
rect 3199 486 3229 508
rect 3314 496 3344 524
rect 2541 425 2571 458
rect 2039 364 2069 391
rect 2147 364 2162 398
rect 2218 364 2248 386
rect 2362 364 2392 386
rect 2448 364 2463 398
rect 2541 364 2571 391
rect 2619 425 2649 458
rect 2734 446 2764 468
rect 3006 446 3036 468
rect 3586 496 3616 524
rect 3701 486 3731 508
rect 3779 486 3809 508
rect 3894 496 3924 524
rect 3121 425 3151 458
rect 2619 364 2649 391
rect 2727 364 2742 398
rect 2798 364 2828 386
rect 2942 364 2972 386
rect 3028 364 3043 398
rect 3121 364 3151 391
rect 3199 425 3229 458
rect 3314 446 3344 468
rect 3586 446 3616 468
rect 4166 496 4196 524
rect 4281 486 4311 508
rect 4359 486 4389 508
rect 4474 496 4504 524
rect 4591 523 6931 524
rect 3701 425 3731 458
rect 3199 364 3229 391
rect 3307 364 3322 398
rect 3378 364 3408 386
rect 3522 364 3552 386
rect 3608 364 3623 398
rect 3701 364 3731 391
rect 3779 425 3809 458
rect 3894 446 3924 468
rect 4166 446 4196 468
rect 4746 495 4776 523
rect 4281 425 4311 458
rect 3779 364 3809 391
rect 3887 364 3902 398
rect 3958 364 3988 386
rect 4102 364 4132 386
rect 4188 364 4203 398
rect 4281 364 4311 391
rect 4359 425 4389 458
rect 4474 446 4504 468
rect 4861 485 4891 507
rect 4939 485 4969 507
rect 5054 495 5084 523
rect 4746 445 4776 467
rect 5326 495 5356 523
rect 5441 485 5471 507
rect 5519 485 5549 507
rect 5634 495 5664 523
rect 4861 424 4891 457
rect 4359 364 4389 391
rect 4467 364 4482 398
rect 4538 364 4568 386
rect 128 350 158 364
rect 392 350 422 364
rect 708 350 738 364
rect 972 350 1002 364
rect 1288 350 1318 364
rect 1552 350 1582 364
rect 1868 350 1898 364
rect 2132 350 2162 364
rect 2448 350 2478 364
rect 2712 350 2742 364
rect 3028 350 3058 364
rect 3292 350 3322 364
rect 3608 350 3638 364
rect 3872 350 3902 364
rect 4188 350 4218 364
rect 4452 350 4482 364
rect 4682 363 4712 385
rect 4768 363 4783 397
rect 4861 363 4891 390
rect 4939 424 4969 457
rect 5054 445 5084 467
rect 5326 445 5356 467
rect 5906 495 5936 523
rect 6021 485 6051 507
rect 6099 485 6129 507
rect 6214 495 6244 523
rect 5441 424 5471 457
rect 4939 363 4969 390
rect 5047 363 5062 397
rect 5118 363 5148 385
rect 5262 363 5292 385
rect 5348 363 5363 397
rect 5441 363 5471 390
rect 5519 424 5549 457
rect 5634 445 5664 467
rect 5906 445 5936 467
rect 6486 495 6516 523
rect 6601 485 6631 507
rect 6679 485 6709 507
rect 6794 495 6824 523
rect 6021 424 6051 457
rect 5519 363 5549 390
rect 5627 363 5642 397
rect 5698 363 5728 385
rect 5842 363 5872 385
rect 5928 363 5943 397
rect 6021 363 6051 390
rect 6099 424 6129 457
rect 6214 445 6244 467
rect 6486 445 6516 467
rect 6601 424 6631 457
rect 6099 363 6129 390
rect 6207 363 6222 397
rect 6278 363 6308 385
rect 6422 363 6452 385
rect 6508 363 6523 397
rect 6601 363 6631 390
rect 6679 424 6709 457
rect 6794 445 6824 467
rect 6679 363 6709 390
rect 6787 363 6802 397
rect 6858 363 6888 385
rect 42 300 72 322
rect 128 300 158 322
rect 221 300 251 322
rect 299 300 329 322
rect 392 300 422 322
rect 478 300 508 322
rect 622 300 652 322
rect 708 300 738 322
rect 801 300 831 322
rect 879 300 909 322
rect 972 300 1002 322
rect 1058 300 1088 322
rect 1202 300 1232 322
rect 1288 300 1318 322
rect 1381 300 1411 322
rect 1459 300 1489 322
rect 1552 300 1582 322
rect 1638 300 1668 322
rect 1782 300 1812 322
rect 1868 300 1898 322
rect 1961 300 1991 322
rect 2039 300 2069 322
rect 2132 300 2162 322
rect 2218 300 2248 322
rect 2362 300 2392 322
rect 2448 300 2478 322
rect 2541 300 2571 322
rect 2619 300 2649 322
rect 2712 300 2742 322
rect 2798 300 2828 322
rect 2942 300 2972 322
rect 3028 300 3058 322
rect 3121 300 3151 322
rect 3199 300 3229 322
rect 3292 300 3322 322
rect 3378 300 3408 322
rect 3522 300 3552 322
rect 3608 300 3638 322
rect 3701 300 3731 322
rect 3779 300 3809 322
rect 3872 300 3902 322
rect 3958 300 3988 322
rect 4102 300 4132 322
rect 4188 300 4218 322
rect 4281 300 4311 322
rect 4359 300 4389 322
rect 4452 300 4482 322
rect 4538 300 4568 322
rect 4768 349 4798 363
rect 5032 349 5062 363
rect 5348 349 5378 363
rect 5612 349 5642 363
rect 5928 349 5958 363
rect 6192 349 6222 363
rect 6508 349 6538 363
rect 6772 349 6802 363
rect 4682 299 4712 321
rect 4768 299 4798 321
rect 4861 299 4891 321
rect 4939 299 4969 321
rect 5032 299 5062 321
rect 5118 299 5148 321
rect 5262 299 5292 321
rect 5348 299 5378 321
rect -1 283 4611 284
rect 5441 299 5471 321
rect 5519 299 5549 321
rect 5612 299 5642 321
rect 5698 299 5728 321
rect 5842 299 5872 321
rect 5928 299 5958 321
rect 6021 299 6051 321
rect 6099 299 6129 321
rect 6192 299 6222 321
rect 6278 299 6308 321
rect 6422 299 6452 321
rect 6508 299 6538 321
rect 6601 299 6631 321
rect 6679 299 6709 321
rect 6772 299 6802 321
rect 6858 299 6888 321
rect -1 254 6931 283
rect 106 226 136 254
rect 221 216 251 238
rect 299 216 329 238
rect 414 226 444 254
rect 106 176 136 198
rect 686 226 716 254
rect 801 216 831 238
rect 879 216 909 238
rect 994 226 1024 254
rect 221 155 251 188
rect 42 94 72 116
rect 128 94 143 128
rect 221 94 251 121
rect 299 155 329 188
rect 414 176 444 198
rect 686 176 716 198
rect 1266 226 1296 254
rect 1381 216 1411 238
rect 1459 216 1489 238
rect 1574 226 1604 254
rect 801 155 831 188
rect 299 94 329 121
rect 407 94 422 128
rect 478 94 508 116
rect 622 94 652 116
rect 708 94 723 128
rect 801 94 831 121
rect 879 155 909 188
rect 994 176 1024 198
rect 1266 176 1296 198
rect 1846 226 1876 254
rect 1961 216 1991 238
rect 2039 216 2069 238
rect 2154 226 2184 254
rect 1381 155 1411 188
rect 879 94 909 121
rect 987 94 1002 128
rect 1058 94 1088 116
rect 1202 94 1232 116
rect 1288 94 1303 128
rect 1381 94 1411 121
rect 1459 155 1489 188
rect 1574 176 1604 198
rect 1846 176 1876 198
rect 2426 226 2456 254
rect 2541 216 2571 238
rect 2619 216 2649 238
rect 2734 226 2764 254
rect 1961 155 1991 188
rect 1459 94 1489 121
rect 1567 94 1582 128
rect 1638 94 1668 116
rect 1782 94 1812 116
rect 1868 94 1883 128
rect 1961 94 1991 121
rect 2039 155 2069 188
rect 2154 176 2184 198
rect 2426 176 2456 198
rect 3006 226 3036 254
rect 3121 216 3151 238
rect 3199 216 3229 238
rect 3314 226 3344 254
rect 2541 155 2571 188
rect 2039 94 2069 121
rect 2147 94 2162 128
rect 2218 94 2248 116
rect 2362 94 2392 116
rect 2448 94 2463 128
rect 2541 94 2571 121
rect 2619 155 2649 188
rect 2734 176 2764 198
rect 3006 176 3036 198
rect 3586 226 3616 254
rect 3701 216 3731 238
rect 3779 216 3809 238
rect 3894 226 3924 254
rect 3121 155 3151 188
rect 2619 94 2649 121
rect 2727 94 2742 128
rect 2798 94 2828 116
rect 2942 94 2972 116
rect 3028 94 3043 128
rect 3121 94 3151 121
rect 3199 155 3229 188
rect 3314 176 3344 198
rect 3586 176 3616 198
rect 4166 226 4196 254
rect 4281 216 4311 238
rect 4359 216 4389 238
rect 4474 226 4504 254
rect 4591 253 6931 254
rect 3701 155 3731 188
rect 3199 94 3229 121
rect 3307 94 3322 128
rect 3378 94 3408 116
rect 3522 94 3552 116
rect 3608 94 3623 128
rect 3701 94 3731 121
rect 3779 155 3809 188
rect 3894 176 3924 198
rect 4166 176 4196 198
rect 4746 225 4776 253
rect 4281 155 4311 188
rect 3779 94 3809 121
rect 3887 94 3902 128
rect 3958 94 3988 116
rect 4102 94 4132 116
rect 4188 94 4203 128
rect 4281 94 4311 121
rect 4359 155 4389 188
rect 4474 176 4504 198
rect 4861 215 4891 237
rect 4939 215 4969 237
rect 5054 225 5084 253
rect 4746 175 4776 197
rect 5326 225 5356 253
rect 5441 215 5471 237
rect 5519 215 5549 237
rect 5634 225 5664 253
rect 4861 154 4891 187
rect 4359 94 4389 121
rect 4467 94 4482 128
rect 4538 94 4568 116
rect 128 80 158 94
rect 392 80 422 94
rect 708 80 738 94
rect 972 80 1002 94
rect 1288 80 1318 94
rect 1552 80 1582 94
rect 1868 80 1898 94
rect 2132 80 2162 94
rect 2448 80 2478 94
rect 2712 80 2742 94
rect 3028 80 3058 94
rect 3292 80 3322 94
rect 3608 80 3638 94
rect 3872 80 3902 94
rect 4188 80 4218 94
rect 4452 80 4482 94
rect 4682 93 4712 115
rect 4768 93 4783 127
rect 4861 93 4891 120
rect 4939 154 4969 187
rect 5054 175 5084 197
rect 5326 175 5356 197
rect 5906 225 5936 253
rect 6021 215 6051 237
rect 6099 215 6129 237
rect 6214 225 6244 253
rect 5441 154 5471 187
rect 4939 93 4969 120
rect 5047 93 5062 127
rect 5118 93 5148 115
rect 5262 93 5292 115
rect 5348 93 5363 127
rect 5441 93 5471 120
rect 5519 154 5549 187
rect 5634 175 5664 197
rect 5906 175 5936 197
rect 6486 225 6516 253
rect 6601 215 6631 237
rect 6679 215 6709 237
rect 6794 225 6824 253
rect 6021 154 6051 187
rect 5519 93 5549 120
rect 5627 93 5642 127
rect 5698 93 5728 115
rect 5842 93 5872 115
rect 5928 93 5943 127
rect 6021 93 6051 120
rect 6099 154 6129 187
rect 6214 175 6244 197
rect 6486 175 6516 197
rect 6601 154 6631 187
rect 6099 93 6129 120
rect 6207 93 6222 127
rect 6278 93 6308 115
rect 6422 93 6452 115
rect 6508 93 6523 127
rect 6601 93 6631 120
rect 6679 154 6709 187
rect 6794 175 6824 197
rect 6679 93 6709 120
rect 6787 93 6802 127
rect 6858 93 6888 115
rect 42 30 72 52
rect 128 30 158 52
rect 221 30 251 52
rect 299 30 329 52
rect 392 30 422 52
rect 478 30 508 52
rect 622 30 652 52
rect 708 30 738 52
rect 801 30 831 52
rect 879 30 909 52
rect 972 30 1002 52
rect 1058 30 1088 52
rect 1202 30 1232 52
rect 1288 30 1318 52
rect 1381 30 1411 52
rect 1459 30 1489 52
rect 1552 30 1582 52
rect 1638 30 1668 52
rect 1782 30 1812 52
rect 1868 30 1898 52
rect 1961 30 1991 52
rect 2039 30 2069 52
rect 2132 30 2162 52
rect 2218 30 2248 52
rect 2362 30 2392 52
rect 2448 30 2478 52
rect 2541 30 2571 52
rect 2619 30 2649 52
rect 2712 30 2742 52
rect 2798 30 2828 52
rect 2942 30 2972 52
rect 3028 30 3058 52
rect 3121 30 3151 52
rect 3199 30 3229 52
rect 3292 30 3322 52
rect 3378 30 3408 52
rect 3522 30 3552 52
rect 3608 30 3638 52
rect 3701 30 3731 52
rect 3779 30 3809 52
rect 3872 30 3902 52
rect 3958 30 3988 52
rect 4102 30 4132 52
rect 4188 30 4218 52
rect 4281 30 4311 52
rect 4359 30 4389 52
rect 4452 30 4482 52
rect 4538 30 4568 52
rect 4768 79 4798 93
rect 5032 79 5062 93
rect 5348 79 5378 93
rect 5612 79 5642 93
rect 5928 79 5958 93
rect 6192 79 6222 93
rect 6508 79 6538 93
rect 6772 79 6802 93
rect 4682 29 4712 51
rect 4768 29 4798 51
rect 4861 29 4891 51
rect 4939 29 4969 51
rect 5032 29 5062 51
rect 5118 29 5148 51
rect 5262 29 5292 51
rect 5348 29 5378 51
rect -1 13 4611 14
rect 5441 29 5471 51
rect 5519 29 5549 51
rect 5612 29 5642 51
rect 5698 29 5728 51
rect 5842 29 5872 51
rect 5928 29 5958 51
rect 6021 29 6051 51
rect 6099 29 6129 51
rect 6192 29 6222 51
rect 6278 29 6308 51
rect 6422 29 6452 51
rect 6508 29 6538 51
rect 6601 29 6631 51
rect 6679 29 6709 51
rect 6772 29 6802 51
rect 6858 29 6888 51
rect -1 -16 6931 13
rect 106 -44 136 -16
rect 221 -54 251 -32
rect 299 -54 329 -32
rect 414 -44 444 -16
rect 106 -94 136 -72
rect 686 -44 716 -16
rect 801 -54 831 -32
rect 879 -54 909 -32
rect 994 -44 1024 -16
rect 221 -115 251 -82
rect 42 -176 72 -154
rect 128 -176 143 -142
rect 221 -176 251 -149
rect 299 -115 329 -82
rect 414 -94 444 -72
rect 686 -94 716 -72
rect 1266 -44 1296 -16
rect 1381 -54 1411 -32
rect 1459 -54 1489 -32
rect 1574 -44 1604 -16
rect 801 -115 831 -82
rect 299 -176 329 -149
rect 407 -176 422 -142
rect 478 -176 508 -154
rect 622 -176 652 -154
rect 708 -176 723 -142
rect 801 -176 831 -149
rect 879 -115 909 -82
rect 994 -94 1024 -72
rect 1266 -94 1296 -72
rect 1846 -44 1876 -16
rect 1961 -54 1991 -32
rect 2039 -54 2069 -32
rect 2154 -44 2184 -16
rect 1381 -115 1411 -82
rect 879 -176 909 -149
rect 987 -176 1002 -142
rect 1058 -176 1088 -154
rect 1202 -176 1232 -154
rect 1288 -176 1303 -142
rect 1381 -176 1411 -149
rect 1459 -115 1489 -82
rect 1574 -94 1604 -72
rect 1846 -94 1876 -72
rect 2426 -44 2456 -16
rect 2541 -54 2571 -32
rect 2619 -54 2649 -32
rect 2734 -44 2764 -16
rect 1961 -115 1991 -82
rect 1459 -176 1489 -149
rect 1567 -176 1582 -142
rect 1638 -176 1668 -154
rect 1782 -176 1812 -154
rect 1868 -176 1883 -142
rect 1961 -176 1991 -149
rect 2039 -115 2069 -82
rect 2154 -94 2184 -72
rect 2426 -94 2456 -72
rect 3006 -44 3036 -16
rect 3121 -54 3151 -32
rect 3199 -54 3229 -32
rect 3314 -44 3344 -16
rect 2541 -115 2571 -82
rect 2039 -176 2069 -149
rect 2147 -176 2162 -142
rect 2218 -176 2248 -154
rect 2362 -176 2392 -154
rect 2448 -176 2463 -142
rect 2541 -176 2571 -149
rect 2619 -115 2649 -82
rect 2734 -94 2764 -72
rect 3006 -94 3036 -72
rect 3586 -44 3616 -16
rect 3701 -54 3731 -32
rect 3779 -54 3809 -32
rect 3894 -44 3924 -16
rect 3121 -115 3151 -82
rect 2619 -176 2649 -149
rect 2727 -176 2742 -142
rect 2798 -176 2828 -154
rect 2942 -176 2972 -154
rect 3028 -176 3043 -142
rect 3121 -176 3151 -149
rect 3199 -115 3229 -82
rect 3314 -94 3344 -72
rect 3586 -94 3616 -72
rect 4166 -44 4196 -16
rect 4281 -54 4311 -32
rect 4359 -54 4389 -32
rect 4474 -44 4504 -16
rect 4591 -17 6931 -16
rect 3701 -115 3731 -82
rect 3199 -176 3229 -149
rect 3307 -176 3322 -142
rect 3378 -176 3408 -154
rect 3522 -176 3552 -154
rect 3608 -176 3623 -142
rect 3701 -176 3731 -149
rect 3779 -115 3809 -82
rect 3894 -94 3924 -72
rect 4166 -94 4196 -72
rect 4746 -45 4776 -17
rect 4281 -115 4311 -82
rect 3779 -176 3809 -149
rect 3887 -176 3902 -142
rect 3958 -176 3988 -154
rect 4102 -176 4132 -154
rect 4188 -176 4203 -142
rect 4281 -176 4311 -149
rect 4359 -115 4389 -82
rect 4474 -94 4504 -72
rect 4861 -55 4891 -33
rect 4939 -55 4969 -33
rect 5054 -45 5084 -17
rect 4746 -95 4776 -73
rect 5326 -45 5356 -17
rect 5441 -55 5471 -33
rect 5519 -55 5549 -33
rect 5634 -45 5664 -17
rect 4861 -116 4891 -83
rect 4359 -176 4389 -149
rect 4467 -176 4482 -142
rect 4538 -176 4568 -154
rect 128 -190 158 -176
rect 392 -190 422 -176
rect 708 -190 738 -176
rect 972 -190 1002 -176
rect 1288 -190 1318 -176
rect 1552 -190 1582 -176
rect 1868 -190 1898 -176
rect 2132 -190 2162 -176
rect 2448 -190 2478 -176
rect 2712 -190 2742 -176
rect 3028 -190 3058 -176
rect 3292 -190 3322 -176
rect 3608 -190 3638 -176
rect 3872 -190 3902 -176
rect 4188 -190 4218 -176
rect 4452 -190 4482 -176
rect 4682 -177 4712 -155
rect 4768 -177 4783 -143
rect 4861 -177 4891 -150
rect 4939 -116 4969 -83
rect 5054 -95 5084 -73
rect 5326 -95 5356 -73
rect 5906 -45 5936 -17
rect 6021 -55 6051 -33
rect 6099 -55 6129 -33
rect 6214 -45 6244 -17
rect 5441 -116 5471 -83
rect 4939 -177 4969 -150
rect 5047 -177 5062 -143
rect 5118 -177 5148 -155
rect 5262 -177 5292 -155
rect 5348 -177 5363 -143
rect 5441 -177 5471 -150
rect 5519 -116 5549 -83
rect 5634 -95 5664 -73
rect 5906 -95 5936 -73
rect 6486 -45 6516 -17
rect 6601 -55 6631 -33
rect 6679 -55 6709 -33
rect 6794 -45 6824 -17
rect 6021 -116 6051 -83
rect 5519 -177 5549 -150
rect 5627 -177 5642 -143
rect 5698 -177 5728 -155
rect 5842 -177 5872 -155
rect 5928 -177 5943 -143
rect 6021 -177 6051 -150
rect 6099 -116 6129 -83
rect 6214 -95 6244 -73
rect 6486 -95 6516 -73
rect 6601 -116 6631 -83
rect 6099 -177 6129 -150
rect 6207 -177 6222 -143
rect 6278 -177 6308 -155
rect 6422 -177 6452 -155
rect 6508 -177 6523 -143
rect 6601 -177 6631 -150
rect 6679 -116 6709 -83
rect 6794 -95 6824 -73
rect 6679 -177 6709 -150
rect 6787 -177 6802 -143
rect 6858 -177 6888 -155
rect 42 -240 72 -218
rect 128 -240 158 -218
rect 221 -240 251 -218
rect 299 -240 329 -218
rect 392 -240 422 -218
rect 478 -240 508 -218
rect 622 -240 652 -218
rect 708 -240 738 -218
rect 801 -240 831 -218
rect 879 -240 909 -218
rect 972 -240 1002 -218
rect 1058 -240 1088 -218
rect 1202 -240 1232 -218
rect 1288 -240 1318 -218
rect 1381 -240 1411 -218
rect 1459 -240 1489 -218
rect 1552 -240 1582 -218
rect 1638 -240 1668 -218
rect 1782 -240 1812 -218
rect 1868 -240 1898 -218
rect 1961 -240 1991 -218
rect 2039 -240 2069 -218
rect 2132 -240 2162 -218
rect 2218 -240 2248 -218
rect 2362 -240 2392 -218
rect 2448 -240 2478 -218
rect 2541 -240 2571 -218
rect 2619 -240 2649 -218
rect 2712 -240 2742 -218
rect 2798 -240 2828 -218
rect 2942 -240 2972 -218
rect 3028 -240 3058 -218
rect 3121 -240 3151 -218
rect 3199 -240 3229 -218
rect 3292 -240 3322 -218
rect 3378 -240 3408 -218
rect 3522 -240 3552 -218
rect 3608 -240 3638 -218
rect 3701 -240 3731 -218
rect 3779 -240 3809 -218
rect 3872 -240 3902 -218
rect 3958 -240 3988 -218
rect 4102 -240 4132 -218
rect 4188 -240 4218 -218
rect 4281 -240 4311 -218
rect 4359 -240 4389 -218
rect 4452 -240 4482 -218
rect 4538 -240 4568 -218
rect 4768 -191 4798 -177
rect 5032 -191 5062 -177
rect 5348 -191 5378 -177
rect 5612 -191 5642 -177
rect 5928 -191 5958 -177
rect 6192 -191 6222 -177
rect 6508 -191 6538 -177
rect 6772 -191 6802 -177
rect 4682 -241 4712 -219
rect 4768 -241 4798 -219
rect 4861 -241 4891 -219
rect 4939 -241 4969 -219
rect 5032 -241 5062 -219
rect 5118 -241 5148 -219
rect 5262 -241 5292 -219
rect 5348 -241 5378 -219
rect -1 -257 4611 -256
rect 5441 -241 5471 -219
rect 5519 -241 5549 -219
rect 5612 -241 5642 -219
rect 5698 -241 5728 -219
rect 5842 -241 5872 -219
rect 5928 -241 5958 -219
rect 6021 -241 6051 -219
rect 6099 -241 6129 -219
rect 6192 -241 6222 -219
rect 6278 -241 6308 -219
rect 6422 -241 6452 -219
rect 6508 -241 6538 -219
rect 6601 -241 6631 -219
rect 6679 -241 6709 -219
rect 6772 -241 6802 -219
rect 6858 -241 6888 -219
rect -1 -286 6931 -257
rect 106 -314 136 -286
rect 221 -324 251 -302
rect 299 -324 329 -302
rect 414 -314 444 -286
rect 106 -364 136 -342
rect 686 -314 716 -286
rect 801 -324 831 -302
rect 879 -324 909 -302
rect 994 -314 1024 -286
rect 221 -385 251 -352
rect 42 -446 72 -424
rect 128 -446 143 -412
rect 221 -446 251 -419
rect 299 -385 329 -352
rect 414 -364 444 -342
rect 686 -364 716 -342
rect 1266 -314 1296 -286
rect 1381 -324 1411 -302
rect 1459 -324 1489 -302
rect 1574 -314 1604 -286
rect 801 -385 831 -352
rect 299 -446 329 -419
rect 407 -446 422 -412
rect 478 -446 508 -424
rect 622 -446 652 -424
rect 708 -446 723 -412
rect 801 -446 831 -419
rect 879 -385 909 -352
rect 994 -364 1024 -342
rect 1266 -364 1296 -342
rect 1846 -314 1876 -286
rect 1961 -324 1991 -302
rect 2039 -324 2069 -302
rect 2154 -314 2184 -286
rect 1381 -385 1411 -352
rect 879 -446 909 -419
rect 987 -446 1002 -412
rect 1058 -446 1088 -424
rect 1202 -446 1232 -424
rect 1288 -446 1303 -412
rect 1381 -446 1411 -419
rect 1459 -385 1489 -352
rect 1574 -364 1604 -342
rect 1846 -364 1876 -342
rect 2426 -314 2456 -286
rect 2541 -324 2571 -302
rect 2619 -324 2649 -302
rect 2734 -314 2764 -286
rect 1961 -385 1991 -352
rect 1459 -446 1489 -419
rect 1567 -446 1582 -412
rect 1638 -446 1668 -424
rect 1782 -446 1812 -424
rect 1868 -446 1883 -412
rect 1961 -446 1991 -419
rect 2039 -385 2069 -352
rect 2154 -364 2184 -342
rect 2426 -364 2456 -342
rect 3006 -314 3036 -286
rect 3121 -324 3151 -302
rect 3199 -324 3229 -302
rect 3314 -314 3344 -286
rect 2541 -385 2571 -352
rect 2039 -446 2069 -419
rect 2147 -446 2162 -412
rect 2218 -446 2248 -424
rect 2362 -446 2392 -424
rect 2448 -446 2463 -412
rect 2541 -446 2571 -419
rect 2619 -385 2649 -352
rect 2734 -364 2764 -342
rect 3006 -364 3036 -342
rect 3586 -314 3616 -286
rect 3701 -324 3731 -302
rect 3779 -324 3809 -302
rect 3894 -314 3924 -286
rect 3121 -385 3151 -352
rect 2619 -446 2649 -419
rect 2727 -446 2742 -412
rect 2798 -446 2828 -424
rect 2942 -446 2972 -424
rect 3028 -446 3043 -412
rect 3121 -446 3151 -419
rect 3199 -385 3229 -352
rect 3314 -364 3344 -342
rect 3586 -364 3616 -342
rect 4166 -314 4196 -286
rect 4281 -324 4311 -302
rect 4359 -324 4389 -302
rect 4474 -314 4504 -286
rect 4591 -287 6931 -286
rect 3701 -385 3731 -352
rect 3199 -446 3229 -419
rect 3307 -446 3322 -412
rect 3378 -446 3408 -424
rect 3522 -446 3552 -424
rect 3608 -446 3623 -412
rect 3701 -446 3731 -419
rect 3779 -385 3809 -352
rect 3894 -364 3924 -342
rect 4166 -364 4196 -342
rect 4746 -315 4776 -287
rect 4281 -385 4311 -352
rect 3779 -446 3809 -419
rect 3887 -446 3902 -412
rect 3958 -446 3988 -424
rect 4102 -446 4132 -424
rect 4188 -446 4203 -412
rect 4281 -446 4311 -419
rect 4359 -385 4389 -352
rect 4474 -364 4504 -342
rect 4861 -325 4891 -303
rect 4939 -325 4969 -303
rect 5054 -315 5084 -287
rect 4746 -365 4776 -343
rect 5326 -315 5356 -287
rect 5441 -325 5471 -303
rect 5519 -325 5549 -303
rect 5634 -315 5664 -287
rect 4861 -386 4891 -353
rect 4359 -446 4389 -419
rect 4467 -446 4482 -412
rect 4538 -446 4568 -424
rect 128 -460 158 -446
rect 392 -460 422 -446
rect 708 -460 738 -446
rect 972 -460 1002 -446
rect 1288 -460 1318 -446
rect 1552 -460 1582 -446
rect 1868 -460 1898 -446
rect 2132 -460 2162 -446
rect 2448 -460 2478 -446
rect 2712 -460 2742 -446
rect 3028 -460 3058 -446
rect 3292 -460 3322 -446
rect 3608 -460 3638 -446
rect 3872 -460 3902 -446
rect 4188 -460 4218 -446
rect 4452 -460 4482 -446
rect 4682 -447 4712 -425
rect 4768 -447 4783 -413
rect 4861 -447 4891 -420
rect 4939 -386 4969 -353
rect 5054 -365 5084 -343
rect 5326 -365 5356 -343
rect 5906 -315 5936 -287
rect 6021 -325 6051 -303
rect 6099 -325 6129 -303
rect 6214 -315 6244 -287
rect 5441 -386 5471 -353
rect 4939 -447 4969 -420
rect 5047 -447 5062 -413
rect 5118 -447 5148 -425
rect 5262 -447 5292 -425
rect 5348 -447 5363 -413
rect 5441 -447 5471 -420
rect 5519 -386 5549 -353
rect 5634 -365 5664 -343
rect 5906 -365 5936 -343
rect 6486 -315 6516 -287
rect 6601 -325 6631 -303
rect 6679 -325 6709 -303
rect 6794 -315 6824 -287
rect 6021 -386 6051 -353
rect 5519 -447 5549 -420
rect 5627 -447 5642 -413
rect 5698 -447 5728 -425
rect 5842 -447 5872 -425
rect 5928 -447 5943 -413
rect 6021 -447 6051 -420
rect 6099 -386 6129 -353
rect 6214 -365 6244 -343
rect 6486 -365 6516 -343
rect 6601 -386 6631 -353
rect 6099 -447 6129 -420
rect 6207 -447 6222 -413
rect 6278 -447 6308 -425
rect 6422 -447 6452 -425
rect 6508 -447 6523 -413
rect 6601 -447 6631 -420
rect 6679 -386 6709 -353
rect 6794 -365 6824 -343
rect 6679 -447 6709 -420
rect 6787 -447 6802 -413
rect 6858 -447 6888 -425
rect 42 -510 72 -488
rect 128 -510 158 -488
rect 221 -510 251 -488
rect 299 -510 329 -488
rect 392 -510 422 -488
rect 478 -510 508 -488
rect 622 -510 652 -488
rect 708 -510 738 -488
rect 801 -510 831 -488
rect 879 -510 909 -488
rect 972 -510 1002 -488
rect 1058 -510 1088 -488
rect 1202 -510 1232 -488
rect 1288 -510 1318 -488
rect 1381 -510 1411 -488
rect 1459 -510 1489 -488
rect 1552 -510 1582 -488
rect 1638 -510 1668 -488
rect 1782 -510 1812 -488
rect 1868 -510 1898 -488
rect 1961 -510 1991 -488
rect 2039 -510 2069 -488
rect 2132 -510 2162 -488
rect 2218 -510 2248 -488
rect 2362 -510 2392 -488
rect 2448 -510 2478 -488
rect 2541 -510 2571 -488
rect 2619 -510 2649 -488
rect 2712 -510 2742 -488
rect 2798 -510 2828 -488
rect 2942 -510 2972 -488
rect 3028 -510 3058 -488
rect 3121 -510 3151 -488
rect 3199 -510 3229 -488
rect 3292 -510 3322 -488
rect 3378 -510 3408 -488
rect 3522 -510 3552 -488
rect 3608 -510 3638 -488
rect 3701 -510 3731 -488
rect 3779 -510 3809 -488
rect 3872 -510 3902 -488
rect 3958 -510 3988 -488
rect 4102 -510 4132 -488
rect 4188 -510 4218 -488
rect 4281 -510 4311 -488
rect 4359 -510 4389 -488
rect 4452 -510 4482 -488
rect 4538 -510 4568 -488
rect 4768 -461 4798 -447
rect 5032 -461 5062 -447
rect 5348 -461 5378 -447
rect 5612 -461 5642 -447
rect 5928 -461 5958 -447
rect 6192 -461 6222 -447
rect 6508 -461 6538 -447
rect 6772 -461 6802 -447
rect 4682 -511 4712 -489
rect 4768 -511 4798 -489
rect 4861 -511 4891 -489
rect 4939 -511 4969 -489
rect 5032 -511 5062 -489
rect 5118 -511 5148 -489
rect 5262 -511 5292 -489
rect 5348 -511 5378 -489
rect -1 -527 4611 -526
rect 5441 -511 5471 -489
rect 5519 -511 5549 -489
rect 5612 -511 5642 -489
rect 5698 -511 5728 -489
rect 5842 -511 5872 -489
rect 5928 -511 5958 -489
rect 6021 -511 6051 -489
rect 6099 -511 6129 -489
rect 6192 -511 6222 -489
rect 6278 -511 6308 -489
rect 6422 -511 6452 -489
rect 6508 -511 6538 -489
rect 6601 -511 6631 -489
rect 6679 -511 6709 -489
rect 6772 -511 6802 -489
rect 6858 -511 6888 -489
rect -1 -556 6931 -527
rect 106 -584 136 -556
rect 221 -594 251 -572
rect 299 -594 329 -572
rect 414 -584 444 -556
rect 106 -634 136 -612
rect 686 -584 716 -556
rect 801 -594 831 -572
rect 879 -594 909 -572
rect 994 -584 1024 -556
rect 221 -655 251 -622
rect 42 -716 72 -694
rect 128 -716 143 -682
rect 221 -716 251 -689
rect 299 -655 329 -622
rect 414 -634 444 -612
rect 686 -634 716 -612
rect 1266 -584 1296 -556
rect 1381 -594 1411 -572
rect 1459 -594 1489 -572
rect 1574 -584 1604 -556
rect 801 -655 831 -622
rect 299 -716 329 -689
rect 407 -716 422 -682
rect 478 -716 508 -694
rect 622 -716 652 -694
rect 708 -716 723 -682
rect 801 -716 831 -689
rect 879 -655 909 -622
rect 994 -634 1024 -612
rect 1266 -634 1296 -612
rect 1846 -584 1876 -556
rect 1961 -594 1991 -572
rect 2039 -594 2069 -572
rect 2154 -584 2184 -556
rect 1381 -655 1411 -622
rect 879 -716 909 -689
rect 987 -716 1002 -682
rect 1058 -716 1088 -694
rect 1202 -716 1232 -694
rect 1288 -716 1303 -682
rect 1381 -716 1411 -689
rect 1459 -655 1489 -622
rect 1574 -634 1604 -612
rect 1846 -634 1876 -612
rect 2426 -584 2456 -556
rect 2541 -594 2571 -572
rect 2619 -594 2649 -572
rect 2734 -584 2764 -556
rect 1961 -655 1991 -622
rect 1459 -716 1489 -689
rect 1567 -716 1582 -682
rect 1638 -716 1668 -694
rect 1782 -716 1812 -694
rect 1868 -716 1883 -682
rect 1961 -716 1991 -689
rect 2039 -655 2069 -622
rect 2154 -634 2184 -612
rect 2426 -634 2456 -612
rect 3006 -584 3036 -556
rect 3121 -594 3151 -572
rect 3199 -594 3229 -572
rect 3314 -584 3344 -556
rect 2541 -655 2571 -622
rect 2039 -716 2069 -689
rect 2147 -716 2162 -682
rect 2218 -716 2248 -694
rect 2362 -716 2392 -694
rect 2448 -716 2463 -682
rect 2541 -716 2571 -689
rect 2619 -655 2649 -622
rect 2734 -634 2764 -612
rect 3006 -634 3036 -612
rect 3586 -584 3616 -556
rect 3701 -594 3731 -572
rect 3779 -594 3809 -572
rect 3894 -584 3924 -556
rect 3121 -655 3151 -622
rect 2619 -716 2649 -689
rect 2727 -716 2742 -682
rect 2798 -716 2828 -694
rect 2942 -716 2972 -694
rect 3028 -716 3043 -682
rect 3121 -716 3151 -689
rect 3199 -655 3229 -622
rect 3314 -634 3344 -612
rect 3586 -634 3616 -612
rect 4166 -584 4196 -556
rect 4281 -594 4311 -572
rect 4359 -594 4389 -572
rect 4474 -584 4504 -556
rect 4591 -557 6931 -556
rect 3701 -655 3731 -622
rect 3199 -716 3229 -689
rect 3307 -716 3322 -682
rect 3378 -716 3408 -694
rect 3522 -716 3552 -694
rect 3608 -716 3623 -682
rect 3701 -716 3731 -689
rect 3779 -655 3809 -622
rect 3894 -634 3924 -612
rect 4166 -634 4196 -612
rect 4746 -585 4776 -557
rect 4281 -655 4311 -622
rect 3779 -716 3809 -689
rect 3887 -716 3902 -682
rect 3958 -716 3988 -694
rect 4102 -716 4132 -694
rect 4188 -716 4203 -682
rect 4281 -716 4311 -689
rect 4359 -655 4389 -622
rect 4474 -634 4504 -612
rect 4861 -595 4891 -573
rect 4939 -595 4969 -573
rect 5054 -585 5084 -557
rect 4746 -635 4776 -613
rect 5326 -585 5356 -557
rect 5441 -595 5471 -573
rect 5519 -595 5549 -573
rect 5634 -585 5664 -557
rect 4861 -656 4891 -623
rect 4359 -716 4389 -689
rect 4467 -716 4482 -682
rect 4538 -716 4568 -694
rect 128 -730 158 -716
rect 392 -730 422 -716
rect 708 -730 738 -716
rect 972 -730 1002 -716
rect 1288 -730 1318 -716
rect 1552 -730 1582 -716
rect 1868 -730 1898 -716
rect 2132 -730 2162 -716
rect 2448 -730 2478 -716
rect 2712 -730 2742 -716
rect 3028 -730 3058 -716
rect 3292 -730 3322 -716
rect 3608 -730 3638 -716
rect 3872 -730 3902 -716
rect 4188 -730 4218 -716
rect 4452 -730 4482 -716
rect 4682 -717 4712 -695
rect 4768 -717 4783 -683
rect 4861 -717 4891 -690
rect 4939 -656 4969 -623
rect 5054 -635 5084 -613
rect 5326 -635 5356 -613
rect 5906 -585 5936 -557
rect 6021 -595 6051 -573
rect 6099 -595 6129 -573
rect 6214 -585 6244 -557
rect 5441 -656 5471 -623
rect 4939 -717 4969 -690
rect 5047 -717 5062 -683
rect 5118 -717 5148 -695
rect 5262 -717 5292 -695
rect 5348 -717 5363 -683
rect 5441 -717 5471 -690
rect 5519 -656 5549 -623
rect 5634 -635 5664 -613
rect 5906 -635 5936 -613
rect 6486 -585 6516 -557
rect 6601 -595 6631 -573
rect 6679 -595 6709 -573
rect 6794 -585 6824 -557
rect 6021 -656 6051 -623
rect 5519 -717 5549 -690
rect 5627 -717 5642 -683
rect 5698 -717 5728 -695
rect 5842 -717 5872 -695
rect 5928 -717 5943 -683
rect 6021 -717 6051 -690
rect 6099 -656 6129 -623
rect 6214 -635 6244 -613
rect 6486 -635 6516 -613
rect 6601 -656 6631 -623
rect 6099 -717 6129 -690
rect 6207 -717 6222 -683
rect 6278 -717 6308 -695
rect 6422 -717 6452 -695
rect 6508 -717 6523 -683
rect 6601 -717 6631 -690
rect 6679 -656 6709 -623
rect 6794 -635 6824 -613
rect 6679 -717 6709 -690
rect 6787 -717 6802 -683
rect 6858 -717 6888 -695
rect 42 -780 72 -758
rect 128 -780 158 -758
rect 221 -780 251 -758
rect 299 -780 329 -758
rect 392 -780 422 -758
rect 478 -780 508 -758
rect 622 -780 652 -758
rect 708 -780 738 -758
rect 801 -780 831 -758
rect 879 -780 909 -758
rect 972 -780 1002 -758
rect 1058 -780 1088 -758
rect 1202 -780 1232 -758
rect 1288 -780 1318 -758
rect 1381 -780 1411 -758
rect 1459 -780 1489 -758
rect 1552 -780 1582 -758
rect 1638 -780 1668 -758
rect 1782 -780 1812 -758
rect 1868 -780 1898 -758
rect 1961 -780 1991 -758
rect 2039 -780 2069 -758
rect 2132 -780 2162 -758
rect 2218 -780 2248 -758
rect 2362 -780 2392 -758
rect 2448 -780 2478 -758
rect 2541 -780 2571 -758
rect 2619 -780 2649 -758
rect 2712 -780 2742 -758
rect 2798 -780 2828 -758
rect 2942 -780 2972 -758
rect 3028 -780 3058 -758
rect 3121 -780 3151 -758
rect 3199 -780 3229 -758
rect 3292 -780 3322 -758
rect 3378 -780 3408 -758
rect 3522 -780 3552 -758
rect 3608 -780 3638 -758
rect 3701 -780 3731 -758
rect 3779 -780 3809 -758
rect 3872 -780 3902 -758
rect 3958 -780 3988 -758
rect 4102 -780 4132 -758
rect 4188 -780 4218 -758
rect 4281 -780 4311 -758
rect 4359 -780 4389 -758
rect 4452 -780 4482 -758
rect 4538 -780 4568 -758
rect 4768 -731 4798 -717
rect 5032 -731 5062 -717
rect 5348 -731 5378 -717
rect 5612 -731 5642 -717
rect 5928 -731 5958 -717
rect 6192 -731 6222 -717
rect 6508 -731 6538 -717
rect 6772 -731 6802 -717
rect 4682 -781 4712 -759
rect 4768 -781 4798 -759
rect 4861 -781 4891 -759
rect 4939 -781 4969 -759
rect 5032 -781 5062 -759
rect 5118 -781 5148 -759
rect 5262 -781 5292 -759
rect 5348 -781 5378 -759
rect -1 -797 4611 -796
rect 5441 -781 5471 -759
rect 5519 -781 5549 -759
rect 5612 -781 5642 -759
rect 5698 -781 5728 -759
rect 5842 -781 5872 -759
rect 5928 -781 5958 -759
rect 6021 -781 6051 -759
rect 6099 -781 6129 -759
rect 6192 -781 6222 -759
rect 6278 -781 6308 -759
rect 6422 -781 6452 -759
rect 6508 -781 6538 -759
rect 6601 -781 6631 -759
rect 6679 -781 6709 -759
rect 6772 -781 6802 -759
rect 6858 -781 6888 -759
rect -1 -826 6931 -797
rect 106 -854 136 -826
rect 221 -864 251 -842
rect 299 -864 329 -842
rect 414 -854 444 -826
rect 106 -904 136 -882
rect 686 -854 716 -826
rect 801 -864 831 -842
rect 879 -864 909 -842
rect 994 -854 1024 -826
rect 221 -925 251 -892
rect 42 -986 72 -964
rect 128 -986 143 -952
rect 221 -986 251 -959
rect 299 -925 329 -892
rect 414 -904 444 -882
rect 686 -904 716 -882
rect 1266 -854 1296 -826
rect 1381 -864 1411 -842
rect 1459 -864 1489 -842
rect 1574 -854 1604 -826
rect 801 -925 831 -892
rect 299 -986 329 -959
rect 407 -986 422 -952
rect 478 -986 508 -964
rect 622 -986 652 -964
rect 708 -986 723 -952
rect 801 -986 831 -959
rect 879 -925 909 -892
rect 994 -904 1024 -882
rect 1266 -904 1296 -882
rect 1846 -854 1876 -826
rect 1961 -864 1991 -842
rect 2039 -864 2069 -842
rect 2154 -854 2184 -826
rect 1381 -925 1411 -892
rect 879 -986 909 -959
rect 987 -986 1002 -952
rect 1058 -986 1088 -964
rect 1202 -986 1232 -964
rect 1288 -986 1303 -952
rect 1381 -986 1411 -959
rect 1459 -925 1489 -892
rect 1574 -904 1604 -882
rect 1846 -904 1876 -882
rect 2426 -854 2456 -826
rect 2541 -864 2571 -842
rect 2619 -864 2649 -842
rect 2734 -854 2764 -826
rect 1961 -925 1991 -892
rect 1459 -986 1489 -959
rect 1567 -986 1582 -952
rect 1638 -986 1668 -964
rect 1782 -986 1812 -964
rect 1868 -986 1883 -952
rect 1961 -986 1991 -959
rect 2039 -925 2069 -892
rect 2154 -904 2184 -882
rect 2426 -904 2456 -882
rect 3006 -854 3036 -826
rect 3121 -864 3151 -842
rect 3199 -864 3229 -842
rect 3314 -854 3344 -826
rect 2541 -925 2571 -892
rect 2039 -986 2069 -959
rect 2147 -986 2162 -952
rect 2218 -986 2248 -964
rect 2362 -986 2392 -964
rect 2448 -986 2463 -952
rect 2541 -986 2571 -959
rect 2619 -925 2649 -892
rect 2734 -904 2764 -882
rect 3006 -904 3036 -882
rect 3586 -854 3616 -826
rect 3701 -864 3731 -842
rect 3779 -864 3809 -842
rect 3894 -854 3924 -826
rect 3121 -925 3151 -892
rect 2619 -986 2649 -959
rect 2727 -986 2742 -952
rect 2798 -986 2828 -964
rect 2942 -986 2972 -964
rect 3028 -986 3043 -952
rect 3121 -986 3151 -959
rect 3199 -925 3229 -892
rect 3314 -904 3344 -882
rect 3586 -904 3616 -882
rect 4166 -854 4196 -826
rect 4281 -864 4311 -842
rect 4359 -864 4389 -842
rect 4474 -854 4504 -826
rect 4591 -827 6931 -826
rect 3701 -925 3731 -892
rect 3199 -986 3229 -959
rect 3307 -986 3322 -952
rect 3378 -986 3408 -964
rect 3522 -986 3552 -964
rect 3608 -986 3623 -952
rect 3701 -986 3731 -959
rect 3779 -925 3809 -892
rect 3894 -904 3924 -882
rect 4166 -904 4196 -882
rect 4746 -855 4776 -827
rect 4281 -925 4311 -892
rect 3779 -986 3809 -959
rect 3887 -986 3902 -952
rect 3958 -986 3988 -964
rect 4102 -986 4132 -964
rect 4188 -986 4203 -952
rect 4281 -986 4311 -959
rect 4359 -925 4389 -892
rect 4474 -904 4504 -882
rect 4861 -865 4891 -843
rect 4939 -865 4969 -843
rect 5054 -855 5084 -827
rect 4746 -905 4776 -883
rect 5326 -855 5356 -827
rect 5441 -865 5471 -843
rect 5519 -865 5549 -843
rect 5634 -855 5664 -827
rect 4861 -926 4891 -893
rect 4359 -986 4389 -959
rect 4467 -986 4482 -952
rect 4538 -986 4568 -964
rect 128 -1000 158 -986
rect 392 -1000 422 -986
rect 708 -1000 738 -986
rect 972 -1000 1002 -986
rect 1288 -1000 1318 -986
rect 1552 -1000 1582 -986
rect 1868 -1000 1898 -986
rect 2132 -1000 2162 -986
rect 2448 -1000 2478 -986
rect 2712 -1000 2742 -986
rect 3028 -1000 3058 -986
rect 3292 -1000 3322 -986
rect 3608 -1000 3638 -986
rect 3872 -1000 3902 -986
rect 4188 -1000 4218 -986
rect 4452 -1000 4482 -986
rect 4682 -987 4712 -965
rect 4768 -987 4783 -953
rect 4861 -987 4891 -960
rect 4939 -926 4969 -893
rect 5054 -905 5084 -883
rect 5326 -905 5356 -883
rect 5906 -855 5936 -827
rect 6021 -865 6051 -843
rect 6099 -865 6129 -843
rect 6214 -855 6244 -827
rect 5441 -926 5471 -893
rect 4939 -987 4969 -960
rect 5047 -987 5062 -953
rect 5118 -987 5148 -965
rect 5262 -987 5292 -965
rect 5348 -987 5363 -953
rect 5441 -987 5471 -960
rect 5519 -926 5549 -893
rect 5634 -905 5664 -883
rect 5906 -905 5936 -883
rect 6486 -855 6516 -827
rect 6601 -865 6631 -843
rect 6679 -865 6709 -843
rect 6794 -855 6824 -827
rect 6021 -926 6051 -893
rect 5519 -987 5549 -960
rect 5627 -987 5642 -953
rect 5698 -987 5728 -965
rect 5842 -987 5872 -965
rect 5928 -987 5943 -953
rect 6021 -987 6051 -960
rect 6099 -926 6129 -893
rect 6214 -905 6244 -883
rect 6486 -905 6516 -883
rect 6601 -926 6631 -893
rect 6099 -987 6129 -960
rect 6207 -987 6222 -953
rect 6278 -987 6308 -965
rect 6422 -987 6452 -965
rect 6508 -987 6523 -953
rect 6601 -987 6631 -960
rect 6679 -926 6709 -893
rect 6794 -905 6824 -883
rect 6679 -987 6709 -960
rect 6787 -987 6802 -953
rect 6858 -987 6888 -965
rect 42 -1050 72 -1028
rect 128 -1050 158 -1028
rect 221 -1050 251 -1028
rect 299 -1050 329 -1028
rect 392 -1050 422 -1028
rect 478 -1050 508 -1028
rect 622 -1050 652 -1028
rect 708 -1050 738 -1028
rect 801 -1050 831 -1028
rect 879 -1050 909 -1028
rect 972 -1050 1002 -1028
rect 1058 -1050 1088 -1028
rect 1202 -1050 1232 -1028
rect 1288 -1050 1318 -1028
rect 1381 -1050 1411 -1028
rect 1459 -1050 1489 -1028
rect 1552 -1050 1582 -1028
rect 1638 -1050 1668 -1028
rect 1782 -1050 1812 -1028
rect 1868 -1050 1898 -1028
rect 1961 -1050 1991 -1028
rect 2039 -1050 2069 -1028
rect 2132 -1050 2162 -1028
rect 2218 -1050 2248 -1028
rect 2362 -1050 2392 -1028
rect 2448 -1050 2478 -1028
rect 2541 -1050 2571 -1028
rect 2619 -1050 2649 -1028
rect 2712 -1050 2742 -1028
rect 2798 -1050 2828 -1028
rect 2942 -1050 2972 -1028
rect 3028 -1050 3058 -1028
rect 3121 -1050 3151 -1028
rect 3199 -1050 3229 -1028
rect 3292 -1050 3322 -1028
rect 3378 -1050 3408 -1028
rect 3522 -1050 3552 -1028
rect 3608 -1050 3638 -1028
rect 3701 -1050 3731 -1028
rect 3779 -1050 3809 -1028
rect 3872 -1050 3902 -1028
rect 3958 -1050 3988 -1028
rect 4102 -1050 4132 -1028
rect 4188 -1050 4218 -1028
rect 4281 -1050 4311 -1028
rect 4359 -1050 4389 -1028
rect 4452 -1050 4482 -1028
rect 4538 -1050 4568 -1028
rect 4768 -1001 4798 -987
rect 5032 -1001 5062 -987
rect 5348 -1001 5378 -987
rect 5612 -1001 5642 -987
rect 5928 -1001 5958 -987
rect 6192 -1001 6222 -987
rect 6508 -1001 6538 -987
rect 6772 -1001 6802 -987
rect 4682 -1051 4712 -1029
rect 4768 -1051 4798 -1029
rect 4861 -1051 4891 -1029
rect 4939 -1051 4969 -1029
rect 5032 -1051 5062 -1029
rect 5118 -1051 5148 -1029
rect 5262 -1051 5292 -1029
rect 5348 -1051 5378 -1029
rect -1 -1067 4611 -1066
rect 5441 -1051 5471 -1029
rect 5519 -1051 5549 -1029
rect 5612 -1051 5642 -1029
rect 5698 -1051 5728 -1029
rect 5842 -1051 5872 -1029
rect 5928 -1051 5958 -1029
rect 6021 -1051 6051 -1029
rect 6099 -1051 6129 -1029
rect 6192 -1051 6222 -1029
rect 6278 -1051 6308 -1029
rect 6422 -1051 6452 -1029
rect 6508 -1051 6538 -1029
rect 6601 -1051 6631 -1029
rect 6679 -1051 6709 -1029
rect 6772 -1051 6802 -1029
rect 6858 -1051 6888 -1029
rect -1 -1096 6931 -1067
rect 106 -1124 136 -1096
rect 221 -1134 251 -1112
rect 299 -1134 329 -1112
rect 414 -1124 444 -1096
rect 106 -1174 136 -1152
rect 686 -1124 716 -1096
rect 801 -1134 831 -1112
rect 879 -1134 909 -1112
rect 994 -1124 1024 -1096
rect 221 -1195 251 -1162
rect 42 -1256 72 -1234
rect 128 -1256 143 -1222
rect 221 -1256 251 -1229
rect 299 -1195 329 -1162
rect 414 -1174 444 -1152
rect 686 -1174 716 -1152
rect 1266 -1124 1296 -1096
rect 1381 -1134 1411 -1112
rect 1459 -1134 1489 -1112
rect 1574 -1124 1604 -1096
rect 801 -1195 831 -1162
rect 299 -1256 329 -1229
rect 407 -1256 422 -1222
rect 478 -1256 508 -1234
rect 622 -1256 652 -1234
rect 708 -1256 723 -1222
rect 801 -1256 831 -1229
rect 879 -1195 909 -1162
rect 994 -1174 1024 -1152
rect 1266 -1174 1296 -1152
rect 1846 -1124 1876 -1096
rect 1961 -1134 1991 -1112
rect 2039 -1134 2069 -1112
rect 2154 -1124 2184 -1096
rect 1381 -1195 1411 -1162
rect 879 -1256 909 -1229
rect 987 -1256 1002 -1222
rect 1058 -1256 1088 -1234
rect 1202 -1256 1232 -1234
rect 1288 -1256 1303 -1222
rect 1381 -1256 1411 -1229
rect 1459 -1195 1489 -1162
rect 1574 -1174 1604 -1152
rect 1846 -1174 1876 -1152
rect 2426 -1124 2456 -1096
rect 2541 -1134 2571 -1112
rect 2619 -1134 2649 -1112
rect 2734 -1124 2764 -1096
rect 1961 -1195 1991 -1162
rect 1459 -1256 1489 -1229
rect 1567 -1256 1582 -1222
rect 1638 -1256 1668 -1234
rect 1782 -1256 1812 -1234
rect 1868 -1256 1883 -1222
rect 1961 -1256 1991 -1229
rect 2039 -1195 2069 -1162
rect 2154 -1174 2184 -1152
rect 2426 -1174 2456 -1152
rect 3006 -1124 3036 -1096
rect 3121 -1134 3151 -1112
rect 3199 -1134 3229 -1112
rect 3314 -1124 3344 -1096
rect 2541 -1195 2571 -1162
rect 2039 -1256 2069 -1229
rect 2147 -1256 2162 -1222
rect 2218 -1256 2248 -1234
rect 2362 -1256 2392 -1234
rect 2448 -1256 2463 -1222
rect 2541 -1256 2571 -1229
rect 2619 -1195 2649 -1162
rect 2734 -1174 2764 -1152
rect 3006 -1174 3036 -1152
rect 3586 -1124 3616 -1096
rect 3701 -1134 3731 -1112
rect 3779 -1134 3809 -1112
rect 3894 -1124 3924 -1096
rect 3121 -1195 3151 -1162
rect 2619 -1256 2649 -1229
rect 2727 -1256 2742 -1222
rect 2798 -1256 2828 -1234
rect 2942 -1256 2972 -1234
rect 3028 -1256 3043 -1222
rect 3121 -1256 3151 -1229
rect 3199 -1195 3229 -1162
rect 3314 -1174 3344 -1152
rect 3586 -1174 3616 -1152
rect 4166 -1124 4196 -1096
rect 4281 -1134 4311 -1112
rect 4359 -1134 4389 -1112
rect 4474 -1124 4504 -1096
rect 4591 -1097 6931 -1096
rect 3701 -1195 3731 -1162
rect 3199 -1256 3229 -1229
rect 3307 -1256 3322 -1222
rect 3378 -1256 3408 -1234
rect 3522 -1256 3552 -1234
rect 3608 -1256 3623 -1222
rect 3701 -1256 3731 -1229
rect 3779 -1195 3809 -1162
rect 3894 -1174 3924 -1152
rect 4166 -1174 4196 -1152
rect 4746 -1125 4776 -1097
rect 4281 -1195 4311 -1162
rect 3779 -1256 3809 -1229
rect 3887 -1256 3902 -1222
rect 3958 -1256 3988 -1234
rect 4102 -1256 4132 -1234
rect 4188 -1256 4203 -1222
rect 4281 -1256 4311 -1229
rect 4359 -1195 4389 -1162
rect 4474 -1174 4504 -1152
rect 4861 -1135 4891 -1113
rect 4939 -1135 4969 -1113
rect 5054 -1125 5084 -1097
rect 4746 -1175 4776 -1153
rect 5326 -1125 5356 -1097
rect 5441 -1135 5471 -1113
rect 5519 -1135 5549 -1113
rect 5634 -1125 5664 -1097
rect 4861 -1196 4891 -1163
rect 4359 -1256 4389 -1229
rect 4467 -1256 4482 -1222
rect 4538 -1256 4568 -1234
rect 128 -1270 158 -1256
rect 392 -1270 422 -1256
rect 708 -1270 738 -1256
rect 972 -1270 1002 -1256
rect 1288 -1270 1318 -1256
rect 1552 -1270 1582 -1256
rect 1868 -1270 1898 -1256
rect 2132 -1270 2162 -1256
rect 2448 -1270 2478 -1256
rect 2712 -1270 2742 -1256
rect 3028 -1270 3058 -1256
rect 3292 -1270 3322 -1256
rect 3608 -1270 3638 -1256
rect 3872 -1270 3902 -1256
rect 4188 -1270 4218 -1256
rect 4452 -1270 4482 -1256
rect 4682 -1257 4712 -1235
rect 4768 -1257 4783 -1223
rect 4861 -1257 4891 -1230
rect 4939 -1196 4969 -1163
rect 5054 -1175 5084 -1153
rect 5326 -1175 5356 -1153
rect 5906 -1125 5936 -1097
rect 6021 -1135 6051 -1113
rect 6099 -1135 6129 -1113
rect 6214 -1125 6244 -1097
rect 5441 -1196 5471 -1163
rect 4939 -1257 4969 -1230
rect 5047 -1257 5062 -1223
rect 5118 -1257 5148 -1235
rect 5262 -1257 5292 -1235
rect 5348 -1257 5363 -1223
rect 5441 -1257 5471 -1230
rect 5519 -1196 5549 -1163
rect 5634 -1175 5664 -1153
rect 5906 -1175 5936 -1153
rect 6486 -1125 6516 -1097
rect 6601 -1135 6631 -1113
rect 6679 -1135 6709 -1113
rect 6794 -1125 6824 -1097
rect 6021 -1196 6051 -1163
rect 5519 -1257 5549 -1230
rect 5627 -1257 5642 -1223
rect 5698 -1257 5728 -1235
rect 5842 -1257 5872 -1235
rect 5928 -1257 5943 -1223
rect 6021 -1257 6051 -1230
rect 6099 -1196 6129 -1163
rect 6214 -1175 6244 -1153
rect 6486 -1175 6516 -1153
rect 6601 -1196 6631 -1163
rect 6099 -1257 6129 -1230
rect 6207 -1257 6222 -1223
rect 6278 -1257 6308 -1235
rect 6422 -1257 6452 -1235
rect 6508 -1257 6523 -1223
rect 6601 -1257 6631 -1230
rect 6679 -1196 6709 -1163
rect 6794 -1175 6824 -1153
rect 6679 -1257 6709 -1230
rect 6787 -1257 6802 -1223
rect 6858 -1257 6888 -1235
rect 42 -1320 72 -1298
rect 128 -1320 158 -1298
rect 221 -1320 251 -1298
rect 299 -1320 329 -1298
rect 392 -1320 422 -1298
rect 478 -1320 508 -1298
rect 622 -1320 652 -1298
rect 708 -1320 738 -1298
rect 801 -1320 831 -1298
rect 879 -1320 909 -1298
rect 972 -1320 1002 -1298
rect 1058 -1320 1088 -1298
rect 1202 -1320 1232 -1298
rect 1288 -1320 1318 -1298
rect 1381 -1320 1411 -1298
rect 1459 -1320 1489 -1298
rect 1552 -1320 1582 -1298
rect 1638 -1320 1668 -1298
rect 1782 -1320 1812 -1298
rect 1868 -1320 1898 -1298
rect 1961 -1320 1991 -1298
rect 2039 -1320 2069 -1298
rect 2132 -1320 2162 -1298
rect 2218 -1320 2248 -1298
rect 2362 -1320 2392 -1298
rect 2448 -1320 2478 -1298
rect 2541 -1320 2571 -1298
rect 2619 -1320 2649 -1298
rect 2712 -1320 2742 -1298
rect 2798 -1320 2828 -1298
rect 2942 -1320 2972 -1298
rect 3028 -1320 3058 -1298
rect 3121 -1320 3151 -1298
rect 3199 -1320 3229 -1298
rect 3292 -1320 3322 -1298
rect 3378 -1320 3408 -1298
rect 3522 -1320 3552 -1298
rect 3608 -1320 3638 -1298
rect 3701 -1320 3731 -1298
rect 3779 -1320 3809 -1298
rect 3872 -1320 3902 -1298
rect 3958 -1320 3988 -1298
rect 4102 -1320 4132 -1298
rect 4188 -1320 4218 -1298
rect 4281 -1320 4311 -1298
rect 4359 -1320 4389 -1298
rect 4452 -1320 4482 -1298
rect 4538 -1320 4568 -1298
rect 4768 -1271 4798 -1257
rect 5032 -1271 5062 -1257
rect 5348 -1271 5378 -1257
rect 5612 -1271 5642 -1257
rect 5928 -1271 5958 -1257
rect 6192 -1271 6222 -1257
rect 6508 -1271 6538 -1257
rect 6772 -1271 6802 -1257
rect 4682 -1321 4712 -1299
rect 4768 -1321 4798 -1299
rect 4861 -1321 4891 -1299
rect 4939 -1321 4969 -1299
rect 5032 -1321 5062 -1299
rect 5118 -1321 5148 -1299
rect 5262 -1321 5292 -1299
rect 5348 -1321 5378 -1299
rect -1 -1337 4611 -1336
rect 5441 -1321 5471 -1299
rect 5519 -1321 5549 -1299
rect 5612 -1321 5642 -1299
rect 5698 -1321 5728 -1299
rect 5842 -1321 5872 -1299
rect 5928 -1321 5958 -1299
rect 6021 -1321 6051 -1299
rect 6099 -1321 6129 -1299
rect 6192 -1321 6222 -1299
rect 6278 -1321 6308 -1299
rect 6422 -1321 6452 -1299
rect 6508 -1321 6538 -1299
rect 6601 -1321 6631 -1299
rect 6679 -1321 6709 -1299
rect 6772 -1321 6802 -1299
rect 6858 -1321 6888 -1299
rect -1 -1366 6931 -1337
rect 106 -1394 136 -1366
rect 221 -1404 251 -1382
rect 299 -1404 329 -1382
rect 414 -1394 444 -1366
rect 106 -1444 136 -1422
rect 686 -1394 716 -1366
rect 801 -1404 831 -1382
rect 879 -1404 909 -1382
rect 994 -1394 1024 -1366
rect 221 -1465 251 -1432
rect 42 -1526 72 -1504
rect 128 -1526 143 -1492
rect 221 -1526 251 -1499
rect 299 -1465 329 -1432
rect 414 -1444 444 -1422
rect 686 -1444 716 -1422
rect 1266 -1394 1296 -1366
rect 1381 -1404 1411 -1382
rect 1459 -1404 1489 -1382
rect 1574 -1394 1604 -1366
rect 801 -1465 831 -1432
rect 299 -1526 329 -1499
rect 407 -1526 422 -1492
rect 478 -1526 508 -1504
rect 622 -1526 652 -1504
rect 708 -1526 723 -1492
rect 801 -1526 831 -1499
rect 879 -1465 909 -1432
rect 994 -1444 1024 -1422
rect 1266 -1444 1296 -1422
rect 1846 -1394 1876 -1366
rect 1961 -1404 1991 -1382
rect 2039 -1404 2069 -1382
rect 2154 -1394 2184 -1366
rect 1381 -1465 1411 -1432
rect 879 -1526 909 -1499
rect 987 -1526 1002 -1492
rect 1058 -1526 1088 -1504
rect 1202 -1526 1232 -1504
rect 1288 -1526 1303 -1492
rect 1381 -1526 1411 -1499
rect 1459 -1465 1489 -1432
rect 1574 -1444 1604 -1422
rect 1846 -1444 1876 -1422
rect 2426 -1394 2456 -1366
rect 2541 -1404 2571 -1382
rect 2619 -1404 2649 -1382
rect 2734 -1394 2764 -1366
rect 1961 -1465 1991 -1432
rect 1459 -1526 1489 -1499
rect 1567 -1526 1582 -1492
rect 1638 -1526 1668 -1504
rect 1782 -1526 1812 -1504
rect 1868 -1526 1883 -1492
rect 1961 -1526 1991 -1499
rect 2039 -1465 2069 -1432
rect 2154 -1444 2184 -1422
rect 2426 -1444 2456 -1422
rect 3006 -1394 3036 -1366
rect 3121 -1404 3151 -1382
rect 3199 -1404 3229 -1382
rect 3314 -1394 3344 -1366
rect 2541 -1465 2571 -1432
rect 2039 -1526 2069 -1499
rect 2147 -1526 2162 -1492
rect 2218 -1526 2248 -1504
rect 2362 -1526 2392 -1504
rect 2448 -1526 2463 -1492
rect 2541 -1526 2571 -1499
rect 2619 -1465 2649 -1432
rect 2734 -1444 2764 -1422
rect 3006 -1444 3036 -1422
rect 3586 -1394 3616 -1366
rect 3701 -1404 3731 -1382
rect 3779 -1404 3809 -1382
rect 3894 -1394 3924 -1366
rect 3121 -1465 3151 -1432
rect 2619 -1526 2649 -1499
rect 2727 -1526 2742 -1492
rect 2798 -1526 2828 -1504
rect 2942 -1526 2972 -1504
rect 3028 -1526 3043 -1492
rect 3121 -1526 3151 -1499
rect 3199 -1465 3229 -1432
rect 3314 -1444 3344 -1422
rect 3586 -1444 3616 -1422
rect 4166 -1394 4196 -1366
rect 4281 -1404 4311 -1382
rect 4359 -1404 4389 -1382
rect 4474 -1394 4504 -1366
rect 4591 -1367 6931 -1366
rect 3701 -1465 3731 -1432
rect 3199 -1526 3229 -1499
rect 3307 -1526 3322 -1492
rect 3378 -1526 3408 -1504
rect 3522 -1526 3552 -1504
rect 3608 -1526 3623 -1492
rect 3701 -1526 3731 -1499
rect 3779 -1465 3809 -1432
rect 3894 -1444 3924 -1422
rect 4166 -1444 4196 -1422
rect 4746 -1395 4776 -1367
rect 4281 -1465 4311 -1432
rect 3779 -1526 3809 -1499
rect 3887 -1526 3902 -1492
rect 3958 -1526 3988 -1504
rect 4102 -1526 4132 -1504
rect 4188 -1526 4203 -1492
rect 4281 -1526 4311 -1499
rect 4359 -1465 4389 -1432
rect 4474 -1444 4504 -1422
rect 4861 -1405 4891 -1383
rect 4939 -1405 4969 -1383
rect 5054 -1395 5084 -1367
rect 4746 -1445 4776 -1423
rect 5326 -1395 5356 -1367
rect 5441 -1405 5471 -1383
rect 5519 -1405 5549 -1383
rect 5634 -1395 5664 -1367
rect 4861 -1466 4891 -1433
rect 4359 -1526 4389 -1499
rect 4467 -1526 4482 -1492
rect 4538 -1526 4568 -1504
rect 128 -1540 158 -1526
rect 392 -1540 422 -1526
rect 708 -1540 738 -1526
rect 972 -1540 1002 -1526
rect 1288 -1540 1318 -1526
rect 1552 -1540 1582 -1526
rect 1868 -1540 1898 -1526
rect 2132 -1540 2162 -1526
rect 2448 -1540 2478 -1526
rect 2712 -1540 2742 -1526
rect 3028 -1540 3058 -1526
rect 3292 -1540 3322 -1526
rect 3608 -1540 3638 -1526
rect 3872 -1540 3902 -1526
rect 4188 -1540 4218 -1526
rect 4452 -1540 4482 -1526
rect 4682 -1527 4712 -1505
rect 4768 -1527 4783 -1493
rect 4861 -1527 4891 -1500
rect 4939 -1466 4969 -1433
rect 5054 -1445 5084 -1423
rect 5326 -1445 5356 -1423
rect 5906 -1395 5936 -1367
rect 6021 -1405 6051 -1383
rect 6099 -1405 6129 -1383
rect 6214 -1395 6244 -1367
rect 5441 -1466 5471 -1433
rect 4939 -1527 4969 -1500
rect 5047 -1527 5062 -1493
rect 5118 -1527 5148 -1505
rect 5262 -1527 5292 -1505
rect 5348 -1527 5363 -1493
rect 5441 -1527 5471 -1500
rect 5519 -1466 5549 -1433
rect 5634 -1445 5664 -1423
rect 5906 -1445 5936 -1423
rect 6486 -1395 6516 -1367
rect 6601 -1405 6631 -1383
rect 6679 -1405 6709 -1383
rect 6794 -1395 6824 -1367
rect 6021 -1466 6051 -1433
rect 5519 -1527 5549 -1500
rect 5627 -1527 5642 -1493
rect 5698 -1527 5728 -1505
rect 5842 -1527 5872 -1505
rect 5928 -1527 5943 -1493
rect 6021 -1527 6051 -1500
rect 6099 -1466 6129 -1433
rect 6214 -1445 6244 -1423
rect 6486 -1445 6516 -1423
rect 6601 -1466 6631 -1433
rect 6099 -1527 6129 -1500
rect 6207 -1527 6222 -1493
rect 6278 -1527 6308 -1505
rect 6422 -1527 6452 -1505
rect 6508 -1527 6523 -1493
rect 6601 -1527 6631 -1500
rect 6679 -1466 6709 -1433
rect 6794 -1445 6824 -1423
rect 6679 -1527 6709 -1500
rect 6787 -1527 6802 -1493
rect 6858 -1527 6888 -1505
rect 42 -1590 72 -1568
rect 128 -1590 158 -1568
rect 221 -1590 251 -1568
rect 299 -1590 329 -1568
rect 392 -1590 422 -1568
rect 478 -1590 508 -1568
rect 622 -1590 652 -1568
rect 708 -1590 738 -1568
rect 801 -1590 831 -1568
rect 879 -1590 909 -1568
rect 972 -1590 1002 -1568
rect 1058 -1590 1088 -1568
rect 1202 -1590 1232 -1568
rect 1288 -1590 1318 -1568
rect 1381 -1590 1411 -1568
rect 1459 -1590 1489 -1568
rect 1552 -1590 1582 -1568
rect 1638 -1590 1668 -1568
rect 1782 -1590 1812 -1568
rect 1868 -1590 1898 -1568
rect 1961 -1590 1991 -1568
rect 2039 -1590 2069 -1568
rect 2132 -1590 2162 -1568
rect 2218 -1590 2248 -1568
rect 2362 -1590 2392 -1568
rect 2448 -1590 2478 -1568
rect 2541 -1590 2571 -1568
rect 2619 -1590 2649 -1568
rect 2712 -1590 2742 -1568
rect 2798 -1590 2828 -1568
rect 2942 -1590 2972 -1568
rect 3028 -1590 3058 -1568
rect 3121 -1590 3151 -1568
rect 3199 -1590 3229 -1568
rect 3292 -1590 3322 -1568
rect 3378 -1590 3408 -1568
rect 3522 -1590 3552 -1568
rect 3608 -1590 3638 -1568
rect 3701 -1590 3731 -1568
rect 3779 -1590 3809 -1568
rect 3872 -1590 3902 -1568
rect 3958 -1590 3988 -1568
rect 4102 -1590 4132 -1568
rect 4188 -1590 4218 -1568
rect 4281 -1590 4311 -1568
rect 4359 -1590 4389 -1568
rect 4452 -1590 4482 -1568
rect 4538 -1590 4568 -1568
rect 4768 -1541 4798 -1527
rect 5032 -1541 5062 -1527
rect 5348 -1541 5378 -1527
rect 5612 -1541 5642 -1527
rect 5928 -1541 5958 -1527
rect 6192 -1541 6222 -1527
rect 6508 -1541 6538 -1527
rect 6772 -1541 6802 -1527
rect 4682 -1591 4712 -1569
rect 4768 -1591 4798 -1569
rect 4861 -1591 4891 -1569
rect 4939 -1591 4969 -1569
rect 5032 -1591 5062 -1569
rect 5118 -1591 5148 -1569
rect 5262 -1591 5292 -1569
rect 5348 -1591 5378 -1569
rect -1 -1607 4611 -1606
rect 5441 -1591 5471 -1569
rect 5519 -1591 5549 -1569
rect 5612 -1591 5642 -1569
rect 5698 -1591 5728 -1569
rect 5842 -1591 5872 -1569
rect 5928 -1591 5958 -1569
rect 6021 -1591 6051 -1569
rect 6099 -1591 6129 -1569
rect 6192 -1591 6222 -1569
rect 6278 -1591 6308 -1569
rect 6422 -1591 6452 -1569
rect 6508 -1591 6538 -1569
rect 6601 -1591 6631 -1569
rect 6679 -1591 6709 -1569
rect 6772 -1591 6802 -1569
rect 6858 -1591 6888 -1569
rect -1 -1636 6931 -1607
rect 106 -1664 136 -1636
rect 221 -1674 251 -1652
rect 299 -1674 329 -1652
rect 414 -1664 444 -1636
rect 106 -1714 136 -1692
rect 686 -1664 716 -1636
rect 801 -1674 831 -1652
rect 879 -1674 909 -1652
rect 994 -1664 1024 -1636
rect 221 -1735 251 -1702
rect 42 -1796 72 -1774
rect 128 -1796 143 -1762
rect 221 -1796 251 -1769
rect 299 -1735 329 -1702
rect 414 -1714 444 -1692
rect 686 -1714 716 -1692
rect 1266 -1664 1296 -1636
rect 1381 -1674 1411 -1652
rect 1459 -1674 1489 -1652
rect 1574 -1664 1604 -1636
rect 801 -1735 831 -1702
rect 299 -1796 329 -1769
rect 407 -1796 422 -1762
rect 478 -1796 508 -1774
rect 622 -1796 652 -1774
rect 708 -1796 723 -1762
rect 801 -1796 831 -1769
rect 879 -1735 909 -1702
rect 994 -1714 1024 -1692
rect 1266 -1714 1296 -1692
rect 1846 -1664 1876 -1636
rect 1961 -1674 1991 -1652
rect 2039 -1674 2069 -1652
rect 2154 -1664 2184 -1636
rect 1381 -1735 1411 -1702
rect 879 -1796 909 -1769
rect 987 -1796 1002 -1762
rect 1058 -1796 1088 -1774
rect 1202 -1796 1232 -1774
rect 1288 -1796 1303 -1762
rect 1381 -1796 1411 -1769
rect 1459 -1735 1489 -1702
rect 1574 -1714 1604 -1692
rect 1846 -1714 1876 -1692
rect 2426 -1664 2456 -1636
rect 2541 -1674 2571 -1652
rect 2619 -1674 2649 -1652
rect 2734 -1664 2764 -1636
rect 1961 -1735 1991 -1702
rect 1459 -1796 1489 -1769
rect 1567 -1796 1582 -1762
rect 1638 -1796 1668 -1774
rect 1782 -1796 1812 -1774
rect 1868 -1796 1883 -1762
rect 1961 -1796 1991 -1769
rect 2039 -1735 2069 -1702
rect 2154 -1714 2184 -1692
rect 2426 -1714 2456 -1692
rect 3006 -1664 3036 -1636
rect 3121 -1674 3151 -1652
rect 3199 -1674 3229 -1652
rect 3314 -1664 3344 -1636
rect 2541 -1735 2571 -1702
rect 2039 -1796 2069 -1769
rect 2147 -1796 2162 -1762
rect 2218 -1796 2248 -1774
rect 2362 -1796 2392 -1774
rect 2448 -1796 2463 -1762
rect 2541 -1796 2571 -1769
rect 2619 -1735 2649 -1702
rect 2734 -1714 2764 -1692
rect 3006 -1714 3036 -1692
rect 3586 -1664 3616 -1636
rect 3701 -1674 3731 -1652
rect 3779 -1674 3809 -1652
rect 3894 -1664 3924 -1636
rect 3121 -1735 3151 -1702
rect 2619 -1796 2649 -1769
rect 2727 -1796 2742 -1762
rect 2798 -1796 2828 -1774
rect 2942 -1796 2972 -1774
rect 3028 -1796 3043 -1762
rect 3121 -1796 3151 -1769
rect 3199 -1735 3229 -1702
rect 3314 -1714 3344 -1692
rect 3586 -1714 3616 -1692
rect 4166 -1664 4196 -1636
rect 4281 -1674 4311 -1652
rect 4359 -1674 4389 -1652
rect 4474 -1664 4504 -1636
rect 4591 -1637 6931 -1636
rect 3701 -1735 3731 -1702
rect 3199 -1796 3229 -1769
rect 3307 -1796 3322 -1762
rect 3378 -1796 3408 -1774
rect 3522 -1796 3552 -1774
rect 3608 -1796 3623 -1762
rect 3701 -1796 3731 -1769
rect 3779 -1735 3809 -1702
rect 3894 -1714 3924 -1692
rect 4166 -1714 4196 -1692
rect 4746 -1665 4776 -1637
rect 4281 -1735 4311 -1702
rect 3779 -1796 3809 -1769
rect 3887 -1796 3902 -1762
rect 3958 -1796 3988 -1774
rect 4102 -1796 4132 -1774
rect 4188 -1796 4203 -1762
rect 4281 -1796 4311 -1769
rect 4359 -1735 4389 -1702
rect 4474 -1714 4504 -1692
rect 4861 -1675 4891 -1653
rect 4939 -1675 4969 -1653
rect 5054 -1665 5084 -1637
rect 4746 -1715 4776 -1693
rect 5326 -1665 5356 -1637
rect 5441 -1675 5471 -1653
rect 5519 -1675 5549 -1653
rect 5634 -1665 5664 -1637
rect 4861 -1736 4891 -1703
rect 4359 -1796 4389 -1769
rect 4467 -1796 4482 -1762
rect 4538 -1796 4568 -1774
rect 128 -1810 158 -1796
rect 392 -1810 422 -1796
rect 708 -1810 738 -1796
rect 972 -1810 1002 -1796
rect 1288 -1810 1318 -1796
rect 1552 -1810 1582 -1796
rect 1868 -1810 1898 -1796
rect 2132 -1810 2162 -1796
rect 2448 -1810 2478 -1796
rect 2712 -1810 2742 -1796
rect 3028 -1810 3058 -1796
rect 3292 -1810 3322 -1796
rect 3608 -1810 3638 -1796
rect 3872 -1810 3902 -1796
rect 4188 -1810 4218 -1796
rect 4452 -1810 4482 -1796
rect 4682 -1797 4712 -1775
rect 4768 -1797 4783 -1763
rect 4861 -1797 4891 -1770
rect 4939 -1736 4969 -1703
rect 5054 -1715 5084 -1693
rect 5326 -1715 5356 -1693
rect 5906 -1665 5936 -1637
rect 6021 -1675 6051 -1653
rect 6099 -1675 6129 -1653
rect 6214 -1665 6244 -1637
rect 5441 -1736 5471 -1703
rect 4939 -1797 4969 -1770
rect 5047 -1797 5062 -1763
rect 5118 -1797 5148 -1775
rect 5262 -1797 5292 -1775
rect 5348 -1797 5363 -1763
rect 5441 -1797 5471 -1770
rect 5519 -1736 5549 -1703
rect 5634 -1715 5664 -1693
rect 5906 -1715 5936 -1693
rect 6486 -1665 6516 -1637
rect 6601 -1675 6631 -1653
rect 6679 -1675 6709 -1653
rect 6794 -1665 6824 -1637
rect 6021 -1736 6051 -1703
rect 5519 -1797 5549 -1770
rect 5627 -1797 5642 -1763
rect 5698 -1797 5728 -1775
rect 5842 -1797 5872 -1775
rect 5928 -1797 5943 -1763
rect 6021 -1797 6051 -1770
rect 6099 -1736 6129 -1703
rect 6214 -1715 6244 -1693
rect 6486 -1715 6516 -1693
rect 6601 -1736 6631 -1703
rect 6099 -1797 6129 -1770
rect 6207 -1797 6222 -1763
rect 6278 -1797 6308 -1775
rect 6422 -1797 6452 -1775
rect 6508 -1797 6523 -1763
rect 6601 -1797 6631 -1770
rect 6679 -1736 6709 -1703
rect 6794 -1715 6824 -1693
rect 6679 -1797 6709 -1770
rect 6787 -1797 6802 -1763
rect 6858 -1797 6888 -1775
rect 42 -1860 72 -1838
rect 128 -1860 158 -1838
rect 221 -1860 251 -1838
rect 299 -1860 329 -1838
rect 392 -1860 422 -1838
rect 478 -1860 508 -1838
rect 622 -1860 652 -1838
rect 708 -1860 738 -1838
rect 801 -1860 831 -1838
rect 879 -1860 909 -1838
rect 972 -1860 1002 -1838
rect 1058 -1860 1088 -1838
rect 1202 -1860 1232 -1838
rect 1288 -1860 1318 -1838
rect 1381 -1860 1411 -1838
rect 1459 -1860 1489 -1838
rect 1552 -1860 1582 -1838
rect 1638 -1860 1668 -1838
rect 1782 -1860 1812 -1838
rect 1868 -1860 1898 -1838
rect 1961 -1860 1991 -1838
rect 2039 -1860 2069 -1838
rect 2132 -1860 2162 -1838
rect 2218 -1860 2248 -1838
rect 2362 -1860 2392 -1838
rect 2448 -1860 2478 -1838
rect 2541 -1860 2571 -1838
rect 2619 -1860 2649 -1838
rect 2712 -1860 2742 -1838
rect 2798 -1860 2828 -1838
rect 2942 -1860 2972 -1838
rect 3028 -1860 3058 -1838
rect 3121 -1860 3151 -1838
rect 3199 -1860 3229 -1838
rect 3292 -1860 3322 -1838
rect 3378 -1860 3408 -1838
rect 3522 -1860 3552 -1838
rect 3608 -1860 3638 -1838
rect 3701 -1860 3731 -1838
rect 3779 -1860 3809 -1838
rect 3872 -1860 3902 -1838
rect 3958 -1860 3988 -1838
rect 4102 -1860 4132 -1838
rect 4188 -1860 4218 -1838
rect 4281 -1860 4311 -1838
rect 4359 -1860 4389 -1838
rect 4452 -1860 4482 -1838
rect 4538 -1860 4568 -1838
rect 4768 -1811 4798 -1797
rect 5032 -1811 5062 -1797
rect 5348 -1811 5378 -1797
rect 5612 -1811 5642 -1797
rect 5928 -1811 5958 -1797
rect 6192 -1811 6222 -1797
rect 6508 -1811 6538 -1797
rect 6772 -1811 6802 -1797
rect 4682 -1861 4712 -1839
rect 4768 -1861 4798 -1839
rect 4861 -1861 4891 -1839
rect 4939 -1861 4969 -1839
rect 5032 -1861 5062 -1839
rect 5118 -1861 5148 -1839
rect 5262 -1861 5292 -1839
rect 5348 -1861 5378 -1839
rect -1 -1877 4611 -1876
rect 5441 -1861 5471 -1839
rect 5519 -1861 5549 -1839
rect 5612 -1861 5642 -1839
rect 5698 -1861 5728 -1839
rect 5842 -1861 5872 -1839
rect 5928 -1861 5958 -1839
rect 6021 -1861 6051 -1839
rect 6099 -1861 6129 -1839
rect 6192 -1861 6222 -1839
rect 6278 -1861 6308 -1839
rect 6422 -1861 6452 -1839
rect 6508 -1861 6538 -1839
rect 6601 -1861 6631 -1839
rect 6679 -1861 6709 -1839
rect 6772 -1861 6802 -1839
rect 6858 -1861 6888 -1839
rect -1 -1906 6931 -1877
rect 106 -1934 136 -1906
rect 221 -1944 251 -1922
rect 299 -1944 329 -1922
rect 414 -1934 444 -1906
rect 106 -1984 136 -1962
rect 686 -1934 716 -1906
rect 801 -1944 831 -1922
rect 879 -1944 909 -1922
rect 994 -1934 1024 -1906
rect 221 -2005 251 -1972
rect 42 -2066 72 -2044
rect 128 -2066 143 -2032
rect 221 -2066 251 -2039
rect 299 -2005 329 -1972
rect 414 -1984 444 -1962
rect 686 -1984 716 -1962
rect 1266 -1934 1296 -1906
rect 1381 -1944 1411 -1922
rect 1459 -1944 1489 -1922
rect 1574 -1934 1604 -1906
rect 801 -2005 831 -1972
rect 299 -2066 329 -2039
rect 407 -2066 422 -2032
rect 478 -2066 508 -2044
rect 622 -2066 652 -2044
rect 708 -2066 723 -2032
rect 801 -2066 831 -2039
rect 879 -2005 909 -1972
rect 994 -1984 1024 -1962
rect 1266 -1984 1296 -1962
rect 1846 -1934 1876 -1906
rect 1961 -1944 1991 -1922
rect 2039 -1944 2069 -1922
rect 2154 -1934 2184 -1906
rect 1381 -2005 1411 -1972
rect 879 -2066 909 -2039
rect 987 -2066 1002 -2032
rect 1058 -2066 1088 -2044
rect 1202 -2066 1232 -2044
rect 1288 -2066 1303 -2032
rect 1381 -2066 1411 -2039
rect 1459 -2005 1489 -1972
rect 1574 -1984 1604 -1962
rect 1846 -1984 1876 -1962
rect 2426 -1934 2456 -1906
rect 2541 -1944 2571 -1922
rect 2619 -1944 2649 -1922
rect 2734 -1934 2764 -1906
rect 1961 -2005 1991 -1972
rect 1459 -2066 1489 -2039
rect 1567 -2066 1582 -2032
rect 1638 -2066 1668 -2044
rect 1782 -2066 1812 -2044
rect 1868 -2066 1883 -2032
rect 1961 -2066 1991 -2039
rect 2039 -2005 2069 -1972
rect 2154 -1984 2184 -1962
rect 2426 -1984 2456 -1962
rect 3006 -1934 3036 -1906
rect 3121 -1944 3151 -1922
rect 3199 -1944 3229 -1922
rect 3314 -1934 3344 -1906
rect 2541 -2005 2571 -1972
rect 2039 -2066 2069 -2039
rect 2147 -2066 2162 -2032
rect 2218 -2066 2248 -2044
rect 2362 -2066 2392 -2044
rect 2448 -2066 2463 -2032
rect 2541 -2066 2571 -2039
rect 2619 -2005 2649 -1972
rect 2734 -1984 2764 -1962
rect 3006 -1984 3036 -1962
rect 3586 -1934 3616 -1906
rect 3701 -1944 3731 -1922
rect 3779 -1944 3809 -1922
rect 3894 -1934 3924 -1906
rect 3121 -2005 3151 -1972
rect 2619 -2066 2649 -2039
rect 2727 -2066 2742 -2032
rect 2798 -2066 2828 -2044
rect 2942 -2066 2972 -2044
rect 3028 -2066 3043 -2032
rect 3121 -2066 3151 -2039
rect 3199 -2005 3229 -1972
rect 3314 -1984 3344 -1962
rect 3586 -1984 3616 -1962
rect 4166 -1934 4196 -1906
rect 4281 -1944 4311 -1922
rect 4359 -1944 4389 -1922
rect 4474 -1934 4504 -1906
rect 4591 -1907 6931 -1906
rect 3701 -2005 3731 -1972
rect 3199 -2066 3229 -2039
rect 3307 -2066 3322 -2032
rect 3378 -2066 3408 -2044
rect 3522 -2066 3552 -2044
rect 3608 -2066 3623 -2032
rect 3701 -2066 3731 -2039
rect 3779 -2005 3809 -1972
rect 3894 -1984 3924 -1962
rect 4166 -1984 4196 -1962
rect 4746 -1935 4776 -1907
rect 4281 -2005 4311 -1972
rect 3779 -2066 3809 -2039
rect 3887 -2066 3902 -2032
rect 3958 -2066 3988 -2044
rect 4102 -2066 4132 -2044
rect 4188 -2066 4203 -2032
rect 4281 -2066 4311 -2039
rect 4359 -2005 4389 -1972
rect 4474 -1984 4504 -1962
rect 4861 -1945 4891 -1923
rect 4939 -1945 4969 -1923
rect 5054 -1935 5084 -1907
rect 4746 -1985 4776 -1963
rect 5326 -1935 5356 -1907
rect 5441 -1945 5471 -1923
rect 5519 -1945 5549 -1923
rect 5634 -1935 5664 -1907
rect 4861 -2006 4891 -1973
rect 4359 -2066 4389 -2039
rect 4467 -2066 4482 -2032
rect 4538 -2066 4568 -2044
rect 128 -2080 158 -2066
rect 392 -2080 422 -2066
rect 708 -2080 738 -2066
rect 972 -2080 1002 -2066
rect 1288 -2080 1318 -2066
rect 1552 -2080 1582 -2066
rect 1868 -2080 1898 -2066
rect 2132 -2080 2162 -2066
rect 2448 -2080 2478 -2066
rect 2712 -2080 2742 -2066
rect 3028 -2080 3058 -2066
rect 3292 -2080 3322 -2066
rect 3608 -2080 3638 -2066
rect 3872 -2080 3902 -2066
rect 4188 -2080 4218 -2066
rect 4452 -2080 4482 -2066
rect 4682 -2067 4712 -2045
rect 4768 -2067 4783 -2033
rect 4861 -2067 4891 -2040
rect 4939 -2006 4969 -1973
rect 5054 -1985 5084 -1963
rect 5326 -1985 5356 -1963
rect 5906 -1935 5936 -1907
rect 6021 -1945 6051 -1923
rect 6099 -1945 6129 -1923
rect 6214 -1935 6244 -1907
rect 5441 -2006 5471 -1973
rect 4939 -2067 4969 -2040
rect 5047 -2067 5062 -2033
rect 5118 -2067 5148 -2045
rect 5262 -2067 5292 -2045
rect 5348 -2067 5363 -2033
rect 5441 -2067 5471 -2040
rect 5519 -2006 5549 -1973
rect 5634 -1985 5664 -1963
rect 5906 -1985 5936 -1963
rect 6486 -1935 6516 -1907
rect 6601 -1945 6631 -1923
rect 6679 -1945 6709 -1923
rect 6794 -1935 6824 -1907
rect 6021 -2006 6051 -1973
rect 5519 -2067 5549 -2040
rect 5627 -2067 5642 -2033
rect 5698 -2067 5728 -2045
rect 5842 -2067 5872 -2045
rect 5928 -2067 5943 -2033
rect 6021 -2067 6051 -2040
rect 6099 -2006 6129 -1973
rect 6214 -1985 6244 -1963
rect 6486 -1985 6516 -1963
rect 6601 -2006 6631 -1973
rect 6099 -2067 6129 -2040
rect 6207 -2067 6222 -2033
rect 6278 -2067 6308 -2045
rect 6422 -2067 6452 -2045
rect 6508 -2067 6523 -2033
rect 6601 -2067 6631 -2040
rect 6679 -2006 6709 -1973
rect 6794 -1985 6824 -1963
rect 6679 -2067 6709 -2040
rect 6787 -2067 6802 -2033
rect 6858 -2067 6888 -2045
rect 42 -2130 72 -2108
rect 128 -2130 158 -2108
rect 221 -2130 251 -2108
rect 299 -2130 329 -2108
rect 392 -2130 422 -2108
rect 478 -2130 508 -2108
rect 622 -2130 652 -2108
rect 708 -2130 738 -2108
rect 801 -2130 831 -2108
rect 879 -2130 909 -2108
rect 972 -2130 1002 -2108
rect 1058 -2130 1088 -2108
rect 1202 -2130 1232 -2108
rect 1288 -2130 1318 -2108
rect 1381 -2130 1411 -2108
rect 1459 -2130 1489 -2108
rect 1552 -2130 1582 -2108
rect 1638 -2130 1668 -2108
rect 1782 -2130 1812 -2108
rect 1868 -2130 1898 -2108
rect 1961 -2130 1991 -2108
rect 2039 -2130 2069 -2108
rect 2132 -2130 2162 -2108
rect 2218 -2130 2248 -2108
rect 2362 -2130 2392 -2108
rect 2448 -2130 2478 -2108
rect 2541 -2130 2571 -2108
rect 2619 -2130 2649 -2108
rect 2712 -2130 2742 -2108
rect 2798 -2130 2828 -2108
rect 2942 -2130 2972 -2108
rect 3028 -2130 3058 -2108
rect 3121 -2130 3151 -2108
rect 3199 -2130 3229 -2108
rect 3292 -2130 3322 -2108
rect 3378 -2130 3408 -2108
rect 3522 -2130 3552 -2108
rect 3608 -2130 3638 -2108
rect 3701 -2130 3731 -2108
rect 3779 -2130 3809 -2108
rect 3872 -2130 3902 -2108
rect 3958 -2130 3988 -2108
rect 4102 -2130 4132 -2108
rect 4188 -2130 4218 -2108
rect 4281 -2130 4311 -2108
rect 4359 -2130 4389 -2108
rect 4452 -2130 4482 -2108
rect 4538 -2130 4568 -2108
rect 4768 -2081 4798 -2067
rect 5032 -2081 5062 -2067
rect 5348 -2081 5378 -2067
rect 5612 -2081 5642 -2067
rect 5928 -2081 5958 -2067
rect 6192 -2081 6222 -2067
rect 6508 -2081 6538 -2067
rect 6772 -2081 6802 -2067
rect 4682 -2131 4712 -2109
rect 4768 -2131 4798 -2109
rect 4861 -2131 4891 -2109
rect 4939 -2131 4969 -2109
rect 5032 -2131 5062 -2109
rect 5118 -2131 5148 -2109
rect 5262 -2131 5292 -2109
rect 5348 -2131 5378 -2109
rect 5441 -2131 5471 -2109
rect 5519 -2131 5549 -2109
rect 5612 -2131 5642 -2109
rect 5698 -2131 5728 -2109
rect 5842 -2131 5872 -2109
rect 5928 -2131 5958 -2109
rect 6021 -2131 6051 -2109
rect 6099 -2131 6129 -2109
rect 6192 -2131 6222 -2109
rect 6278 -2131 6308 -2109
rect 6422 -2131 6452 -2109
rect 6508 -2131 6538 -2109
rect 6601 -2131 6631 -2109
rect 6679 -2131 6709 -2109
rect 6772 -2131 6802 -2109
rect 6858 -2131 6888 -2109
<< polycont >>
rect 42 2006 72 2040
rect 143 1984 173 2018
rect 221 2011 251 2045
rect 299 2011 329 2045
rect 377 1984 407 2018
rect 478 2006 508 2040
rect 622 2006 652 2040
rect 723 1984 753 2018
rect 801 2011 831 2045
rect 879 2011 909 2045
rect 957 1984 987 2018
rect 1058 2006 1088 2040
rect 1202 2006 1232 2040
rect 1303 1984 1333 2018
rect 1381 2011 1411 2045
rect 1459 2011 1489 2045
rect 1537 1984 1567 2018
rect 1638 2006 1668 2040
rect 1782 2006 1812 2040
rect 1883 1984 1913 2018
rect 1961 2011 1991 2045
rect 2039 2011 2069 2045
rect 2117 1984 2147 2018
rect 2218 2006 2248 2040
rect 2362 2006 2392 2040
rect 2463 1984 2493 2018
rect 2541 2011 2571 2045
rect 2619 2011 2649 2045
rect 2697 1984 2727 2018
rect 2798 2006 2828 2040
rect 2942 2006 2972 2040
rect 3043 1984 3073 2018
rect 3121 2011 3151 2045
rect 3199 2011 3229 2045
rect 3277 1984 3307 2018
rect 3378 2006 3408 2040
rect 3522 2006 3552 2040
rect 3623 1984 3653 2018
rect 3701 2011 3731 2045
rect 3779 2011 3809 2045
rect 3857 1984 3887 2018
rect 3958 2006 3988 2040
rect 4102 2006 4132 2040
rect 4203 1984 4233 2018
rect 4281 2011 4311 2045
rect 4359 2011 4389 2045
rect 4437 1984 4467 2018
rect 4538 2006 4568 2040
rect 4682 2006 4712 2040
rect 4783 1984 4813 2018
rect 4861 2011 4891 2045
rect 4939 2011 4969 2045
rect 5017 1984 5047 2018
rect 5118 2006 5148 2040
rect 5262 2006 5292 2040
rect 5363 1984 5393 2018
rect 5441 2011 5471 2045
rect 5519 2011 5549 2045
rect 5597 1984 5627 2018
rect 5698 2006 5728 2040
rect 5842 2006 5872 2040
rect 5943 1984 5973 2018
rect 6021 2011 6051 2045
rect 6099 2011 6129 2045
rect 6177 1984 6207 2018
rect 6278 2006 6308 2040
rect 6422 2006 6452 2040
rect 6523 1984 6553 2018
rect 6601 2011 6631 2045
rect 6679 2011 6709 2045
rect 6757 1984 6787 2018
rect 6858 2006 6888 2040
rect 42 1736 72 1770
rect 143 1714 173 1748
rect 221 1741 251 1775
rect 299 1741 329 1775
rect 377 1714 407 1748
rect 478 1736 508 1770
rect 622 1736 652 1770
rect 723 1714 753 1748
rect 801 1741 831 1775
rect 879 1741 909 1775
rect 957 1714 987 1748
rect 1058 1736 1088 1770
rect 1202 1736 1232 1770
rect 1303 1714 1333 1748
rect 1381 1741 1411 1775
rect 1459 1741 1489 1775
rect 1537 1714 1567 1748
rect 1638 1736 1668 1770
rect 1782 1736 1812 1770
rect 1883 1714 1913 1748
rect 1961 1741 1991 1775
rect 2039 1741 2069 1775
rect 2117 1714 2147 1748
rect 2218 1736 2248 1770
rect 2362 1736 2392 1770
rect 2463 1714 2493 1748
rect 2541 1741 2571 1775
rect 2619 1741 2649 1775
rect 2697 1714 2727 1748
rect 2798 1736 2828 1770
rect 2942 1736 2972 1770
rect 3043 1714 3073 1748
rect 3121 1741 3151 1775
rect 3199 1741 3229 1775
rect 3277 1714 3307 1748
rect 3378 1736 3408 1770
rect 3522 1736 3552 1770
rect 3623 1714 3653 1748
rect 3701 1741 3731 1775
rect 3779 1741 3809 1775
rect 3857 1714 3887 1748
rect 3958 1736 3988 1770
rect 4102 1736 4132 1770
rect 4203 1714 4233 1748
rect 4281 1741 4311 1775
rect 4359 1741 4389 1775
rect 4437 1714 4467 1748
rect 4538 1736 4568 1770
rect 4682 1736 4712 1770
rect 4783 1714 4813 1748
rect 4861 1741 4891 1775
rect 4939 1741 4969 1775
rect 5017 1714 5047 1748
rect 5118 1736 5148 1770
rect 5262 1736 5292 1770
rect 5363 1714 5393 1748
rect 5441 1741 5471 1775
rect 5519 1741 5549 1775
rect 5597 1714 5627 1748
rect 5698 1736 5728 1770
rect 5842 1736 5872 1770
rect 5943 1714 5973 1748
rect 6021 1741 6051 1775
rect 6099 1741 6129 1775
rect 6177 1714 6207 1748
rect 6278 1736 6308 1770
rect 6422 1736 6452 1770
rect 6523 1714 6553 1748
rect 6601 1741 6631 1775
rect 6679 1741 6709 1775
rect 6757 1714 6787 1748
rect 6858 1736 6888 1770
rect 42 1466 72 1500
rect 143 1444 173 1478
rect 221 1471 251 1505
rect 299 1471 329 1505
rect 377 1444 407 1478
rect 478 1466 508 1500
rect 622 1466 652 1500
rect 723 1444 753 1478
rect 801 1471 831 1505
rect 879 1471 909 1505
rect 957 1444 987 1478
rect 1058 1466 1088 1500
rect 1202 1466 1232 1500
rect 1303 1444 1333 1478
rect 1381 1471 1411 1505
rect 1459 1471 1489 1505
rect 1537 1444 1567 1478
rect 1638 1466 1668 1500
rect 1782 1466 1812 1500
rect 1883 1444 1913 1478
rect 1961 1471 1991 1505
rect 2039 1471 2069 1505
rect 2117 1444 2147 1478
rect 2218 1466 2248 1500
rect 2362 1466 2392 1500
rect 2463 1444 2493 1478
rect 2541 1471 2571 1505
rect 2619 1471 2649 1505
rect 2697 1444 2727 1478
rect 2798 1466 2828 1500
rect 2942 1466 2972 1500
rect 3043 1444 3073 1478
rect 3121 1471 3151 1505
rect 3199 1471 3229 1505
rect 3277 1444 3307 1478
rect 3378 1466 3408 1500
rect 3522 1466 3552 1500
rect 3623 1444 3653 1478
rect 3701 1471 3731 1505
rect 3779 1471 3809 1505
rect 3857 1444 3887 1478
rect 3958 1466 3988 1500
rect 4102 1466 4132 1500
rect 4203 1444 4233 1478
rect 4281 1471 4311 1505
rect 4359 1471 4389 1505
rect 4437 1444 4467 1478
rect 4538 1466 4568 1500
rect 4682 1466 4712 1500
rect 4783 1444 4813 1478
rect 4861 1471 4891 1505
rect 4939 1471 4969 1505
rect 5017 1444 5047 1478
rect 5118 1466 5148 1500
rect 5262 1466 5292 1500
rect 5363 1444 5393 1478
rect 5441 1471 5471 1505
rect 5519 1471 5549 1505
rect 5597 1444 5627 1478
rect 5698 1466 5728 1500
rect 5842 1466 5872 1500
rect 5943 1444 5973 1478
rect 6021 1471 6051 1505
rect 6099 1471 6129 1505
rect 6177 1444 6207 1478
rect 6278 1466 6308 1500
rect 6422 1466 6452 1500
rect 6523 1444 6553 1478
rect 6601 1471 6631 1505
rect 6679 1471 6709 1505
rect 6757 1444 6787 1478
rect 6858 1466 6888 1500
rect 42 1196 72 1230
rect 143 1174 173 1208
rect 221 1201 251 1235
rect 299 1201 329 1235
rect 377 1174 407 1208
rect 478 1196 508 1230
rect 622 1196 652 1230
rect 723 1174 753 1208
rect 801 1201 831 1235
rect 879 1201 909 1235
rect 957 1174 987 1208
rect 1058 1196 1088 1230
rect 1202 1196 1232 1230
rect 1303 1174 1333 1208
rect 1381 1201 1411 1235
rect 1459 1201 1489 1235
rect 1537 1174 1567 1208
rect 1638 1196 1668 1230
rect 1782 1196 1812 1230
rect 1883 1174 1913 1208
rect 1961 1201 1991 1235
rect 2039 1201 2069 1235
rect 2117 1174 2147 1208
rect 2218 1196 2248 1230
rect 2362 1196 2392 1230
rect 2463 1174 2493 1208
rect 2541 1201 2571 1235
rect 2619 1201 2649 1235
rect 2697 1174 2727 1208
rect 2798 1196 2828 1230
rect 2942 1196 2972 1230
rect 3043 1174 3073 1208
rect 3121 1201 3151 1235
rect 3199 1201 3229 1235
rect 3277 1174 3307 1208
rect 3378 1196 3408 1230
rect 3522 1196 3552 1230
rect 3623 1174 3653 1208
rect 3701 1201 3731 1235
rect 3779 1201 3809 1235
rect 3857 1174 3887 1208
rect 3958 1196 3988 1230
rect 4102 1196 4132 1230
rect 4203 1174 4233 1208
rect 4281 1201 4311 1235
rect 4359 1201 4389 1235
rect 4437 1174 4467 1208
rect 4538 1196 4568 1230
rect 4682 1196 4712 1230
rect 4783 1174 4813 1208
rect 4861 1201 4891 1235
rect 4939 1201 4969 1235
rect 5017 1174 5047 1208
rect 5118 1196 5148 1230
rect 5262 1196 5292 1230
rect 5363 1174 5393 1208
rect 5441 1201 5471 1235
rect 5519 1201 5549 1235
rect 5597 1174 5627 1208
rect 5698 1196 5728 1230
rect 5842 1196 5872 1230
rect 5943 1174 5973 1208
rect 6021 1201 6051 1235
rect 6099 1201 6129 1235
rect 6177 1174 6207 1208
rect 6278 1196 6308 1230
rect 6422 1196 6452 1230
rect 6523 1174 6553 1208
rect 6601 1201 6631 1235
rect 6679 1201 6709 1235
rect 6757 1174 6787 1208
rect 6858 1196 6888 1230
rect 42 926 72 960
rect 143 904 173 938
rect 221 931 251 965
rect 299 931 329 965
rect 377 904 407 938
rect 478 926 508 960
rect 622 926 652 960
rect 723 904 753 938
rect 801 931 831 965
rect 879 931 909 965
rect 957 904 987 938
rect 1058 926 1088 960
rect 1202 926 1232 960
rect 1303 904 1333 938
rect 1381 931 1411 965
rect 1459 931 1489 965
rect 1537 904 1567 938
rect 1638 926 1668 960
rect 1782 926 1812 960
rect 1883 904 1913 938
rect 1961 931 1991 965
rect 2039 931 2069 965
rect 2117 904 2147 938
rect 2218 926 2248 960
rect 2362 926 2392 960
rect 2463 904 2493 938
rect 2541 931 2571 965
rect 2619 931 2649 965
rect 2697 904 2727 938
rect 2798 926 2828 960
rect 2942 926 2972 960
rect 3043 904 3073 938
rect 3121 931 3151 965
rect 3199 931 3229 965
rect 3277 904 3307 938
rect 3378 926 3408 960
rect 3522 926 3552 960
rect 3623 904 3653 938
rect 3701 931 3731 965
rect 3779 931 3809 965
rect 3857 904 3887 938
rect 3958 926 3988 960
rect 4102 926 4132 960
rect 4203 904 4233 938
rect 4281 931 4311 965
rect 4359 931 4389 965
rect 4437 904 4467 938
rect 4538 926 4568 960
rect 4682 925 4712 959
rect 4783 903 4813 937
rect 4861 930 4891 964
rect 4939 930 4969 964
rect 5017 903 5047 937
rect 5118 925 5148 959
rect 5262 925 5292 959
rect 5363 903 5393 937
rect 5441 930 5471 964
rect 5519 930 5549 964
rect 5597 903 5627 937
rect 5698 925 5728 959
rect 5842 925 5872 959
rect 5943 903 5973 937
rect 6021 930 6051 964
rect 6099 930 6129 964
rect 6177 903 6207 937
rect 6278 925 6308 959
rect 6422 925 6452 959
rect 6523 903 6553 937
rect 6601 930 6631 964
rect 6679 930 6709 964
rect 6757 903 6787 937
rect 6858 925 6888 959
rect 42 656 72 690
rect 143 634 173 668
rect 221 661 251 695
rect 299 661 329 695
rect 377 634 407 668
rect 478 656 508 690
rect 622 656 652 690
rect 723 634 753 668
rect 801 661 831 695
rect 879 661 909 695
rect 957 634 987 668
rect 1058 656 1088 690
rect 1202 656 1232 690
rect 1303 634 1333 668
rect 1381 661 1411 695
rect 1459 661 1489 695
rect 1537 634 1567 668
rect 1638 656 1668 690
rect 1782 656 1812 690
rect 1883 634 1913 668
rect 1961 661 1991 695
rect 2039 661 2069 695
rect 2117 634 2147 668
rect 2218 656 2248 690
rect 2362 656 2392 690
rect 2463 634 2493 668
rect 2541 661 2571 695
rect 2619 661 2649 695
rect 2697 634 2727 668
rect 2798 656 2828 690
rect 2942 656 2972 690
rect 3043 634 3073 668
rect 3121 661 3151 695
rect 3199 661 3229 695
rect 3277 634 3307 668
rect 3378 656 3408 690
rect 3522 656 3552 690
rect 3623 634 3653 668
rect 3701 661 3731 695
rect 3779 661 3809 695
rect 3857 634 3887 668
rect 3958 656 3988 690
rect 4102 656 4132 690
rect 4203 634 4233 668
rect 4281 661 4311 695
rect 4359 661 4389 695
rect 4437 634 4467 668
rect 4538 656 4568 690
rect 4682 655 4712 689
rect 4783 633 4813 667
rect 4861 660 4891 694
rect 4939 660 4969 694
rect 5017 633 5047 667
rect 5118 655 5148 689
rect 5262 655 5292 689
rect 5363 633 5393 667
rect 5441 660 5471 694
rect 5519 660 5549 694
rect 5597 633 5627 667
rect 5698 655 5728 689
rect 5842 655 5872 689
rect 5943 633 5973 667
rect 6021 660 6051 694
rect 6099 660 6129 694
rect 6177 633 6207 667
rect 6278 655 6308 689
rect 6422 655 6452 689
rect 6523 633 6553 667
rect 6601 660 6631 694
rect 6679 660 6709 694
rect 6757 633 6787 667
rect 6858 655 6888 689
rect 42 386 72 420
rect 143 364 173 398
rect 221 391 251 425
rect 299 391 329 425
rect 377 364 407 398
rect 478 386 508 420
rect 622 386 652 420
rect 723 364 753 398
rect 801 391 831 425
rect 879 391 909 425
rect 957 364 987 398
rect 1058 386 1088 420
rect 1202 386 1232 420
rect 1303 364 1333 398
rect 1381 391 1411 425
rect 1459 391 1489 425
rect 1537 364 1567 398
rect 1638 386 1668 420
rect 1782 386 1812 420
rect 1883 364 1913 398
rect 1961 391 1991 425
rect 2039 391 2069 425
rect 2117 364 2147 398
rect 2218 386 2248 420
rect 2362 386 2392 420
rect 2463 364 2493 398
rect 2541 391 2571 425
rect 2619 391 2649 425
rect 2697 364 2727 398
rect 2798 386 2828 420
rect 2942 386 2972 420
rect 3043 364 3073 398
rect 3121 391 3151 425
rect 3199 391 3229 425
rect 3277 364 3307 398
rect 3378 386 3408 420
rect 3522 386 3552 420
rect 3623 364 3653 398
rect 3701 391 3731 425
rect 3779 391 3809 425
rect 3857 364 3887 398
rect 3958 386 3988 420
rect 4102 386 4132 420
rect 4203 364 4233 398
rect 4281 391 4311 425
rect 4359 391 4389 425
rect 4437 364 4467 398
rect 4538 386 4568 420
rect 4682 385 4712 419
rect 4783 363 4813 397
rect 4861 390 4891 424
rect 4939 390 4969 424
rect 5017 363 5047 397
rect 5118 385 5148 419
rect 5262 385 5292 419
rect 5363 363 5393 397
rect 5441 390 5471 424
rect 5519 390 5549 424
rect 5597 363 5627 397
rect 5698 385 5728 419
rect 5842 385 5872 419
rect 5943 363 5973 397
rect 6021 390 6051 424
rect 6099 390 6129 424
rect 6177 363 6207 397
rect 6278 385 6308 419
rect 6422 385 6452 419
rect 6523 363 6553 397
rect 6601 390 6631 424
rect 6679 390 6709 424
rect 6757 363 6787 397
rect 6858 385 6888 419
rect 42 116 72 150
rect 143 94 173 128
rect 221 121 251 155
rect 299 121 329 155
rect 377 94 407 128
rect 478 116 508 150
rect 622 116 652 150
rect 723 94 753 128
rect 801 121 831 155
rect 879 121 909 155
rect 957 94 987 128
rect 1058 116 1088 150
rect 1202 116 1232 150
rect 1303 94 1333 128
rect 1381 121 1411 155
rect 1459 121 1489 155
rect 1537 94 1567 128
rect 1638 116 1668 150
rect 1782 116 1812 150
rect 1883 94 1913 128
rect 1961 121 1991 155
rect 2039 121 2069 155
rect 2117 94 2147 128
rect 2218 116 2248 150
rect 2362 116 2392 150
rect 2463 94 2493 128
rect 2541 121 2571 155
rect 2619 121 2649 155
rect 2697 94 2727 128
rect 2798 116 2828 150
rect 2942 116 2972 150
rect 3043 94 3073 128
rect 3121 121 3151 155
rect 3199 121 3229 155
rect 3277 94 3307 128
rect 3378 116 3408 150
rect 3522 116 3552 150
rect 3623 94 3653 128
rect 3701 121 3731 155
rect 3779 121 3809 155
rect 3857 94 3887 128
rect 3958 116 3988 150
rect 4102 116 4132 150
rect 4203 94 4233 128
rect 4281 121 4311 155
rect 4359 121 4389 155
rect 4437 94 4467 128
rect 4538 116 4568 150
rect 4682 115 4712 149
rect 4783 93 4813 127
rect 4861 120 4891 154
rect 4939 120 4969 154
rect 5017 93 5047 127
rect 5118 115 5148 149
rect 5262 115 5292 149
rect 5363 93 5393 127
rect 5441 120 5471 154
rect 5519 120 5549 154
rect 5597 93 5627 127
rect 5698 115 5728 149
rect 5842 115 5872 149
rect 5943 93 5973 127
rect 6021 120 6051 154
rect 6099 120 6129 154
rect 6177 93 6207 127
rect 6278 115 6308 149
rect 6422 115 6452 149
rect 6523 93 6553 127
rect 6601 120 6631 154
rect 6679 120 6709 154
rect 6757 93 6787 127
rect 6858 115 6888 149
rect 42 -154 72 -120
rect 143 -176 173 -142
rect 221 -149 251 -115
rect 299 -149 329 -115
rect 377 -176 407 -142
rect 478 -154 508 -120
rect 622 -154 652 -120
rect 723 -176 753 -142
rect 801 -149 831 -115
rect 879 -149 909 -115
rect 957 -176 987 -142
rect 1058 -154 1088 -120
rect 1202 -154 1232 -120
rect 1303 -176 1333 -142
rect 1381 -149 1411 -115
rect 1459 -149 1489 -115
rect 1537 -176 1567 -142
rect 1638 -154 1668 -120
rect 1782 -154 1812 -120
rect 1883 -176 1913 -142
rect 1961 -149 1991 -115
rect 2039 -149 2069 -115
rect 2117 -176 2147 -142
rect 2218 -154 2248 -120
rect 2362 -154 2392 -120
rect 2463 -176 2493 -142
rect 2541 -149 2571 -115
rect 2619 -149 2649 -115
rect 2697 -176 2727 -142
rect 2798 -154 2828 -120
rect 2942 -154 2972 -120
rect 3043 -176 3073 -142
rect 3121 -149 3151 -115
rect 3199 -149 3229 -115
rect 3277 -176 3307 -142
rect 3378 -154 3408 -120
rect 3522 -154 3552 -120
rect 3623 -176 3653 -142
rect 3701 -149 3731 -115
rect 3779 -149 3809 -115
rect 3857 -176 3887 -142
rect 3958 -154 3988 -120
rect 4102 -154 4132 -120
rect 4203 -176 4233 -142
rect 4281 -149 4311 -115
rect 4359 -149 4389 -115
rect 4437 -176 4467 -142
rect 4538 -154 4568 -120
rect 4682 -155 4712 -121
rect 4783 -177 4813 -143
rect 4861 -150 4891 -116
rect 4939 -150 4969 -116
rect 5017 -177 5047 -143
rect 5118 -155 5148 -121
rect 5262 -155 5292 -121
rect 5363 -177 5393 -143
rect 5441 -150 5471 -116
rect 5519 -150 5549 -116
rect 5597 -177 5627 -143
rect 5698 -155 5728 -121
rect 5842 -155 5872 -121
rect 5943 -177 5973 -143
rect 6021 -150 6051 -116
rect 6099 -150 6129 -116
rect 6177 -177 6207 -143
rect 6278 -155 6308 -121
rect 6422 -155 6452 -121
rect 6523 -177 6553 -143
rect 6601 -150 6631 -116
rect 6679 -150 6709 -116
rect 6757 -177 6787 -143
rect 6858 -155 6888 -121
rect 42 -424 72 -390
rect 143 -446 173 -412
rect 221 -419 251 -385
rect 299 -419 329 -385
rect 377 -446 407 -412
rect 478 -424 508 -390
rect 622 -424 652 -390
rect 723 -446 753 -412
rect 801 -419 831 -385
rect 879 -419 909 -385
rect 957 -446 987 -412
rect 1058 -424 1088 -390
rect 1202 -424 1232 -390
rect 1303 -446 1333 -412
rect 1381 -419 1411 -385
rect 1459 -419 1489 -385
rect 1537 -446 1567 -412
rect 1638 -424 1668 -390
rect 1782 -424 1812 -390
rect 1883 -446 1913 -412
rect 1961 -419 1991 -385
rect 2039 -419 2069 -385
rect 2117 -446 2147 -412
rect 2218 -424 2248 -390
rect 2362 -424 2392 -390
rect 2463 -446 2493 -412
rect 2541 -419 2571 -385
rect 2619 -419 2649 -385
rect 2697 -446 2727 -412
rect 2798 -424 2828 -390
rect 2942 -424 2972 -390
rect 3043 -446 3073 -412
rect 3121 -419 3151 -385
rect 3199 -419 3229 -385
rect 3277 -446 3307 -412
rect 3378 -424 3408 -390
rect 3522 -424 3552 -390
rect 3623 -446 3653 -412
rect 3701 -419 3731 -385
rect 3779 -419 3809 -385
rect 3857 -446 3887 -412
rect 3958 -424 3988 -390
rect 4102 -424 4132 -390
rect 4203 -446 4233 -412
rect 4281 -419 4311 -385
rect 4359 -419 4389 -385
rect 4437 -446 4467 -412
rect 4538 -424 4568 -390
rect 4682 -425 4712 -391
rect 4783 -447 4813 -413
rect 4861 -420 4891 -386
rect 4939 -420 4969 -386
rect 5017 -447 5047 -413
rect 5118 -425 5148 -391
rect 5262 -425 5292 -391
rect 5363 -447 5393 -413
rect 5441 -420 5471 -386
rect 5519 -420 5549 -386
rect 5597 -447 5627 -413
rect 5698 -425 5728 -391
rect 5842 -425 5872 -391
rect 5943 -447 5973 -413
rect 6021 -420 6051 -386
rect 6099 -420 6129 -386
rect 6177 -447 6207 -413
rect 6278 -425 6308 -391
rect 6422 -425 6452 -391
rect 6523 -447 6553 -413
rect 6601 -420 6631 -386
rect 6679 -420 6709 -386
rect 6757 -447 6787 -413
rect 6858 -425 6888 -391
rect 42 -694 72 -660
rect 143 -716 173 -682
rect 221 -689 251 -655
rect 299 -689 329 -655
rect 377 -716 407 -682
rect 478 -694 508 -660
rect 622 -694 652 -660
rect 723 -716 753 -682
rect 801 -689 831 -655
rect 879 -689 909 -655
rect 957 -716 987 -682
rect 1058 -694 1088 -660
rect 1202 -694 1232 -660
rect 1303 -716 1333 -682
rect 1381 -689 1411 -655
rect 1459 -689 1489 -655
rect 1537 -716 1567 -682
rect 1638 -694 1668 -660
rect 1782 -694 1812 -660
rect 1883 -716 1913 -682
rect 1961 -689 1991 -655
rect 2039 -689 2069 -655
rect 2117 -716 2147 -682
rect 2218 -694 2248 -660
rect 2362 -694 2392 -660
rect 2463 -716 2493 -682
rect 2541 -689 2571 -655
rect 2619 -689 2649 -655
rect 2697 -716 2727 -682
rect 2798 -694 2828 -660
rect 2942 -694 2972 -660
rect 3043 -716 3073 -682
rect 3121 -689 3151 -655
rect 3199 -689 3229 -655
rect 3277 -716 3307 -682
rect 3378 -694 3408 -660
rect 3522 -694 3552 -660
rect 3623 -716 3653 -682
rect 3701 -689 3731 -655
rect 3779 -689 3809 -655
rect 3857 -716 3887 -682
rect 3958 -694 3988 -660
rect 4102 -694 4132 -660
rect 4203 -716 4233 -682
rect 4281 -689 4311 -655
rect 4359 -689 4389 -655
rect 4437 -716 4467 -682
rect 4538 -694 4568 -660
rect 4682 -695 4712 -661
rect 4783 -717 4813 -683
rect 4861 -690 4891 -656
rect 4939 -690 4969 -656
rect 5017 -717 5047 -683
rect 5118 -695 5148 -661
rect 5262 -695 5292 -661
rect 5363 -717 5393 -683
rect 5441 -690 5471 -656
rect 5519 -690 5549 -656
rect 5597 -717 5627 -683
rect 5698 -695 5728 -661
rect 5842 -695 5872 -661
rect 5943 -717 5973 -683
rect 6021 -690 6051 -656
rect 6099 -690 6129 -656
rect 6177 -717 6207 -683
rect 6278 -695 6308 -661
rect 6422 -695 6452 -661
rect 6523 -717 6553 -683
rect 6601 -690 6631 -656
rect 6679 -690 6709 -656
rect 6757 -717 6787 -683
rect 6858 -695 6888 -661
rect 42 -964 72 -930
rect 143 -986 173 -952
rect 221 -959 251 -925
rect 299 -959 329 -925
rect 377 -986 407 -952
rect 478 -964 508 -930
rect 622 -964 652 -930
rect 723 -986 753 -952
rect 801 -959 831 -925
rect 879 -959 909 -925
rect 957 -986 987 -952
rect 1058 -964 1088 -930
rect 1202 -964 1232 -930
rect 1303 -986 1333 -952
rect 1381 -959 1411 -925
rect 1459 -959 1489 -925
rect 1537 -986 1567 -952
rect 1638 -964 1668 -930
rect 1782 -964 1812 -930
rect 1883 -986 1913 -952
rect 1961 -959 1991 -925
rect 2039 -959 2069 -925
rect 2117 -986 2147 -952
rect 2218 -964 2248 -930
rect 2362 -964 2392 -930
rect 2463 -986 2493 -952
rect 2541 -959 2571 -925
rect 2619 -959 2649 -925
rect 2697 -986 2727 -952
rect 2798 -964 2828 -930
rect 2942 -964 2972 -930
rect 3043 -986 3073 -952
rect 3121 -959 3151 -925
rect 3199 -959 3229 -925
rect 3277 -986 3307 -952
rect 3378 -964 3408 -930
rect 3522 -964 3552 -930
rect 3623 -986 3653 -952
rect 3701 -959 3731 -925
rect 3779 -959 3809 -925
rect 3857 -986 3887 -952
rect 3958 -964 3988 -930
rect 4102 -964 4132 -930
rect 4203 -986 4233 -952
rect 4281 -959 4311 -925
rect 4359 -959 4389 -925
rect 4437 -986 4467 -952
rect 4538 -964 4568 -930
rect 4682 -965 4712 -931
rect 4783 -987 4813 -953
rect 4861 -960 4891 -926
rect 4939 -960 4969 -926
rect 5017 -987 5047 -953
rect 5118 -965 5148 -931
rect 5262 -965 5292 -931
rect 5363 -987 5393 -953
rect 5441 -960 5471 -926
rect 5519 -960 5549 -926
rect 5597 -987 5627 -953
rect 5698 -965 5728 -931
rect 5842 -965 5872 -931
rect 5943 -987 5973 -953
rect 6021 -960 6051 -926
rect 6099 -960 6129 -926
rect 6177 -987 6207 -953
rect 6278 -965 6308 -931
rect 6422 -965 6452 -931
rect 6523 -987 6553 -953
rect 6601 -960 6631 -926
rect 6679 -960 6709 -926
rect 6757 -987 6787 -953
rect 6858 -965 6888 -931
rect 42 -1234 72 -1200
rect 143 -1256 173 -1222
rect 221 -1229 251 -1195
rect 299 -1229 329 -1195
rect 377 -1256 407 -1222
rect 478 -1234 508 -1200
rect 622 -1234 652 -1200
rect 723 -1256 753 -1222
rect 801 -1229 831 -1195
rect 879 -1229 909 -1195
rect 957 -1256 987 -1222
rect 1058 -1234 1088 -1200
rect 1202 -1234 1232 -1200
rect 1303 -1256 1333 -1222
rect 1381 -1229 1411 -1195
rect 1459 -1229 1489 -1195
rect 1537 -1256 1567 -1222
rect 1638 -1234 1668 -1200
rect 1782 -1234 1812 -1200
rect 1883 -1256 1913 -1222
rect 1961 -1229 1991 -1195
rect 2039 -1229 2069 -1195
rect 2117 -1256 2147 -1222
rect 2218 -1234 2248 -1200
rect 2362 -1234 2392 -1200
rect 2463 -1256 2493 -1222
rect 2541 -1229 2571 -1195
rect 2619 -1229 2649 -1195
rect 2697 -1256 2727 -1222
rect 2798 -1234 2828 -1200
rect 2942 -1234 2972 -1200
rect 3043 -1256 3073 -1222
rect 3121 -1229 3151 -1195
rect 3199 -1229 3229 -1195
rect 3277 -1256 3307 -1222
rect 3378 -1234 3408 -1200
rect 3522 -1234 3552 -1200
rect 3623 -1256 3653 -1222
rect 3701 -1229 3731 -1195
rect 3779 -1229 3809 -1195
rect 3857 -1256 3887 -1222
rect 3958 -1234 3988 -1200
rect 4102 -1234 4132 -1200
rect 4203 -1256 4233 -1222
rect 4281 -1229 4311 -1195
rect 4359 -1229 4389 -1195
rect 4437 -1256 4467 -1222
rect 4538 -1234 4568 -1200
rect 4682 -1235 4712 -1201
rect 4783 -1257 4813 -1223
rect 4861 -1230 4891 -1196
rect 4939 -1230 4969 -1196
rect 5017 -1257 5047 -1223
rect 5118 -1235 5148 -1201
rect 5262 -1235 5292 -1201
rect 5363 -1257 5393 -1223
rect 5441 -1230 5471 -1196
rect 5519 -1230 5549 -1196
rect 5597 -1257 5627 -1223
rect 5698 -1235 5728 -1201
rect 5842 -1235 5872 -1201
rect 5943 -1257 5973 -1223
rect 6021 -1230 6051 -1196
rect 6099 -1230 6129 -1196
rect 6177 -1257 6207 -1223
rect 6278 -1235 6308 -1201
rect 6422 -1235 6452 -1201
rect 6523 -1257 6553 -1223
rect 6601 -1230 6631 -1196
rect 6679 -1230 6709 -1196
rect 6757 -1257 6787 -1223
rect 6858 -1235 6888 -1201
rect 42 -1504 72 -1470
rect 143 -1526 173 -1492
rect 221 -1499 251 -1465
rect 299 -1499 329 -1465
rect 377 -1526 407 -1492
rect 478 -1504 508 -1470
rect 622 -1504 652 -1470
rect 723 -1526 753 -1492
rect 801 -1499 831 -1465
rect 879 -1499 909 -1465
rect 957 -1526 987 -1492
rect 1058 -1504 1088 -1470
rect 1202 -1504 1232 -1470
rect 1303 -1526 1333 -1492
rect 1381 -1499 1411 -1465
rect 1459 -1499 1489 -1465
rect 1537 -1526 1567 -1492
rect 1638 -1504 1668 -1470
rect 1782 -1504 1812 -1470
rect 1883 -1526 1913 -1492
rect 1961 -1499 1991 -1465
rect 2039 -1499 2069 -1465
rect 2117 -1526 2147 -1492
rect 2218 -1504 2248 -1470
rect 2362 -1504 2392 -1470
rect 2463 -1526 2493 -1492
rect 2541 -1499 2571 -1465
rect 2619 -1499 2649 -1465
rect 2697 -1526 2727 -1492
rect 2798 -1504 2828 -1470
rect 2942 -1504 2972 -1470
rect 3043 -1526 3073 -1492
rect 3121 -1499 3151 -1465
rect 3199 -1499 3229 -1465
rect 3277 -1526 3307 -1492
rect 3378 -1504 3408 -1470
rect 3522 -1504 3552 -1470
rect 3623 -1526 3653 -1492
rect 3701 -1499 3731 -1465
rect 3779 -1499 3809 -1465
rect 3857 -1526 3887 -1492
rect 3958 -1504 3988 -1470
rect 4102 -1504 4132 -1470
rect 4203 -1526 4233 -1492
rect 4281 -1499 4311 -1465
rect 4359 -1499 4389 -1465
rect 4437 -1526 4467 -1492
rect 4538 -1504 4568 -1470
rect 4682 -1505 4712 -1471
rect 4783 -1527 4813 -1493
rect 4861 -1500 4891 -1466
rect 4939 -1500 4969 -1466
rect 5017 -1527 5047 -1493
rect 5118 -1505 5148 -1471
rect 5262 -1505 5292 -1471
rect 5363 -1527 5393 -1493
rect 5441 -1500 5471 -1466
rect 5519 -1500 5549 -1466
rect 5597 -1527 5627 -1493
rect 5698 -1505 5728 -1471
rect 5842 -1505 5872 -1471
rect 5943 -1527 5973 -1493
rect 6021 -1500 6051 -1466
rect 6099 -1500 6129 -1466
rect 6177 -1527 6207 -1493
rect 6278 -1505 6308 -1471
rect 6422 -1505 6452 -1471
rect 6523 -1527 6553 -1493
rect 6601 -1500 6631 -1466
rect 6679 -1500 6709 -1466
rect 6757 -1527 6787 -1493
rect 6858 -1505 6888 -1471
rect 42 -1774 72 -1740
rect 143 -1796 173 -1762
rect 221 -1769 251 -1735
rect 299 -1769 329 -1735
rect 377 -1796 407 -1762
rect 478 -1774 508 -1740
rect 622 -1774 652 -1740
rect 723 -1796 753 -1762
rect 801 -1769 831 -1735
rect 879 -1769 909 -1735
rect 957 -1796 987 -1762
rect 1058 -1774 1088 -1740
rect 1202 -1774 1232 -1740
rect 1303 -1796 1333 -1762
rect 1381 -1769 1411 -1735
rect 1459 -1769 1489 -1735
rect 1537 -1796 1567 -1762
rect 1638 -1774 1668 -1740
rect 1782 -1774 1812 -1740
rect 1883 -1796 1913 -1762
rect 1961 -1769 1991 -1735
rect 2039 -1769 2069 -1735
rect 2117 -1796 2147 -1762
rect 2218 -1774 2248 -1740
rect 2362 -1774 2392 -1740
rect 2463 -1796 2493 -1762
rect 2541 -1769 2571 -1735
rect 2619 -1769 2649 -1735
rect 2697 -1796 2727 -1762
rect 2798 -1774 2828 -1740
rect 2942 -1774 2972 -1740
rect 3043 -1796 3073 -1762
rect 3121 -1769 3151 -1735
rect 3199 -1769 3229 -1735
rect 3277 -1796 3307 -1762
rect 3378 -1774 3408 -1740
rect 3522 -1774 3552 -1740
rect 3623 -1796 3653 -1762
rect 3701 -1769 3731 -1735
rect 3779 -1769 3809 -1735
rect 3857 -1796 3887 -1762
rect 3958 -1774 3988 -1740
rect 4102 -1774 4132 -1740
rect 4203 -1796 4233 -1762
rect 4281 -1769 4311 -1735
rect 4359 -1769 4389 -1735
rect 4437 -1796 4467 -1762
rect 4538 -1774 4568 -1740
rect 4682 -1775 4712 -1741
rect 4783 -1797 4813 -1763
rect 4861 -1770 4891 -1736
rect 4939 -1770 4969 -1736
rect 5017 -1797 5047 -1763
rect 5118 -1775 5148 -1741
rect 5262 -1775 5292 -1741
rect 5363 -1797 5393 -1763
rect 5441 -1770 5471 -1736
rect 5519 -1770 5549 -1736
rect 5597 -1797 5627 -1763
rect 5698 -1775 5728 -1741
rect 5842 -1775 5872 -1741
rect 5943 -1797 5973 -1763
rect 6021 -1770 6051 -1736
rect 6099 -1770 6129 -1736
rect 6177 -1797 6207 -1763
rect 6278 -1775 6308 -1741
rect 6422 -1775 6452 -1741
rect 6523 -1797 6553 -1763
rect 6601 -1770 6631 -1736
rect 6679 -1770 6709 -1736
rect 6757 -1797 6787 -1763
rect 6858 -1775 6888 -1741
rect 42 -2044 72 -2010
rect 143 -2066 173 -2032
rect 221 -2039 251 -2005
rect 299 -2039 329 -2005
rect 377 -2066 407 -2032
rect 478 -2044 508 -2010
rect 622 -2044 652 -2010
rect 723 -2066 753 -2032
rect 801 -2039 831 -2005
rect 879 -2039 909 -2005
rect 957 -2066 987 -2032
rect 1058 -2044 1088 -2010
rect 1202 -2044 1232 -2010
rect 1303 -2066 1333 -2032
rect 1381 -2039 1411 -2005
rect 1459 -2039 1489 -2005
rect 1537 -2066 1567 -2032
rect 1638 -2044 1668 -2010
rect 1782 -2044 1812 -2010
rect 1883 -2066 1913 -2032
rect 1961 -2039 1991 -2005
rect 2039 -2039 2069 -2005
rect 2117 -2066 2147 -2032
rect 2218 -2044 2248 -2010
rect 2362 -2044 2392 -2010
rect 2463 -2066 2493 -2032
rect 2541 -2039 2571 -2005
rect 2619 -2039 2649 -2005
rect 2697 -2066 2727 -2032
rect 2798 -2044 2828 -2010
rect 2942 -2044 2972 -2010
rect 3043 -2066 3073 -2032
rect 3121 -2039 3151 -2005
rect 3199 -2039 3229 -2005
rect 3277 -2066 3307 -2032
rect 3378 -2044 3408 -2010
rect 3522 -2044 3552 -2010
rect 3623 -2066 3653 -2032
rect 3701 -2039 3731 -2005
rect 3779 -2039 3809 -2005
rect 3857 -2066 3887 -2032
rect 3958 -2044 3988 -2010
rect 4102 -2044 4132 -2010
rect 4203 -2066 4233 -2032
rect 4281 -2039 4311 -2005
rect 4359 -2039 4389 -2005
rect 4437 -2066 4467 -2032
rect 4538 -2044 4568 -2010
rect 4682 -2045 4712 -2011
rect 4783 -2067 4813 -2033
rect 4861 -2040 4891 -2006
rect 4939 -2040 4969 -2006
rect 5017 -2067 5047 -2033
rect 5118 -2045 5148 -2011
rect 5262 -2045 5292 -2011
rect 5363 -2067 5393 -2033
rect 5441 -2040 5471 -2006
rect 5519 -2040 5549 -2006
rect 5597 -2067 5627 -2033
rect 5698 -2045 5728 -2011
rect 5842 -2045 5872 -2011
rect 5943 -2067 5973 -2033
rect 6021 -2040 6051 -2006
rect 6099 -2040 6129 -2006
rect 6177 -2067 6207 -2033
rect 6278 -2045 6308 -2011
rect 6422 -2045 6452 -2011
rect 6523 -2067 6553 -2033
rect 6601 -2040 6631 -2006
rect 6679 -2040 6709 -2006
rect 6757 -2067 6787 -2033
rect 6858 -2045 6888 -2011
<< corelocali >>
rect -1 1984 14 2174
tri 79 2138 101 2160 se
rect 101 2153 116 2174
tri 101 2138 116 2153 nw
rect 435 2153 450 2174
tri 73 2132 79 2138 se
rect 79 2132 88 2138
rect 73 2116 88 2132
tri 88 2125 101 2138 nw
rect 242 2130 259 2144
rect 291 2130 308 2144
tri 435 2138 450 2153 ne
tri 450 2138 472 2160 sw
rect 73 2080 88 2088
rect 154 2116 214 2130
rect 169 2106 214 2116
rect 169 2088 197 2106
tri 73 2065 88 2080 ne
tri 88 2065 110 2087 sw
rect 154 2078 197 2088
rect 212 2102 214 2106
rect 336 2116 396 2130
tri 450 2125 463 2138 ne
rect 463 2132 472 2138
tri 472 2132 478 2138 sw
rect 336 2106 381 2116
rect 212 2078 286 2102
rect 154 2074 286 2078
tri 286 2074 314 2102 sw
rect 336 2092 338 2106
tri 336 2090 338 2092 ne
rect 350 2088 381 2106
rect 350 2078 396 2088
rect 463 2117 478 2132
tri 88 2053 100 2065 ne
rect 100 2060 110 2065
tri 110 2060 115 2065 sw
rect -1 1714 14 1942
rect 100 1904 115 2060
rect 154 2018 182 2074
tri 274 2056 292 2074 ne
rect 292 2054 314 2074
tri 314 2054 334 2074 sw
tri 350 2060 368 2078 ne
rect 173 1984 182 2018
rect 216 2045 258 2046
rect 216 2011 221 2045
rect 251 2011 258 2045
rect 216 2002 258 2011
rect 292 2045 334 2054
rect 292 2011 299 2045
rect 329 2011 334 2045
rect 292 2006 334 2011
rect 368 2018 396 2078
tri 441 2065 463 2087 se
rect 463 2080 478 2088
tri 463 2065 478 2080 nw
tri 435 2059 441 2065 se
rect 441 2059 450 2065
rect 154 1974 182 1984
tri 182 1974 206 1998 sw
rect 154 1942 196 1974
tri 213 1966 214 1967 sw
rect 213 1942 214 1966
tri 216 1965 253 2002 ne
rect 253 1974 258 2002
tri 258 1974 284 2000 sw
rect 368 1984 377 2018
rect 368 1974 396 1984
rect 253 1965 337 1974
tri 253 1946 272 1965 ne
rect 272 1946 337 1965
rect 154 1920 214 1942
rect 336 1942 337 1946
rect 354 1942 396 1974
rect 336 1920 396 1942
rect 242 1904 259 1918
rect 291 1904 308 1918
tri 79 1868 101 1890 se
rect 101 1883 116 1904
tri 101 1868 116 1883 nw
rect 435 1883 450 2059
tri 450 2052 463 2065 nw
rect 536 1984 551 2174
tri 73 1862 79 1868 se
rect 79 1862 88 1868
rect 73 1846 88 1862
tri 88 1855 101 1868 nw
rect 242 1860 259 1874
rect 291 1860 308 1874
tri 435 1868 450 1883 ne
tri 450 1868 472 1890 sw
rect 73 1810 88 1818
rect 154 1846 214 1860
rect 169 1836 214 1846
rect 169 1818 197 1836
tri 73 1795 88 1810 ne
tri 88 1795 110 1817 sw
rect 154 1808 197 1818
rect 212 1832 214 1836
rect 336 1846 396 1860
tri 450 1855 463 1868 ne
rect 463 1862 472 1868
tri 472 1862 478 1868 sw
rect 336 1836 381 1846
rect 212 1808 286 1832
rect 154 1804 286 1808
tri 286 1804 314 1832 sw
rect 336 1822 338 1836
tri 336 1820 338 1822 ne
rect 350 1818 381 1836
rect 350 1808 396 1818
rect 463 1847 478 1862
tri 88 1783 100 1795 ne
rect 100 1790 110 1795
tri 110 1790 115 1795 sw
rect -1 1444 14 1672
rect 100 1634 115 1790
rect 154 1748 182 1804
tri 274 1786 292 1804 ne
rect 292 1784 314 1804
tri 314 1784 334 1804 sw
tri 350 1790 368 1808 ne
rect 173 1714 182 1748
rect 216 1775 258 1776
rect 216 1741 221 1775
rect 251 1741 258 1775
rect 216 1732 258 1741
rect 292 1775 334 1784
rect 292 1741 299 1775
rect 329 1741 334 1775
rect 292 1736 334 1741
rect 368 1748 396 1808
tri 441 1795 463 1817 se
rect 463 1810 478 1818
tri 463 1795 478 1810 nw
tri 435 1789 441 1795 se
rect 441 1789 450 1795
rect 154 1704 182 1714
tri 182 1704 206 1728 sw
rect 154 1672 196 1704
tri 213 1696 214 1697 sw
rect 213 1672 214 1696
tri 216 1695 253 1732 ne
rect 253 1704 258 1732
tri 258 1704 284 1730 sw
rect 368 1714 377 1748
rect 368 1704 396 1714
rect 253 1695 337 1704
tri 253 1676 272 1695 ne
rect 272 1676 337 1695
rect 154 1650 214 1672
rect 336 1672 337 1676
rect 354 1672 396 1704
rect 336 1650 396 1672
rect 242 1634 259 1648
rect 291 1634 308 1648
tri 79 1598 101 1620 se
rect 101 1613 116 1634
tri 101 1598 116 1613 nw
rect 435 1613 450 1789
tri 450 1782 463 1795 nw
rect 536 1714 551 1942
tri 73 1592 79 1598 se
rect 79 1592 88 1598
rect 73 1576 88 1592
tri 88 1585 101 1598 nw
rect 242 1590 259 1604
rect 291 1590 308 1604
tri 435 1598 450 1613 ne
tri 450 1598 472 1620 sw
rect 73 1540 88 1548
rect 154 1576 214 1590
rect 169 1566 214 1576
rect 169 1548 197 1566
tri 73 1525 88 1540 ne
tri 88 1525 110 1547 sw
rect 154 1538 197 1548
rect 212 1562 214 1566
rect 336 1576 396 1590
tri 450 1585 463 1598 ne
rect 463 1592 472 1598
tri 472 1592 478 1598 sw
rect 336 1566 381 1576
rect 212 1538 286 1562
rect 154 1534 286 1538
tri 286 1534 314 1562 sw
rect 336 1552 338 1566
tri 336 1550 338 1552 ne
rect 350 1548 381 1566
rect 350 1538 396 1548
rect 463 1577 478 1592
tri 88 1513 100 1525 ne
rect 100 1520 110 1525
tri 110 1520 115 1525 sw
rect -1 1174 14 1402
rect 100 1364 115 1520
rect 154 1478 182 1534
tri 274 1516 292 1534 ne
rect 292 1514 314 1534
tri 314 1514 334 1534 sw
tri 350 1520 368 1538 ne
rect 173 1444 182 1478
rect 216 1505 258 1506
rect 216 1471 221 1505
rect 251 1471 258 1505
rect 216 1462 258 1471
rect 292 1505 334 1514
rect 292 1471 299 1505
rect 329 1471 334 1505
rect 292 1466 334 1471
rect 368 1478 396 1538
tri 441 1525 463 1547 se
rect 463 1540 478 1548
tri 463 1525 478 1540 nw
tri 435 1519 441 1525 se
rect 441 1519 450 1525
rect 154 1434 182 1444
tri 182 1434 206 1458 sw
rect 154 1402 196 1434
tri 213 1426 214 1427 sw
rect 213 1402 214 1426
tri 216 1425 253 1462 ne
rect 253 1434 258 1462
tri 258 1434 284 1460 sw
rect 368 1444 377 1478
rect 368 1434 396 1444
rect 253 1425 337 1434
tri 253 1406 272 1425 ne
rect 272 1406 337 1425
rect 154 1380 214 1402
rect 336 1402 337 1406
rect 354 1402 396 1434
rect 336 1380 396 1402
rect 242 1364 259 1378
rect 291 1364 308 1378
tri 79 1328 101 1350 se
rect 101 1343 116 1364
tri 101 1328 116 1343 nw
rect 435 1343 450 1519
tri 450 1512 463 1525 nw
rect 536 1444 551 1672
tri 73 1322 79 1328 se
rect 79 1322 88 1328
rect 73 1306 88 1322
tri 88 1315 101 1328 nw
rect 242 1320 259 1334
rect 291 1320 308 1334
tri 435 1328 450 1343 ne
tri 450 1328 472 1350 sw
rect 73 1270 88 1278
rect 154 1306 214 1320
rect 169 1296 214 1306
rect 169 1278 197 1296
tri 73 1255 88 1270 ne
tri 88 1255 110 1277 sw
rect 154 1268 197 1278
rect 212 1292 214 1296
rect 336 1306 396 1320
tri 450 1315 463 1328 ne
rect 463 1322 472 1328
tri 472 1322 478 1328 sw
rect 336 1296 381 1306
rect 212 1268 286 1292
rect 154 1264 286 1268
tri 286 1264 314 1292 sw
rect 336 1282 338 1296
tri 336 1280 338 1282 ne
rect 350 1278 381 1296
rect 350 1268 396 1278
rect 463 1307 478 1322
tri 88 1243 100 1255 ne
rect 100 1250 110 1255
tri 110 1250 115 1255 sw
rect -1 904 14 1132
rect 100 1094 115 1250
rect 154 1208 182 1264
tri 274 1246 292 1264 ne
rect 292 1244 314 1264
tri 314 1244 334 1264 sw
tri 350 1250 368 1268 ne
rect 173 1174 182 1208
rect 216 1235 258 1236
rect 216 1201 221 1235
rect 251 1201 258 1235
rect 216 1192 258 1201
rect 292 1235 334 1244
rect 292 1201 299 1235
rect 329 1201 334 1235
rect 292 1196 334 1201
rect 368 1208 396 1268
tri 441 1255 463 1277 se
rect 463 1270 478 1278
tri 463 1255 478 1270 nw
tri 435 1249 441 1255 se
rect 441 1249 450 1255
rect 154 1164 182 1174
tri 182 1164 206 1188 sw
rect 154 1132 196 1164
tri 213 1156 214 1157 sw
rect 213 1132 214 1156
tri 216 1155 253 1192 ne
rect 253 1164 258 1192
tri 258 1164 284 1190 sw
rect 368 1174 377 1208
rect 368 1164 396 1174
rect 253 1155 337 1164
tri 253 1136 272 1155 ne
rect 272 1136 337 1155
rect 154 1110 214 1132
rect 336 1132 337 1136
rect 354 1132 396 1164
rect 336 1110 396 1132
rect 242 1094 259 1108
rect 291 1094 308 1108
tri 79 1058 101 1080 se
rect 101 1073 116 1094
tri 101 1058 116 1073 nw
rect 435 1073 450 1249
tri 450 1242 463 1255 nw
rect 536 1174 551 1402
tri 73 1052 79 1058 se
rect 79 1052 88 1058
rect 73 1036 88 1052
tri 88 1045 101 1058 nw
rect 242 1050 259 1064
rect 291 1050 308 1064
tri 435 1058 450 1073 ne
tri 450 1058 472 1080 sw
rect 73 1000 88 1008
rect 154 1036 214 1050
rect 169 1026 214 1036
rect 169 1008 197 1026
tri 73 985 88 1000 ne
tri 88 985 110 1007 sw
rect 154 998 197 1008
rect 212 1022 214 1026
rect 336 1036 396 1050
tri 450 1045 463 1058 ne
rect 463 1052 472 1058
tri 472 1052 478 1058 sw
rect 336 1026 381 1036
rect 212 998 286 1022
rect 154 994 286 998
tri 286 994 314 1022 sw
rect 336 1012 338 1026
tri 336 1010 338 1012 ne
rect 350 1008 381 1026
rect 350 998 396 1008
rect 463 1037 478 1052
tri 88 973 100 985 ne
rect 100 980 110 985
tri 110 980 115 985 sw
rect -1 634 14 862
rect 100 824 115 980
rect 154 938 182 994
tri 274 976 292 994 ne
rect 292 974 314 994
tri 314 974 334 994 sw
tri 350 980 368 998 ne
rect 173 904 182 938
rect 216 965 258 966
rect 216 931 221 965
rect 251 931 258 965
rect 216 922 258 931
rect 292 965 334 974
rect 292 931 299 965
rect 329 931 334 965
rect 292 926 334 931
rect 368 938 396 998
tri 441 985 463 1007 se
rect 463 1000 478 1008
tri 463 985 478 1000 nw
tri 435 979 441 985 se
rect 441 979 450 985
rect 154 894 182 904
tri 182 894 206 918 sw
rect 154 862 196 894
tri 213 886 214 887 sw
rect 213 862 214 886
tri 216 885 253 922 ne
rect 253 894 258 922
tri 258 894 284 920 sw
rect 368 904 377 938
rect 368 894 396 904
rect 253 885 337 894
tri 253 866 272 885 ne
rect 272 866 337 885
rect 154 840 214 862
rect 336 862 337 866
rect 354 862 396 894
rect 336 840 396 862
rect 242 824 259 838
rect 291 824 308 838
tri 79 788 101 810 se
rect 101 803 116 824
tri 101 788 116 803 nw
rect 435 803 450 979
tri 450 972 463 985 nw
rect 536 904 551 1132
tri 73 782 79 788 se
rect 79 782 88 788
rect 73 766 88 782
tri 88 775 101 788 nw
rect 242 780 259 794
rect 291 780 308 794
tri 435 788 450 803 ne
tri 450 788 472 810 sw
rect 73 730 88 738
rect 154 766 214 780
rect 169 756 214 766
rect 169 738 197 756
tri 73 715 88 730 ne
tri 88 715 110 737 sw
rect 154 728 197 738
rect 212 752 214 756
rect 336 766 396 780
tri 450 775 463 788 ne
rect 463 782 472 788
tri 472 782 478 788 sw
rect 336 756 381 766
rect 212 728 286 752
rect 154 724 286 728
tri 286 724 314 752 sw
rect 336 742 338 756
tri 336 740 338 742 ne
rect 350 738 381 756
rect 350 728 396 738
rect 463 767 478 782
tri 88 703 100 715 ne
rect 100 710 110 715
tri 110 710 115 715 sw
rect -1 364 14 592
rect 100 554 115 710
rect 154 668 182 724
tri 274 706 292 724 ne
rect 292 704 314 724
tri 314 704 334 724 sw
tri 350 710 368 728 ne
rect 173 634 182 668
rect 216 695 258 696
rect 216 661 221 695
rect 251 661 258 695
rect 216 652 258 661
rect 292 695 334 704
rect 292 661 299 695
rect 329 661 334 695
rect 292 656 334 661
rect 368 668 396 728
tri 441 715 463 737 se
rect 463 730 478 738
tri 463 715 478 730 nw
tri 435 709 441 715 se
rect 441 709 450 715
rect 154 624 182 634
tri 182 624 206 648 sw
rect 154 592 196 624
tri 213 616 214 617 sw
rect 213 592 214 616
tri 216 615 253 652 ne
rect 253 624 258 652
tri 258 624 284 650 sw
rect 368 634 377 668
rect 368 624 396 634
rect 253 615 337 624
tri 253 596 272 615 ne
rect 272 596 337 615
rect 154 570 214 592
rect 336 592 337 596
rect 354 592 396 624
rect 336 570 396 592
rect 242 554 259 568
rect 291 554 308 568
tri 79 518 101 540 se
rect 101 533 116 554
tri 101 518 116 533 nw
rect 435 533 450 709
tri 450 702 463 715 nw
rect 536 634 551 862
tri 73 512 79 518 se
rect 79 512 88 518
rect 73 496 88 512
tri 88 505 101 518 nw
rect 242 510 259 524
rect 291 510 308 524
tri 435 518 450 533 ne
tri 450 518 472 540 sw
rect 73 460 88 468
rect 154 496 214 510
rect 169 486 214 496
rect 169 468 197 486
tri 73 445 88 460 ne
tri 88 445 110 467 sw
rect 154 458 197 468
rect 212 482 214 486
rect 336 496 396 510
tri 450 505 463 518 ne
rect 463 512 472 518
tri 472 512 478 518 sw
rect 336 486 381 496
rect 212 458 286 482
rect 154 454 286 458
tri 286 454 314 482 sw
rect 336 472 338 486
tri 336 470 338 472 ne
rect 350 468 381 486
rect 350 458 396 468
rect 463 497 478 512
tri 88 433 100 445 ne
rect 100 440 110 445
tri 110 440 115 445 sw
rect -1 94 14 322
rect 100 284 115 440
rect 154 398 182 454
tri 274 436 292 454 ne
rect 292 434 314 454
tri 314 434 334 454 sw
tri 350 440 368 458 ne
rect 173 364 182 398
rect 216 425 258 426
rect 216 391 221 425
rect 251 391 258 425
rect 216 382 258 391
rect 292 425 334 434
rect 292 391 299 425
rect 329 391 334 425
rect 292 386 334 391
rect 368 398 396 458
tri 441 445 463 467 se
rect 463 460 478 468
tri 463 445 478 460 nw
tri 435 439 441 445 se
rect 441 439 450 445
rect 154 354 182 364
tri 182 354 206 378 sw
rect 154 322 196 354
tri 213 346 214 347 sw
rect 213 322 214 346
tri 216 345 253 382 ne
rect 253 354 258 382
tri 258 354 284 380 sw
rect 368 364 377 398
rect 368 354 396 364
rect 253 345 337 354
tri 253 326 272 345 ne
rect 272 326 337 345
rect 154 300 214 322
rect 336 322 337 326
rect 354 322 396 354
rect 336 300 396 322
rect 242 284 259 298
rect 291 284 308 298
tri 79 248 101 270 se
rect 101 263 116 284
tri 101 248 116 263 nw
rect 435 263 450 439
tri 450 432 463 445 nw
rect 536 364 551 592
tri 73 242 79 248 se
rect 79 242 88 248
rect 73 226 88 242
tri 88 235 101 248 nw
rect 242 240 259 254
rect 291 240 308 254
tri 435 248 450 263 ne
tri 450 248 472 270 sw
rect 73 190 88 198
rect 154 226 214 240
rect 169 216 214 226
rect 169 198 197 216
tri 73 175 88 190 ne
tri 88 175 110 197 sw
rect 154 188 197 198
rect 212 212 214 216
rect 336 226 396 240
tri 450 235 463 248 ne
rect 463 242 472 248
tri 472 242 478 248 sw
rect 336 216 381 226
rect 212 188 286 212
rect 154 184 286 188
tri 286 184 314 212 sw
rect 336 202 338 216
tri 336 200 338 202 ne
rect 350 198 381 216
rect 350 188 396 198
rect 463 227 478 242
tri 88 163 100 175 ne
rect 100 170 110 175
tri 110 170 115 175 sw
rect -1 -176 14 52
rect 100 14 115 170
rect 154 128 182 184
tri 274 166 292 184 ne
rect 292 164 314 184
tri 314 164 334 184 sw
tri 350 170 368 188 ne
rect 173 94 182 128
rect 216 155 258 156
rect 216 121 221 155
rect 251 121 258 155
rect 216 112 258 121
rect 292 155 334 164
rect 292 121 299 155
rect 329 121 334 155
rect 292 116 334 121
rect 368 128 396 188
tri 441 175 463 197 se
rect 463 190 478 198
tri 463 175 478 190 nw
tri 435 169 441 175 se
rect 441 169 450 175
rect 154 84 182 94
tri 182 84 206 108 sw
rect 154 52 196 84
tri 213 76 214 77 sw
rect 213 52 214 76
tri 216 75 253 112 ne
rect 253 84 258 112
tri 258 84 284 110 sw
rect 368 94 377 128
rect 368 84 396 94
rect 253 75 337 84
tri 253 56 272 75 ne
rect 272 56 337 75
rect 154 30 214 52
rect 336 52 337 56
rect 354 52 396 84
rect 336 30 396 52
rect 242 14 259 28
rect 291 14 308 28
tri 79 -22 101 0 se
rect 101 -7 116 14
tri 101 -22 116 -7 nw
rect 435 -7 450 169
tri 450 162 463 175 nw
rect 536 94 551 322
tri 73 -28 79 -22 se
rect 79 -28 88 -22
rect 73 -44 88 -28
tri 88 -35 101 -22 nw
rect 242 -30 259 -16
rect 291 -30 308 -16
tri 435 -22 450 -7 ne
tri 450 -22 472 0 sw
rect 73 -80 88 -72
rect 154 -44 214 -30
rect 169 -54 214 -44
rect 169 -72 197 -54
tri 73 -95 88 -80 ne
tri 88 -95 110 -73 sw
rect 154 -82 197 -72
rect 212 -58 214 -54
rect 336 -44 396 -30
tri 450 -35 463 -22 ne
rect 463 -28 472 -22
tri 472 -28 478 -22 sw
rect 336 -54 381 -44
rect 212 -82 286 -58
rect 154 -86 286 -82
tri 286 -86 314 -58 sw
rect 336 -68 338 -54
tri 336 -70 338 -68 ne
rect 350 -72 381 -54
rect 350 -82 396 -72
rect 463 -43 478 -28
tri 88 -107 100 -95 ne
rect 100 -100 110 -95
tri 110 -100 115 -95 sw
rect -1 -446 14 -218
rect 100 -256 115 -100
rect 154 -142 182 -86
tri 274 -104 292 -86 ne
rect 292 -106 314 -86
tri 314 -106 334 -86 sw
tri 350 -100 368 -82 ne
rect 173 -176 182 -142
rect 216 -115 258 -114
rect 216 -149 221 -115
rect 251 -149 258 -115
rect 216 -158 258 -149
rect 292 -115 334 -106
rect 292 -149 299 -115
rect 329 -149 334 -115
rect 292 -154 334 -149
rect 368 -142 396 -82
tri 441 -95 463 -73 se
rect 463 -80 478 -72
tri 463 -95 478 -80 nw
tri 435 -101 441 -95 se
rect 441 -101 450 -95
rect 154 -186 182 -176
tri 182 -186 206 -162 sw
rect 154 -218 196 -186
tri 213 -194 214 -193 sw
rect 213 -218 214 -194
tri 216 -195 253 -158 ne
rect 253 -186 258 -158
tri 258 -186 284 -160 sw
rect 368 -176 377 -142
rect 368 -186 396 -176
rect 253 -195 337 -186
tri 253 -214 272 -195 ne
rect 272 -214 337 -195
rect 154 -240 214 -218
rect 336 -218 337 -214
rect 354 -218 396 -186
rect 336 -240 396 -218
rect 242 -256 259 -242
rect 291 -256 308 -242
tri 79 -292 101 -270 se
rect 101 -277 116 -256
tri 101 -292 116 -277 nw
rect 435 -277 450 -101
tri 450 -108 463 -95 nw
rect 536 -176 551 52
tri 73 -298 79 -292 se
rect 79 -298 88 -292
rect 73 -314 88 -298
tri 88 -305 101 -292 nw
rect 242 -300 259 -286
rect 291 -300 308 -286
tri 435 -292 450 -277 ne
tri 450 -292 472 -270 sw
rect 73 -350 88 -342
rect 154 -314 214 -300
rect 169 -324 214 -314
rect 169 -342 197 -324
tri 73 -365 88 -350 ne
tri 88 -365 110 -343 sw
rect 154 -352 197 -342
rect 212 -328 214 -324
rect 336 -314 396 -300
tri 450 -305 463 -292 ne
rect 463 -298 472 -292
tri 472 -298 478 -292 sw
rect 336 -324 381 -314
rect 212 -352 286 -328
rect 154 -356 286 -352
tri 286 -356 314 -328 sw
rect 336 -338 338 -324
tri 336 -340 338 -338 ne
rect 350 -342 381 -324
rect 350 -352 396 -342
rect 463 -313 478 -298
tri 88 -377 100 -365 ne
rect 100 -370 110 -365
tri 110 -370 115 -365 sw
rect -1 -716 14 -488
rect 100 -526 115 -370
rect 154 -412 182 -356
tri 274 -374 292 -356 ne
rect 292 -376 314 -356
tri 314 -376 334 -356 sw
tri 350 -370 368 -352 ne
rect 173 -446 182 -412
rect 216 -385 258 -384
rect 216 -419 221 -385
rect 251 -419 258 -385
rect 216 -428 258 -419
rect 292 -385 334 -376
rect 292 -419 299 -385
rect 329 -419 334 -385
rect 292 -424 334 -419
rect 368 -412 396 -352
tri 441 -365 463 -343 se
rect 463 -350 478 -342
tri 463 -365 478 -350 nw
tri 435 -371 441 -365 se
rect 441 -371 450 -365
rect 154 -456 182 -446
tri 182 -456 206 -432 sw
rect 154 -488 196 -456
tri 213 -464 214 -463 sw
rect 213 -488 214 -464
tri 216 -465 253 -428 ne
rect 253 -456 258 -428
tri 258 -456 284 -430 sw
rect 368 -446 377 -412
rect 368 -456 396 -446
rect 253 -465 337 -456
tri 253 -484 272 -465 ne
rect 272 -484 337 -465
rect 154 -510 214 -488
rect 336 -488 337 -484
rect 354 -488 396 -456
rect 336 -510 396 -488
rect 242 -526 259 -512
rect 291 -526 308 -512
tri 79 -562 101 -540 se
rect 101 -547 116 -526
tri 101 -562 116 -547 nw
rect 435 -547 450 -371
tri 450 -378 463 -365 nw
rect 536 -446 551 -218
tri 73 -568 79 -562 se
rect 79 -568 88 -562
rect 73 -584 88 -568
tri 88 -575 101 -562 nw
rect 242 -570 259 -556
rect 291 -570 308 -556
tri 435 -562 450 -547 ne
tri 450 -562 472 -540 sw
rect 73 -620 88 -612
rect 154 -584 214 -570
rect 169 -594 214 -584
rect 169 -612 197 -594
tri 73 -635 88 -620 ne
tri 88 -635 110 -613 sw
rect 154 -622 197 -612
rect 212 -598 214 -594
rect 336 -584 396 -570
tri 450 -575 463 -562 ne
rect 463 -568 472 -562
tri 472 -568 478 -562 sw
rect 336 -594 381 -584
rect 212 -622 286 -598
rect 154 -626 286 -622
tri 286 -626 314 -598 sw
rect 336 -608 338 -594
tri 336 -610 338 -608 ne
rect 350 -612 381 -594
rect 350 -622 396 -612
rect 463 -583 478 -568
tri 88 -647 100 -635 ne
rect 100 -640 110 -635
tri 110 -640 115 -635 sw
rect -1 -986 14 -758
rect 100 -796 115 -640
rect 154 -682 182 -626
tri 274 -644 292 -626 ne
rect 292 -646 314 -626
tri 314 -646 334 -626 sw
tri 350 -640 368 -622 ne
rect 173 -716 182 -682
rect 216 -655 258 -654
rect 216 -689 221 -655
rect 251 -689 258 -655
rect 216 -698 258 -689
rect 292 -655 334 -646
rect 292 -689 299 -655
rect 329 -689 334 -655
rect 292 -694 334 -689
rect 368 -682 396 -622
tri 441 -635 463 -613 se
rect 463 -620 478 -612
tri 463 -635 478 -620 nw
tri 435 -641 441 -635 se
rect 441 -641 450 -635
rect 154 -726 182 -716
tri 182 -726 206 -702 sw
rect 154 -758 196 -726
tri 213 -734 214 -733 sw
rect 213 -758 214 -734
tri 216 -735 253 -698 ne
rect 253 -726 258 -698
tri 258 -726 284 -700 sw
rect 368 -716 377 -682
rect 368 -726 396 -716
rect 253 -735 337 -726
tri 253 -754 272 -735 ne
rect 272 -754 337 -735
rect 154 -780 214 -758
rect 336 -758 337 -754
rect 354 -758 396 -726
rect 336 -780 396 -758
rect 242 -796 259 -782
rect 291 -796 308 -782
tri 79 -832 101 -810 se
rect 101 -817 116 -796
tri 101 -832 116 -817 nw
rect 435 -817 450 -641
tri 450 -648 463 -635 nw
rect 536 -716 551 -488
tri 73 -838 79 -832 se
rect 79 -838 88 -832
rect 73 -854 88 -838
tri 88 -845 101 -832 nw
rect 242 -840 259 -826
rect 291 -840 308 -826
tri 435 -832 450 -817 ne
tri 450 -832 472 -810 sw
rect 73 -890 88 -882
rect 154 -854 214 -840
rect 169 -864 214 -854
rect 169 -882 197 -864
tri 73 -905 88 -890 ne
tri 88 -905 110 -883 sw
rect 154 -892 197 -882
rect 212 -868 214 -864
rect 336 -854 396 -840
tri 450 -845 463 -832 ne
rect 463 -838 472 -832
tri 472 -838 478 -832 sw
rect 336 -864 381 -854
rect 212 -892 286 -868
rect 154 -896 286 -892
tri 286 -896 314 -868 sw
rect 336 -878 338 -864
tri 336 -880 338 -878 ne
rect 350 -882 381 -864
rect 350 -892 396 -882
rect 463 -853 478 -838
tri 88 -917 100 -905 ne
rect 100 -910 110 -905
tri 110 -910 115 -905 sw
rect -1 -1256 14 -1028
rect 100 -1066 115 -910
rect 154 -952 182 -896
tri 274 -914 292 -896 ne
rect 292 -916 314 -896
tri 314 -916 334 -896 sw
tri 350 -910 368 -892 ne
rect 173 -986 182 -952
rect 216 -925 258 -924
rect 216 -959 221 -925
rect 251 -959 258 -925
rect 216 -968 258 -959
rect 292 -925 334 -916
rect 292 -959 299 -925
rect 329 -959 334 -925
rect 292 -964 334 -959
rect 368 -952 396 -892
tri 441 -905 463 -883 se
rect 463 -890 478 -882
tri 463 -905 478 -890 nw
tri 435 -911 441 -905 se
rect 441 -911 450 -905
rect 154 -996 182 -986
tri 182 -996 206 -972 sw
rect 154 -1028 196 -996
tri 213 -1004 214 -1003 sw
rect 213 -1028 214 -1004
tri 216 -1005 253 -968 ne
rect 253 -996 258 -968
tri 258 -996 284 -970 sw
rect 368 -986 377 -952
rect 368 -996 396 -986
rect 253 -1005 337 -996
tri 253 -1024 272 -1005 ne
rect 272 -1024 337 -1005
rect 154 -1050 214 -1028
rect 336 -1028 337 -1024
rect 354 -1028 396 -996
rect 336 -1050 396 -1028
rect 242 -1066 259 -1052
rect 291 -1066 308 -1052
tri 79 -1102 101 -1080 se
rect 101 -1087 116 -1066
tri 101 -1102 116 -1087 nw
rect 435 -1087 450 -911
tri 450 -918 463 -905 nw
rect 536 -986 551 -758
tri 73 -1108 79 -1102 se
rect 79 -1108 88 -1102
rect 73 -1124 88 -1108
tri 88 -1115 101 -1102 nw
rect 242 -1110 259 -1096
rect 291 -1110 308 -1096
tri 435 -1102 450 -1087 ne
tri 450 -1102 472 -1080 sw
rect 73 -1160 88 -1152
rect 154 -1124 214 -1110
rect 169 -1134 214 -1124
rect 169 -1152 197 -1134
tri 73 -1175 88 -1160 ne
tri 88 -1175 110 -1153 sw
rect 154 -1162 197 -1152
rect 212 -1138 214 -1134
rect 336 -1124 396 -1110
tri 450 -1115 463 -1102 ne
rect 463 -1108 472 -1102
tri 472 -1108 478 -1102 sw
rect 336 -1134 381 -1124
rect 212 -1162 286 -1138
rect 154 -1166 286 -1162
tri 286 -1166 314 -1138 sw
rect 336 -1148 338 -1134
tri 336 -1150 338 -1148 ne
rect 350 -1152 381 -1134
rect 350 -1162 396 -1152
rect 463 -1123 478 -1108
tri 88 -1187 100 -1175 ne
rect 100 -1180 110 -1175
tri 110 -1180 115 -1175 sw
rect -1 -1526 14 -1298
rect 100 -1336 115 -1180
rect 154 -1222 182 -1166
tri 274 -1184 292 -1166 ne
rect 292 -1186 314 -1166
tri 314 -1186 334 -1166 sw
tri 350 -1180 368 -1162 ne
rect 173 -1256 182 -1222
rect 216 -1195 258 -1194
rect 216 -1229 221 -1195
rect 251 -1229 258 -1195
rect 216 -1238 258 -1229
rect 292 -1195 334 -1186
rect 292 -1229 299 -1195
rect 329 -1229 334 -1195
rect 292 -1234 334 -1229
rect 368 -1222 396 -1162
tri 441 -1175 463 -1153 se
rect 463 -1160 478 -1152
tri 463 -1175 478 -1160 nw
tri 435 -1181 441 -1175 se
rect 441 -1181 450 -1175
rect 154 -1266 182 -1256
tri 182 -1266 206 -1242 sw
rect 154 -1298 196 -1266
tri 213 -1274 214 -1273 sw
rect 213 -1298 214 -1274
tri 216 -1275 253 -1238 ne
rect 253 -1266 258 -1238
tri 258 -1266 284 -1240 sw
rect 368 -1256 377 -1222
rect 368 -1266 396 -1256
rect 253 -1275 337 -1266
tri 253 -1294 272 -1275 ne
rect 272 -1294 337 -1275
rect 154 -1320 214 -1298
rect 336 -1298 337 -1294
rect 354 -1298 396 -1266
rect 336 -1320 396 -1298
rect 242 -1336 259 -1322
rect 291 -1336 308 -1322
tri 79 -1372 101 -1350 se
rect 101 -1357 116 -1336
tri 101 -1372 116 -1357 nw
rect 435 -1357 450 -1181
tri 450 -1188 463 -1175 nw
rect 536 -1256 551 -1028
tri 73 -1378 79 -1372 se
rect 79 -1378 88 -1372
rect 73 -1394 88 -1378
tri 88 -1385 101 -1372 nw
rect 242 -1380 259 -1366
rect 291 -1380 308 -1366
tri 435 -1372 450 -1357 ne
tri 450 -1372 472 -1350 sw
rect 73 -1430 88 -1422
rect 154 -1394 214 -1380
rect 169 -1404 214 -1394
rect 169 -1422 197 -1404
tri 73 -1445 88 -1430 ne
tri 88 -1445 110 -1423 sw
rect 154 -1432 197 -1422
rect 212 -1408 214 -1404
rect 336 -1394 396 -1380
tri 450 -1385 463 -1372 ne
rect 463 -1378 472 -1372
tri 472 -1378 478 -1372 sw
rect 336 -1404 381 -1394
rect 212 -1432 286 -1408
rect 154 -1436 286 -1432
tri 286 -1436 314 -1408 sw
rect 336 -1418 338 -1404
tri 336 -1420 338 -1418 ne
rect 350 -1422 381 -1404
rect 350 -1432 396 -1422
rect 463 -1393 478 -1378
tri 88 -1457 100 -1445 ne
rect 100 -1450 110 -1445
tri 110 -1450 115 -1445 sw
rect -1 -1796 14 -1568
rect 100 -1606 115 -1450
rect 154 -1492 182 -1436
tri 274 -1454 292 -1436 ne
rect 292 -1456 314 -1436
tri 314 -1456 334 -1436 sw
tri 350 -1450 368 -1432 ne
rect 173 -1526 182 -1492
rect 216 -1465 258 -1464
rect 216 -1499 221 -1465
rect 251 -1499 258 -1465
rect 216 -1508 258 -1499
rect 292 -1465 334 -1456
rect 292 -1499 299 -1465
rect 329 -1499 334 -1465
rect 292 -1504 334 -1499
rect 368 -1492 396 -1432
tri 441 -1445 463 -1423 se
rect 463 -1430 478 -1422
tri 463 -1445 478 -1430 nw
tri 435 -1451 441 -1445 se
rect 441 -1451 450 -1445
rect 154 -1536 182 -1526
tri 182 -1536 206 -1512 sw
rect 154 -1568 196 -1536
tri 213 -1544 214 -1543 sw
rect 213 -1568 214 -1544
tri 216 -1545 253 -1508 ne
rect 253 -1536 258 -1508
tri 258 -1536 284 -1510 sw
rect 368 -1526 377 -1492
rect 368 -1536 396 -1526
rect 253 -1545 337 -1536
tri 253 -1564 272 -1545 ne
rect 272 -1564 337 -1545
rect 154 -1590 214 -1568
rect 336 -1568 337 -1564
rect 354 -1568 396 -1536
rect 336 -1590 396 -1568
rect 242 -1606 259 -1592
rect 291 -1606 308 -1592
tri 79 -1642 101 -1620 se
rect 101 -1627 116 -1606
tri 101 -1642 116 -1627 nw
rect 435 -1627 450 -1451
tri 450 -1458 463 -1445 nw
rect 536 -1526 551 -1298
tri 73 -1648 79 -1642 se
rect 79 -1648 88 -1642
rect 73 -1664 88 -1648
tri 88 -1655 101 -1642 nw
rect 242 -1650 259 -1636
rect 291 -1650 308 -1636
tri 435 -1642 450 -1627 ne
tri 450 -1642 472 -1620 sw
rect 73 -1700 88 -1692
rect 154 -1664 214 -1650
rect 169 -1674 214 -1664
rect 169 -1692 197 -1674
tri 73 -1715 88 -1700 ne
tri 88 -1715 110 -1693 sw
rect 154 -1702 197 -1692
rect 212 -1678 214 -1674
rect 336 -1664 396 -1650
tri 450 -1655 463 -1642 ne
rect 463 -1648 472 -1642
tri 472 -1648 478 -1642 sw
rect 336 -1674 381 -1664
rect 212 -1702 286 -1678
rect 154 -1706 286 -1702
tri 286 -1706 314 -1678 sw
rect 336 -1688 338 -1674
tri 336 -1690 338 -1688 ne
rect 350 -1692 381 -1674
rect 350 -1702 396 -1692
rect 463 -1663 478 -1648
tri 88 -1727 100 -1715 ne
rect 100 -1720 110 -1715
tri 110 -1720 115 -1715 sw
rect -1 -2066 14 -1838
rect 100 -1876 115 -1720
rect 154 -1762 182 -1706
tri 274 -1724 292 -1706 ne
rect 292 -1726 314 -1706
tri 314 -1726 334 -1706 sw
tri 350 -1720 368 -1702 ne
rect 173 -1796 182 -1762
rect 216 -1735 258 -1734
rect 216 -1769 221 -1735
rect 251 -1769 258 -1735
rect 216 -1778 258 -1769
rect 292 -1735 334 -1726
rect 292 -1769 299 -1735
rect 329 -1769 334 -1735
rect 292 -1774 334 -1769
rect 368 -1762 396 -1702
tri 441 -1715 463 -1693 se
rect 463 -1700 478 -1692
tri 463 -1715 478 -1700 nw
tri 435 -1721 441 -1715 se
rect 441 -1721 450 -1715
rect 154 -1806 182 -1796
tri 182 -1806 206 -1782 sw
rect 154 -1838 196 -1806
tri 213 -1814 214 -1813 sw
rect 213 -1838 214 -1814
tri 216 -1815 253 -1778 ne
rect 253 -1806 258 -1778
tri 258 -1806 284 -1780 sw
rect 368 -1796 377 -1762
rect 368 -1806 396 -1796
rect 253 -1815 337 -1806
tri 253 -1834 272 -1815 ne
rect 272 -1834 337 -1815
rect 154 -1860 214 -1838
rect 336 -1838 337 -1834
rect 354 -1838 396 -1806
rect 336 -1860 396 -1838
rect 242 -1876 259 -1862
rect 291 -1876 308 -1862
tri 79 -1912 101 -1890 se
rect 101 -1897 116 -1876
tri 101 -1912 116 -1897 nw
rect 435 -1897 450 -1721
tri 450 -1728 463 -1715 nw
rect 536 -1796 551 -1568
tri 73 -1918 79 -1912 se
rect 79 -1918 88 -1912
rect 73 -1934 88 -1918
tri 88 -1925 101 -1912 nw
rect 242 -1920 259 -1906
rect 291 -1920 308 -1906
tri 435 -1912 450 -1897 ne
tri 450 -1912 472 -1890 sw
rect 73 -1970 88 -1962
rect 154 -1934 214 -1920
rect 169 -1944 214 -1934
rect 169 -1962 197 -1944
tri 73 -1985 88 -1970 ne
tri 88 -1985 110 -1963 sw
rect 154 -1972 197 -1962
rect 212 -1948 214 -1944
rect 336 -1934 396 -1920
tri 450 -1925 463 -1912 ne
rect 463 -1918 472 -1912
tri 472 -1918 478 -1912 sw
rect 336 -1944 381 -1934
rect 212 -1972 286 -1948
rect 154 -1976 286 -1972
tri 286 -1976 314 -1948 sw
rect 336 -1958 338 -1944
tri 336 -1960 338 -1958 ne
rect 350 -1962 381 -1944
rect 350 -1972 396 -1962
rect 463 -1933 478 -1918
tri 88 -1997 100 -1985 ne
rect 100 -1990 110 -1985
tri 110 -1990 115 -1985 sw
rect -1 -2146 14 -2108
rect 100 -2146 115 -1990
rect 154 -2032 182 -1976
tri 274 -1994 292 -1976 ne
rect 292 -1996 314 -1976
tri 314 -1996 334 -1976 sw
tri 350 -1990 368 -1972 ne
rect 173 -2066 182 -2032
rect 216 -2005 258 -2004
rect 216 -2039 221 -2005
rect 251 -2039 258 -2005
rect 216 -2048 258 -2039
rect 292 -2005 334 -1996
rect 292 -2039 299 -2005
rect 329 -2039 334 -2005
rect 292 -2044 334 -2039
rect 368 -2032 396 -1972
tri 441 -1985 463 -1963 se
rect 463 -1970 478 -1962
tri 463 -1985 478 -1970 nw
tri 435 -1991 441 -1985 se
rect 441 -1991 450 -1985
rect 154 -2076 182 -2066
tri 182 -2076 206 -2052 sw
rect 154 -2108 196 -2076
tri 213 -2084 214 -2083 sw
rect 213 -2108 214 -2084
tri 216 -2085 253 -2048 ne
rect 253 -2076 258 -2048
tri 258 -2076 284 -2050 sw
rect 368 -2066 377 -2032
rect 368 -2076 396 -2066
rect 253 -2085 337 -2076
tri 253 -2104 272 -2085 ne
rect 272 -2104 337 -2085
rect 154 -2130 214 -2108
rect 336 -2108 337 -2104
rect 354 -2108 396 -2076
rect 336 -2130 396 -2108
rect 242 -2146 259 -2132
rect 291 -2146 308 -2132
rect 435 -2146 450 -1991
tri 450 -1998 463 -1985 nw
rect 536 -2066 551 -1838
rect 536 -2146 551 -2108
rect 579 1984 594 2174
tri 659 2138 681 2160 se
rect 681 2153 696 2174
tri 681 2138 696 2153 nw
rect 1015 2153 1030 2174
tri 653 2132 659 2138 se
rect 659 2132 668 2138
rect 653 2116 668 2132
tri 668 2125 681 2138 nw
rect 822 2130 839 2144
rect 871 2130 888 2144
tri 1015 2138 1030 2153 ne
tri 1030 2138 1052 2160 sw
rect 653 2080 668 2088
rect 734 2116 794 2130
rect 749 2106 794 2116
rect 749 2088 777 2106
tri 653 2065 668 2080 ne
tri 668 2065 690 2087 sw
rect 734 2078 777 2088
rect 792 2102 794 2106
rect 916 2116 976 2130
tri 1030 2125 1043 2138 ne
rect 1043 2132 1052 2138
tri 1052 2132 1058 2138 sw
rect 916 2106 961 2116
rect 792 2078 866 2102
rect 734 2074 866 2078
tri 866 2074 894 2102 sw
rect 916 2092 918 2106
tri 916 2090 918 2092 ne
rect 930 2088 961 2106
rect 930 2078 976 2088
rect 1043 2117 1058 2132
tri 668 2053 680 2065 ne
rect 680 2060 690 2065
tri 690 2060 695 2065 sw
rect 579 1714 594 1942
rect 680 1904 695 2060
rect 734 2018 762 2074
tri 854 2056 872 2074 ne
rect 872 2054 894 2074
tri 894 2054 914 2074 sw
tri 930 2060 948 2078 ne
rect 753 1984 762 2018
rect 796 2045 838 2046
rect 796 2011 801 2045
rect 831 2011 838 2045
rect 796 2002 838 2011
rect 872 2045 914 2054
rect 872 2011 879 2045
rect 909 2011 914 2045
rect 872 2006 914 2011
rect 948 2018 976 2078
tri 1021 2065 1043 2087 se
rect 1043 2080 1058 2088
tri 1043 2065 1058 2080 nw
tri 1015 2059 1021 2065 se
rect 1021 2059 1030 2065
rect 734 1974 762 1984
tri 762 1974 786 1998 sw
rect 734 1942 776 1974
tri 793 1966 794 1967 sw
rect 793 1942 794 1966
tri 796 1965 833 2002 ne
rect 833 1974 838 2002
tri 838 1974 864 2000 sw
rect 948 1984 957 2018
rect 948 1974 976 1984
rect 833 1965 917 1974
tri 833 1946 852 1965 ne
rect 852 1946 917 1965
rect 734 1920 794 1942
rect 916 1942 917 1946
rect 934 1942 976 1974
rect 916 1920 976 1942
rect 822 1904 839 1918
rect 871 1904 888 1918
tri 659 1868 681 1890 se
rect 681 1883 696 1904
tri 681 1868 696 1883 nw
rect 1015 1883 1030 2059
tri 1030 2052 1043 2065 nw
rect 1116 1984 1131 2174
tri 653 1862 659 1868 se
rect 659 1862 668 1868
rect 653 1846 668 1862
tri 668 1855 681 1868 nw
rect 822 1860 839 1874
rect 871 1860 888 1874
tri 1015 1868 1030 1883 ne
tri 1030 1868 1052 1890 sw
rect 653 1810 668 1818
rect 734 1846 794 1860
rect 749 1836 794 1846
rect 749 1818 777 1836
tri 653 1795 668 1810 ne
tri 668 1795 690 1817 sw
rect 734 1808 777 1818
rect 792 1832 794 1836
rect 916 1846 976 1860
tri 1030 1855 1043 1868 ne
rect 1043 1862 1052 1868
tri 1052 1862 1058 1868 sw
rect 916 1836 961 1846
rect 792 1808 866 1832
rect 734 1804 866 1808
tri 866 1804 894 1832 sw
rect 916 1822 918 1836
tri 916 1820 918 1822 ne
rect 930 1818 961 1836
rect 930 1808 976 1818
rect 1043 1847 1058 1862
tri 668 1783 680 1795 ne
rect 680 1790 690 1795
tri 690 1790 695 1795 sw
rect 579 1444 594 1672
rect 680 1634 695 1790
rect 734 1748 762 1804
tri 854 1786 872 1804 ne
rect 872 1784 894 1804
tri 894 1784 914 1804 sw
tri 930 1790 948 1808 ne
rect 753 1714 762 1748
rect 796 1775 838 1776
rect 796 1741 801 1775
rect 831 1741 838 1775
rect 796 1732 838 1741
rect 872 1775 914 1784
rect 872 1741 879 1775
rect 909 1741 914 1775
rect 872 1736 914 1741
rect 948 1748 976 1808
tri 1021 1795 1043 1817 se
rect 1043 1810 1058 1818
tri 1043 1795 1058 1810 nw
tri 1015 1789 1021 1795 se
rect 1021 1789 1030 1795
rect 734 1704 762 1714
tri 762 1704 786 1728 sw
rect 734 1672 776 1704
tri 793 1696 794 1697 sw
rect 793 1672 794 1696
tri 796 1695 833 1732 ne
rect 833 1704 838 1732
tri 838 1704 864 1730 sw
rect 948 1714 957 1748
rect 948 1704 976 1714
rect 833 1695 917 1704
tri 833 1676 852 1695 ne
rect 852 1676 917 1695
rect 734 1650 794 1672
rect 916 1672 917 1676
rect 934 1672 976 1704
rect 916 1650 976 1672
rect 822 1634 839 1648
rect 871 1634 888 1648
tri 659 1598 681 1620 se
rect 681 1613 696 1634
tri 681 1598 696 1613 nw
rect 1015 1613 1030 1789
tri 1030 1782 1043 1795 nw
rect 1116 1714 1131 1942
tri 653 1592 659 1598 se
rect 659 1592 668 1598
rect 653 1576 668 1592
tri 668 1585 681 1598 nw
rect 822 1590 839 1604
rect 871 1590 888 1604
tri 1015 1598 1030 1613 ne
tri 1030 1598 1052 1620 sw
rect 653 1540 668 1548
rect 734 1576 794 1590
rect 749 1566 794 1576
rect 749 1548 777 1566
tri 653 1525 668 1540 ne
tri 668 1525 690 1547 sw
rect 734 1538 777 1548
rect 792 1562 794 1566
rect 916 1576 976 1590
tri 1030 1585 1043 1598 ne
rect 1043 1592 1052 1598
tri 1052 1592 1058 1598 sw
rect 916 1566 961 1576
rect 792 1538 866 1562
rect 734 1534 866 1538
tri 866 1534 894 1562 sw
rect 916 1552 918 1566
tri 916 1550 918 1552 ne
rect 930 1548 961 1566
rect 930 1538 976 1548
rect 1043 1577 1058 1592
tri 668 1513 680 1525 ne
rect 680 1520 690 1525
tri 690 1520 695 1525 sw
rect 579 1174 594 1402
rect 680 1364 695 1520
rect 734 1478 762 1534
tri 854 1516 872 1534 ne
rect 872 1514 894 1534
tri 894 1514 914 1534 sw
tri 930 1520 948 1538 ne
rect 753 1444 762 1478
rect 796 1505 838 1506
rect 796 1471 801 1505
rect 831 1471 838 1505
rect 796 1462 838 1471
rect 872 1505 914 1514
rect 872 1471 879 1505
rect 909 1471 914 1505
rect 872 1466 914 1471
rect 948 1478 976 1538
tri 1021 1525 1043 1547 se
rect 1043 1540 1058 1548
tri 1043 1525 1058 1540 nw
tri 1015 1519 1021 1525 se
rect 1021 1519 1030 1525
rect 734 1434 762 1444
tri 762 1434 786 1458 sw
rect 734 1402 776 1434
tri 793 1426 794 1427 sw
rect 793 1402 794 1426
tri 796 1425 833 1462 ne
rect 833 1434 838 1462
tri 838 1434 864 1460 sw
rect 948 1444 957 1478
rect 948 1434 976 1444
rect 833 1425 917 1434
tri 833 1406 852 1425 ne
rect 852 1406 917 1425
rect 734 1380 794 1402
rect 916 1402 917 1406
rect 934 1402 976 1434
rect 916 1380 976 1402
rect 822 1364 839 1378
rect 871 1364 888 1378
tri 659 1328 681 1350 se
rect 681 1343 696 1364
tri 681 1328 696 1343 nw
rect 1015 1343 1030 1519
tri 1030 1512 1043 1525 nw
rect 1116 1444 1131 1672
tri 653 1322 659 1328 se
rect 659 1322 668 1328
rect 653 1306 668 1322
tri 668 1315 681 1328 nw
rect 822 1320 839 1334
rect 871 1320 888 1334
tri 1015 1328 1030 1343 ne
tri 1030 1328 1052 1350 sw
rect 653 1270 668 1278
rect 734 1306 794 1320
rect 749 1296 794 1306
rect 749 1278 777 1296
tri 653 1255 668 1270 ne
tri 668 1255 690 1277 sw
rect 734 1268 777 1278
rect 792 1292 794 1296
rect 916 1306 976 1320
tri 1030 1315 1043 1328 ne
rect 1043 1322 1052 1328
tri 1052 1322 1058 1328 sw
rect 916 1296 961 1306
rect 792 1268 866 1292
rect 734 1264 866 1268
tri 866 1264 894 1292 sw
rect 916 1282 918 1296
tri 916 1280 918 1282 ne
rect 930 1278 961 1296
rect 930 1268 976 1278
rect 1043 1307 1058 1322
tri 668 1243 680 1255 ne
rect 680 1250 690 1255
tri 690 1250 695 1255 sw
rect 579 904 594 1132
rect 680 1094 695 1250
rect 734 1208 762 1264
tri 854 1246 872 1264 ne
rect 872 1244 894 1264
tri 894 1244 914 1264 sw
tri 930 1250 948 1268 ne
rect 753 1174 762 1208
rect 796 1235 838 1236
rect 796 1201 801 1235
rect 831 1201 838 1235
rect 796 1192 838 1201
rect 872 1235 914 1244
rect 872 1201 879 1235
rect 909 1201 914 1235
rect 872 1196 914 1201
rect 948 1208 976 1268
tri 1021 1255 1043 1277 se
rect 1043 1270 1058 1278
tri 1043 1255 1058 1270 nw
tri 1015 1249 1021 1255 se
rect 1021 1249 1030 1255
rect 734 1164 762 1174
tri 762 1164 786 1188 sw
rect 734 1132 776 1164
tri 793 1156 794 1157 sw
rect 793 1132 794 1156
tri 796 1155 833 1192 ne
rect 833 1164 838 1192
tri 838 1164 864 1190 sw
rect 948 1174 957 1208
rect 948 1164 976 1174
rect 833 1155 917 1164
tri 833 1136 852 1155 ne
rect 852 1136 917 1155
rect 734 1110 794 1132
rect 916 1132 917 1136
rect 934 1132 976 1164
rect 916 1110 976 1132
rect 822 1094 839 1108
rect 871 1094 888 1108
tri 659 1058 681 1080 se
rect 681 1073 696 1094
tri 681 1058 696 1073 nw
rect 1015 1073 1030 1249
tri 1030 1242 1043 1255 nw
rect 1116 1174 1131 1402
tri 653 1052 659 1058 se
rect 659 1052 668 1058
rect 653 1036 668 1052
tri 668 1045 681 1058 nw
rect 822 1050 839 1064
rect 871 1050 888 1064
tri 1015 1058 1030 1073 ne
tri 1030 1058 1052 1080 sw
rect 653 1000 668 1008
rect 734 1036 794 1050
rect 749 1026 794 1036
rect 749 1008 777 1026
tri 653 985 668 1000 ne
tri 668 985 690 1007 sw
rect 734 998 777 1008
rect 792 1022 794 1026
rect 916 1036 976 1050
tri 1030 1045 1043 1058 ne
rect 1043 1052 1052 1058
tri 1052 1052 1058 1058 sw
rect 916 1026 961 1036
rect 792 998 866 1022
rect 734 994 866 998
tri 866 994 894 1022 sw
rect 916 1012 918 1026
tri 916 1010 918 1012 ne
rect 930 1008 961 1026
rect 930 998 976 1008
rect 1043 1037 1058 1052
tri 668 973 680 985 ne
rect 680 980 690 985
tri 690 980 695 985 sw
rect 579 634 594 862
rect 680 824 695 980
rect 734 938 762 994
tri 854 976 872 994 ne
rect 872 974 894 994
tri 894 974 914 994 sw
tri 930 980 948 998 ne
rect 753 904 762 938
rect 796 965 838 966
rect 796 931 801 965
rect 831 931 838 965
rect 796 922 838 931
rect 872 965 914 974
rect 872 931 879 965
rect 909 931 914 965
rect 872 926 914 931
rect 948 938 976 998
tri 1021 985 1043 1007 se
rect 1043 1000 1058 1008
tri 1043 985 1058 1000 nw
tri 1015 979 1021 985 se
rect 1021 979 1030 985
rect 734 894 762 904
tri 762 894 786 918 sw
rect 734 862 776 894
tri 793 886 794 887 sw
rect 793 862 794 886
tri 796 885 833 922 ne
rect 833 894 838 922
tri 838 894 864 920 sw
rect 948 904 957 938
rect 948 894 976 904
rect 833 885 917 894
tri 833 866 852 885 ne
rect 852 866 917 885
rect 734 840 794 862
rect 916 862 917 866
rect 934 862 976 894
rect 916 840 976 862
rect 822 824 839 838
rect 871 824 888 838
tri 659 788 681 810 se
rect 681 803 696 824
tri 681 788 696 803 nw
rect 1015 803 1030 979
tri 1030 972 1043 985 nw
rect 1116 904 1131 1132
tri 653 782 659 788 se
rect 659 782 668 788
rect 653 766 668 782
tri 668 775 681 788 nw
rect 822 780 839 794
rect 871 780 888 794
tri 1015 788 1030 803 ne
tri 1030 788 1052 810 sw
rect 653 730 668 738
rect 734 766 794 780
rect 749 756 794 766
rect 749 738 777 756
tri 653 715 668 730 ne
tri 668 715 690 737 sw
rect 734 728 777 738
rect 792 752 794 756
rect 916 766 976 780
tri 1030 775 1043 788 ne
rect 1043 782 1052 788
tri 1052 782 1058 788 sw
rect 916 756 961 766
rect 792 728 866 752
rect 734 724 866 728
tri 866 724 894 752 sw
rect 916 742 918 756
tri 916 740 918 742 ne
rect 930 738 961 756
rect 930 728 976 738
rect 1043 767 1058 782
tri 668 703 680 715 ne
rect 680 710 690 715
tri 690 710 695 715 sw
rect 579 364 594 592
rect 680 554 695 710
rect 734 668 762 724
tri 854 706 872 724 ne
rect 872 704 894 724
tri 894 704 914 724 sw
tri 930 710 948 728 ne
rect 753 634 762 668
rect 796 695 838 696
rect 796 661 801 695
rect 831 661 838 695
rect 796 652 838 661
rect 872 695 914 704
rect 872 661 879 695
rect 909 661 914 695
rect 872 656 914 661
rect 948 668 976 728
tri 1021 715 1043 737 se
rect 1043 730 1058 738
tri 1043 715 1058 730 nw
tri 1015 709 1021 715 se
rect 1021 709 1030 715
rect 734 624 762 634
tri 762 624 786 648 sw
rect 734 592 776 624
tri 793 616 794 617 sw
rect 793 592 794 616
tri 796 615 833 652 ne
rect 833 624 838 652
tri 838 624 864 650 sw
rect 948 634 957 668
rect 948 624 976 634
rect 833 615 917 624
tri 833 596 852 615 ne
rect 852 596 917 615
rect 734 570 794 592
rect 916 592 917 596
rect 934 592 976 624
rect 916 570 976 592
rect 822 554 839 568
rect 871 554 888 568
tri 659 518 681 540 se
rect 681 533 696 554
tri 681 518 696 533 nw
rect 1015 533 1030 709
tri 1030 702 1043 715 nw
rect 1116 634 1131 862
tri 653 512 659 518 se
rect 659 512 668 518
rect 653 496 668 512
tri 668 505 681 518 nw
rect 822 510 839 524
rect 871 510 888 524
tri 1015 518 1030 533 ne
tri 1030 518 1052 540 sw
rect 653 460 668 468
rect 734 496 794 510
rect 749 486 794 496
rect 749 468 777 486
tri 653 445 668 460 ne
tri 668 445 690 467 sw
rect 734 458 777 468
rect 792 482 794 486
rect 916 496 976 510
tri 1030 505 1043 518 ne
rect 1043 512 1052 518
tri 1052 512 1058 518 sw
rect 916 486 961 496
rect 792 458 866 482
rect 734 454 866 458
tri 866 454 894 482 sw
rect 916 472 918 486
tri 916 470 918 472 ne
rect 930 468 961 486
rect 930 458 976 468
rect 1043 497 1058 512
tri 668 433 680 445 ne
rect 680 440 690 445
tri 690 440 695 445 sw
rect 579 94 594 322
rect 680 284 695 440
rect 734 398 762 454
tri 854 436 872 454 ne
rect 872 434 894 454
tri 894 434 914 454 sw
tri 930 440 948 458 ne
rect 753 364 762 398
rect 796 425 838 426
rect 796 391 801 425
rect 831 391 838 425
rect 796 382 838 391
rect 872 425 914 434
rect 872 391 879 425
rect 909 391 914 425
rect 872 386 914 391
rect 948 398 976 458
tri 1021 445 1043 467 se
rect 1043 460 1058 468
tri 1043 445 1058 460 nw
tri 1015 439 1021 445 se
rect 1021 439 1030 445
rect 734 354 762 364
tri 762 354 786 378 sw
rect 734 322 776 354
tri 793 346 794 347 sw
rect 793 322 794 346
tri 796 345 833 382 ne
rect 833 354 838 382
tri 838 354 864 380 sw
rect 948 364 957 398
rect 948 354 976 364
rect 833 345 917 354
tri 833 326 852 345 ne
rect 852 326 917 345
rect 734 300 794 322
rect 916 322 917 326
rect 934 322 976 354
rect 916 300 976 322
rect 822 284 839 298
rect 871 284 888 298
tri 659 248 681 270 se
rect 681 263 696 284
tri 681 248 696 263 nw
rect 1015 263 1030 439
tri 1030 432 1043 445 nw
rect 1116 364 1131 592
tri 653 242 659 248 se
rect 659 242 668 248
rect 653 226 668 242
tri 668 235 681 248 nw
rect 822 240 839 254
rect 871 240 888 254
tri 1015 248 1030 263 ne
tri 1030 248 1052 270 sw
rect 653 190 668 198
rect 734 226 794 240
rect 749 216 794 226
rect 749 198 777 216
tri 653 175 668 190 ne
tri 668 175 690 197 sw
rect 734 188 777 198
rect 792 212 794 216
rect 916 226 976 240
tri 1030 235 1043 248 ne
rect 1043 242 1052 248
tri 1052 242 1058 248 sw
rect 916 216 961 226
rect 792 188 866 212
rect 734 184 866 188
tri 866 184 894 212 sw
rect 916 202 918 216
tri 916 200 918 202 ne
rect 930 198 961 216
rect 930 188 976 198
rect 1043 227 1058 242
tri 668 163 680 175 ne
rect 680 170 690 175
tri 690 170 695 175 sw
rect 579 -176 594 52
rect 680 14 695 170
rect 734 128 762 184
tri 854 166 872 184 ne
rect 872 164 894 184
tri 894 164 914 184 sw
tri 930 170 948 188 ne
rect 753 94 762 128
rect 796 155 838 156
rect 796 121 801 155
rect 831 121 838 155
rect 796 112 838 121
rect 872 155 914 164
rect 872 121 879 155
rect 909 121 914 155
rect 872 116 914 121
rect 948 128 976 188
tri 1021 175 1043 197 se
rect 1043 190 1058 198
tri 1043 175 1058 190 nw
tri 1015 169 1021 175 se
rect 1021 169 1030 175
rect 734 84 762 94
tri 762 84 786 108 sw
rect 734 52 776 84
tri 793 76 794 77 sw
rect 793 52 794 76
tri 796 75 833 112 ne
rect 833 84 838 112
tri 838 84 864 110 sw
rect 948 94 957 128
rect 948 84 976 94
rect 833 75 917 84
tri 833 56 852 75 ne
rect 852 56 917 75
rect 734 30 794 52
rect 916 52 917 56
rect 934 52 976 84
rect 916 30 976 52
rect 822 14 839 28
rect 871 14 888 28
tri 659 -22 681 0 se
rect 681 -7 696 14
tri 681 -22 696 -7 nw
rect 1015 -7 1030 169
tri 1030 162 1043 175 nw
rect 1116 94 1131 322
tri 653 -28 659 -22 se
rect 659 -28 668 -22
rect 653 -44 668 -28
tri 668 -35 681 -22 nw
rect 822 -30 839 -16
rect 871 -30 888 -16
tri 1015 -22 1030 -7 ne
tri 1030 -22 1052 0 sw
rect 653 -80 668 -72
rect 734 -44 794 -30
rect 749 -54 794 -44
rect 749 -72 777 -54
tri 653 -95 668 -80 ne
tri 668 -95 690 -73 sw
rect 734 -82 777 -72
rect 792 -58 794 -54
rect 916 -44 976 -30
tri 1030 -35 1043 -22 ne
rect 1043 -28 1052 -22
tri 1052 -28 1058 -22 sw
rect 916 -54 961 -44
rect 792 -82 866 -58
rect 734 -86 866 -82
tri 866 -86 894 -58 sw
rect 916 -68 918 -54
tri 916 -70 918 -68 ne
rect 930 -72 961 -54
rect 930 -82 976 -72
rect 1043 -43 1058 -28
tri 668 -107 680 -95 ne
rect 680 -100 690 -95
tri 690 -100 695 -95 sw
rect 579 -446 594 -218
rect 680 -256 695 -100
rect 734 -142 762 -86
tri 854 -104 872 -86 ne
rect 872 -106 894 -86
tri 894 -106 914 -86 sw
tri 930 -100 948 -82 ne
rect 753 -176 762 -142
rect 796 -115 838 -114
rect 796 -149 801 -115
rect 831 -149 838 -115
rect 796 -158 838 -149
rect 872 -115 914 -106
rect 872 -149 879 -115
rect 909 -149 914 -115
rect 872 -154 914 -149
rect 948 -142 976 -82
tri 1021 -95 1043 -73 se
rect 1043 -80 1058 -72
tri 1043 -95 1058 -80 nw
tri 1015 -101 1021 -95 se
rect 1021 -101 1030 -95
rect 734 -186 762 -176
tri 762 -186 786 -162 sw
rect 734 -218 776 -186
tri 793 -194 794 -193 sw
rect 793 -218 794 -194
tri 796 -195 833 -158 ne
rect 833 -186 838 -158
tri 838 -186 864 -160 sw
rect 948 -176 957 -142
rect 948 -186 976 -176
rect 833 -195 917 -186
tri 833 -214 852 -195 ne
rect 852 -214 917 -195
rect 734 -240 794 -218
rect 916 -218 917 -214
rect 934 -218 976 -186
rect 916 -240 976 -218
rect 822 -256 839 -242
rect 871 -256 888 -242
tri 659 -292 681 -270 se
rect 681 -277 696 -256
tri 681 -292 696 -277 nw
rect 1015 -277 1030 -101
tri 1030 -108 1043 -95 nw
rect 1116 -176 1131 52
tri 653 -298 659 -292 se
rect 659 -298 668 -292
rect 653 -314 668 -298
tri 668 -305 681 -292 nw
rect 822 -300 839 -286
rect 871 -300 888 -286
tri 1015 -292 1030 -277 ne
tri 1030 -292 1052 -270 sw
rect 653 -350 668 -342
rect 734 -314 794 -300
rect 749 -324 794 -314
rect 749 -342 777 -324
tri 653 -365 668 -350 ne
tri 668 -365 690 -343 sw
rect 734 -352 777 -342
rect 792 -328 794 -324
rect 916 -314 976 -300
tri 1030 -305 1043 -292 ne
rect 1043 -298 1052 -292
tri 1052 -298 1058 -292 sw
rect 916 -324 961 -314
rect 792 -352 866 -328
rect 734 -356 866 -352
tri 866 -356 894 -328 sw
rect 916 -338 918 -324
tri 916 -340 918 -338 ne
rect 930 -342 961 -324
rect 930 -352 976 -342
rect 1043 -313 1058 -298
tri 668 -377 680 -365 ne
rect 680 -370 690 -365
tri 690 -370 695 -365 sw
rect 579 -716 594 -488
rect 680 -526 695 -370
rect 734 -412 762 -356
tri 854 -374 872 -356 ne
rect 872 -376 894 -356
tri 894 -376 914 -356 sw
tri 930 -370 948 -352 ne
rect 753 -446 762 -412
rect 796 -385 838 -384
rect 796 -419 801 -385
rect 831 -419 838 -385
rect 796 -428 838 -419
rect 872 -385 914 -376
rect 872 -419 879 -385
rect 909 -419 914 -385
rect 872 -424 914 -419
rect 948 -412 976 -352
tri 1021 -365 1043 -343 se
rect 1043 -350 1058 -342
tri 1043 -365 1058 -350 nw
tri 1015 -371 1021 -365 se
rect 1021 -371 1030 -365
rect 734 -456 762 -446
tri 762 -456 786 -432 sw
rect 734 -488 776 -456
tri 793 -464 794 -463 sw
rect 793 -488 794 -464
tri 796 -465 833 -428 ne
rect 833 -456 838 -428
tri 838 -456 864 -430 sw
rect 948 -446 957 -412
rect 948 -456 976 -446
rect 833 -465 917 -456
tri 833 -484 852 -465 ne
rect 852 -484 917 -465
rect 734 -510 794 -488
rect 916 -488 917 -484
rect 934 -488 976 -456
rect 916 -510 976 -488
rect 822 -526 839 -512
rect 871 -526 888 -512
tri 659 -562 681 -540 se
rect 681 -547 696 -526
tri 681 -562 696 -547 nw
rect 1015 -547 1030 -371
tri 1030 -378 1043 -365 nw
rect 1116 -446 1131 -218
tri 653 -568 659 -562 se
rect 659 -568 668 -562
rect 653 -584 668 -568
tri 668 -575 681 -562 nw
rect 822 -570 839 -556
rect 871 -570 888 -556
tri 1015 -562 1030 -547 ne
tri 1030 -562 1052 -540 sw
rect 653 -620 668 -612
rect 734 -584 794 -570
rect 749 -594 794 -584
rect 749 -612 777 -594
tri 653 -635 668 -620 ne
tri 668 -635 690 -613 sw
rect 734 -622 777 -612
rect 792 -598 794 -594
rect 916 -584 976 -570
tri 1030 -575 1043 -562 ne
rect 1043 -568 1052 -562
tri 1052 -568 1058 -562 sw
rect 916 -594 961 -584
rect 792 -622 866 -598
rect 734 -626 866 -622
tri 866 -626 894 -598 sw
rect 916 -608 918 -594
tri 916 -610 918 -608 ne
rect 930 -612 961 -594
rect 930 -622 976 -612
rect 1043 -583 1058 -568
tri 668 -647 680 -635 ne
rect 680 -640 690 -635
tri 690 -640 695 -635 sw
rect 579 -986 594 -758
rect 680 -796 695 -640
rect 734 -682 762 -626
tri 854 -644 872 -626 ne
rect 872 -646 894 -626
tri 894 -646 914 -626 sw
tri 930 -640 948 -622 ne
rect 753 -716 762 -682
rect 796 -655 838 -654
rect 796 -689 801 -655
rect 831 -689 838 -655
rect 796 -698 838 -689
rect 872 -655 914 -646
rect 872 -689 879 -655
rect 909 -689 914 -655
rect 872 -694 914 -689
rect 948 -682 976 -622
tri 1021 -635 1043 -613 se
rect 1043 -620 1058 -612
tri 1043 -635 1058 -620 nw
tri 1015 -641 1021 -635 se
rect 1021 -641 1030 -635
rect 734 -726 762 -716
tri 762 -726 786 -702 sw
rect 734 -758 776 -726
tri 793 -734 794 -733 sw
rect 793 -758 794 -734
tri 796 -735 833 -698 ne
rect 833 -726 838 -698
tri 838 -726 864 -700 sw
rect 948 -716 957 -682
rect 948 -726 976 -716
rect 833 -735 917 -726
tri 833 -754 852 -735 ne
rect 852 -754 917 -735
rect 734 -780 794 -758
rect 916 -758 917 -754
rect 934 -758 976 -726
rect 916 -780 976 -758
rect 822 -796 839 -782
rect 871 -796 888 -782
tri 659 -832 681 -810 se
rect 681 -817 696 -796
tri 681 -832 696 -817 nw
rect 1015 -817 1030 -641
tri 1030 -648 1043 -635 nw
rect 1116 -716 1131 -488
tri 653 -838 659 -832 se
rect 659 -838 668 -832
rect 653 -854 668 -838
tri 668 -845 681 -832 nw
rect 822 -840 839 -826
rect 871 -840 888 -826
tri 1015 -832 1030 -817 ne
tri 1030 -832 1052 -810 sw
rect 653 -890 668 -882
rect 734 -854 794 -840
rect 749 -864 794 -854
rect 749 -882 777 -864
tri 653 -905 668 -890 ne
tri 668 -905 690 -883 sw
rect 734 -892 777 -882
rect 792 -868 794 -864
rect 916 -854 976 -840
tri 1030 -845 1043 -832 ne
rect 1043 -838 1052 -832
tri 1052 -838 1058 -832 sw
rect 916 -864 961 -854
rect 792 -892 866 -868
rect 734 -896 866 -892
tri 866 -896 894 -868 sw
rect 916 -878 918 -864
tri 916 -880 918 -878 ne
rect 930 -882 961 -864
rect 930 -892 976 -882
rect 1043 -853 1058 -838
tri 668 -917 680 -905 ne
rect 680 -910 690 -905
tri 690 -910 695 -905 sw
rect 579 -1256 594 -1028
rect 680 -1066 695 -910
rect 734 -952 762 -896
tri 854 -914 872 -896 ne
rect 872 -916 894 -896
tri 894 -916 914 -896 sw
tri 930 -910 948 -892 ne
rect 753 -986 762 -952
rect 796 -925 838 -924
rect 796 -959 801 -925
rect 831 -959 838 -925
rect 796 -968 838 -959
rect 872 -925 914 -916
rect 872 -959 879 -925
rect 909 -959 914 -925
rect 872 -964 914 -959
rect 948 -952 976 -892
tri 1021 -905 1043 -883 se
rect 1043 -890 1058 -882
tri 1043 -905 1058 -890 nw
tri 1015 -911 1021 -905 se
rect 1021 -911 1030 -905
rect 734 -996 762 -986
tri 762 -996 786 -972 sw
rect 734 -1028 776 -996
tri 793 -1004 794 -1003 sw
rect 793 -1028 794 -1004
tri 796 -1005 833 -968 ne
rect 833 -996 838 -968
tri 838 -996 864 -970 sw
rect 948 -986 957 -952
rect 948 -996 976 -986
rect 833 -1005 917 -996
tri 833 -1024 852 -1005 ne
rect 852 -1024 917 -1005
rect 734 -1050 794 -1028
rect 916 -1028 917 -1024
rect 934 -1028 976 -996
rect 916 -1050 976 -1028
rect 822 -1066 839 -1052
rect 871 -1066 888 -1052
tri 659 -1102 681 -1080 se
rect 681 -1087 696 -1066
tri 681 -1102 696 -1087 nw
rect 1015 -1087 1030 -911
tri 1030 -918 1043 -905 nw
rect 1116 -986 1131 -758
tri 653 -1108 659 -1102 se
rect 659 -1108 668 -1102
rect 653 -1124 668 -1108
tri 668 -1115 681 -1102 nw
rect 822 -1110 839 -1096
rect 871 -1110 888 -1096
tri 1015 -1102 1030 -1087 ne
tri 1030 -1102 1052 -1080 sw
rect 653 -1160 668 -1152
rect 734 -1124 794 -1110
rect 749 -1134 794 -1124
rect 749 -1152 777 -1134
tri 653 -1175 668 -1160 ne
tri 668 -1175 690 -1153 sw
rect 734 -1162 777 -1152
rect 792 -1138 794 -1134
rect 916 -1124 976 -1110
tri 1030 -1115 1043 -1102 ne
rect 1043 -1108 1052 -1102
tri 1052 -1108 1058 -1102 sw
rect 916 -1134 961 -1124
rect 792 -1162 866 -1138
rect 734 -1166 866 -1162
tri 866 -1166 894 -1138 sw
rect 916 -1148 918 -1134
tri 916 -1150 918 -1148 ne
rect 930 -1152 961 -1134
rect 930 -1162 976 -1152
rect 1043 -1123 1058 -1108
tri 668 -1187 680 -1175 ne
rect 680 -1180 690 -1175
tri 690 -1180 695 -1175 sw
rect 579 -1526 594 -1298
rect 680 -1336 695 -1180
rect 734 -1222 762 -1166
tri 854 -1184 872 -1166 ne
rect 872 -1186 894 -1166
tri 894 -1186 914 -1166 sw
tri 930 -1180 948 -1162 ne
rect 753 -1256 762 -1222
rect 796 -1195 838 -1194
rect 796 -1229 801 -1195
rect 831 -1229 838 -1195
rect 796 -1238 838 -1229
rect 872 -1195 914 -1186
rect 872 -1229 879 -1195
rect 909 -1229 914 -1195
rect 872 -1234 914 -1229
rect 948 -1222 976 -1162
tri 1021 -1175 1043 -1153 se
rect 1043 -1160 1058 -1152
tri 1043 -1175 1058 -1160 nw
tri 1015 -1181 1021 -1175 se
rect 1021 -1181 1030 -1175
rect 734 -1266 762 -1256
tri 762 -1266 786 -1242 sw
rect 734 -1298 776 -1266
tri 793 -1274 794 -1273 sw
rect 793 -1298 794 -1274
tri 796 -1275 833 -1238 ne
rect 833 -1266 838 -1238
tri 838 -1266 864 -1240 sw
rect 948 -1256 957 -1222
rect 948 -1266 976 -1256
rect 833 -1275 917 -1266
tri 833 -1294 852 -1275 ne
rect 852 -1294 917 -1275
rect 734 -1320 794 -1298
rect 916 -1298 917 -1294
rect 934 -1298 976 -1266
rect 916 -1320 976 -1298
rect 822 -1336 839 -1322
rect 871 -1336 888 -1322
tri 659 -1372 681 -1350 se
rect 681 -1357 696 -1336
tri 681 -1372 696 -1357 nw
rect 1015 -1357 1030 -1181
tri 1030 -1188 1043 -1175 nw
rect 1116 -1256 1131 -1028
tri 653 -1378 659 -1372 se
rect 659 -1378 668 -1372
rect 653 -1394 668 -1378
tri 668 -1385 681 -1372 nw
rect 822 -1380 839 -1366
rect 871 -1380 888 -1366
tri 1015 -1372 1030 -1357 ne
tri 1030 -1372 1052 -1350 sw
rect 653 -1430 668 -1422
rect 734 -1394 794 -1380
rect 749 -1404 794 -1394
rect 749 -1422 777 -1404
tri 653 -1445 668 -1430 ne
tri 668 -1445 690 -1423 sw
rect 734 -1432 777 -1422
rect 792 -1408 794 -1404
rect 916 -1394 976 -1380
tri 1030 -1385 1043 -1372 ne
rect 1043 -1378 1052 -1372
tri 1052 -1378 1058 -1372 sw
rect 916 -1404 961 -1394
rect 792 -1432 866 -1408
rect 734 -1436 866 -1432
tri 866 -1436 894 -1408 sw
rect 916 -1418 918 -1404
tri 916 -1420 918 -1418 ne
rect 930 -1422 961 -1404
rect 930 -1432 976 -1422
rect 1043 -1393 1058 -1378
tri 668 -1457 680 -1445 ne
rect 680 -1450 690 -1445
tri 690 -1450 695 -1445 sw
rect 579 -1796 594 -1568
rect 680 -1606 695 -1450
rect 734 -1492 762 -1436
tri 854 -1454 872 -1436 ne
rect 872 -1456 894 -1436
tri 894 -1456 914 -1436 sw
tri 930 -1450 948 -1432 ne
rect 753 -1526 762 -1492
rect 796 -1465 838 -1464
rect 796 -1499 801 -1465
rect 831 -1499 838 -1465
rect 796 -1508 838 -1499
rect 872 -1465 914 -1456
rect 872 -1499 879 -1465
rect 909 -1499 914 -1465
rect 872 -1504 914 -1499
rect 948 -1492 976 -1432
tri 1021 -1445 1043 -1423 se
rect 1043 -1430 1058 -1422
tri 1043 -1445 1058 -1430 nw
tri 1015 -1451 1021 -1445 se
rect 1021 -1451 1030 -1445
rect 734 -1536 762 -1526
tri 762 -1536 786 -1512 sw
rect 734 -1568 776 -1536
tri 793 -1544 794 -1543 sw
rect 793 -1568 794 -1544
tri 796 -1545 833 -1508 ne
rect 833 -1536 838 -1508
tri 838 -1536 864 -1510 sw
rect 948 -1526 957 -1492
rect 948 -1536 976 -1526
rect 833 -1545 917 -1536
tri 833 -1564 852 -1545 ne
rect 852 -1564 917 -1545
rect 734 -1590 794 -1568
rect 916 -1568 917 -1564
rect 934 -1568 976 -1536
rect 916 -1590 976 -1568
rect 822 -1606 839 -1592
rect 871 -1606 888 -1592
tri 659 -1642 681 -1620 se
rect 681 -1627 696 -1606
tri 681 -1642 696 -1627 nw
rect 1015 -1627 1030 -1451
tri 1030 -1458 1043 -1445 nw
rect 1116 -1526 1131 -1298
tri 653 -1648 659 -1642 se
rect 659 -1648 668 -1642
rect 653 -1664 668 -1648
tri 668 -1655 681 -1642 nw
rect 822 -1650 839 -1636
rect 871 -1650 888 -1636
tri 1015 -1642 1030 -1627 ne
tri 1030 -1642 1052 -1620 sw
rect 653 -1700 668 -1692
rect 734 -1664 794 -1650
rect 749 -1674 794 -1664
rect 749 -1692 777 -1674
tri 653 -1715 668 -1700 ne
tri 668 -1715 690 -1693 sw
rect 734 -1702 777 -1692
rect 792 -1678 794 -1674
rect 916 -1664 976 -1650
tri 1030 -1655 1043 -1642 ne
rect 1043 -1648 1052 -1642
tri 1052 -1648 1058 -1642 sw
rect 916 -1674 961 -1664
rect 792 -1702 866 -1678
rect 734 -1706 866 -1702
tri 866 -1706 894 -1678 sw
rect 916 -1688 918 -1674
tri 916 -1690 918 -1688 ne
rect 930 -1692 961 -1674
rect 930 -1702 976 -1692
rect 1043 -1663 1058 -1648
tri 668 -1727 680 -1715 ne
rect 680 -1720 690 -1715
tri 690 -1720 695 -1715 sw
rect 579 -2066 594 -1838
rect 680 -1876 695 -1720
rect 734 -1762 762 -1706
tri 854 -1724 872 -1706 ne
rect 872 -1726 894 -1706
tri 894 -1726 914 -1706 sw
tri 930 -1720 948 -1702 ne
rect 753 -1796 762 -1762
rect 796 -1735 838 -1734
rect 796 -1769 801 -1735
rect 831 -1769 838 -1735
rect 796 -1778 838 -1769
rect 872 -1735 914 -1726
rect 872 -1769 879 -1735
rect 909 -1769 914 -1735
rect 872 -1774 914 -1769
rect 948 -1762 976 -1702
tri 1021 -1715 1043 -1693 se
rect 1043 -1700 1058 -1692
tri 1043 -1715 1058 -1700 nw
tri 1015 -1721 1021 -1715 se
rect 1021 -1721 1030 -1715
rect 734 -1806 762 -1796
tri 762 -1806 786 -1782 sw
rect 734 -1838 776 -1806
tri 793 -1814 794 -1813 sw
rect 793 -1838 794 -1814
tri 796 -1815 833 -1778 ne
rect 833 -1806 838 -1778
tri 838 -1806 864 -1780 sw
rect 948 -1796 957 -1762
rect 948 -1806 976 -1796
rect 833 -1815 917 -1806
tri 833 -1834 852 -1815 ne
rect 852 -1834 917 -1815
rect 734 -1860 794 -1838
rect 916 -1838 917 -1834
rect 934 -1838 976 -1806
rect 916 -1860 976 -1838
rect 822 -1876 839 -1862
rect 871 -1876 888 -1862
tri 659 -1912 681 -1890 se
rect 681 -1897 696 -1876
tri 681 -1912 696 -1897 nw
rect 1015 -1897 1030 -1721
tri 1030 -1728 1043 -1715 nw
rect 1116 -1796 1131 -1568
tri 653 -1918 659 -1912 se
rect 659 -1918 668 -1912
rect 653 -1934 668 -1918
tri 668 -1925 681 -1912 nw
rect 822 -1920 839 -1906
rect 871 -1920 888 -1906
tri 1015 -1912 1030 -1897 ne
tri 1030 -1912 1052 -1890 sw
rect 653 -1970 668 -1962
rect 734 -1934 794 -1920
rect 749 -1944 794 -1934
rect 749 -1962 777 -1944
tri 653 -1985 668 -1970 ne
tri 668 -1985 690 -1963 sw
rect 734 -1972 777 -1962
rect 792 -1948 794 -1944
rect 916 -1934 976 -1920
tri 1030 -1925 1043 -1912 ne
rect 1043 -1918 1052 -1912
tri 1052 -1918 1058 -1912 sw
rect 916 -1944 961 -1934
rect 792 -1972 866 -1948
rect 734 -1976 866 -1972
tri 866 -1976 894 -1948 sw
rect 916 -1958 918 -1944
tri 916 -1960 918 -1958 ne
rect 930 -1962 961 -1944
rect 930 -1972 976 -1962
rect 1043 -1933 1058 -1918
tri 668 -1997 680 -1985 ne
rect 680 -1990 690 -1985
tri 690 -1990 695 -1985 sw
rect 579 -2146 594 -2108
rect 680 -2146 695 -1990
rect 734 -2032 762 -1976
tri 854 -1994 872 -1976 ne
rect 872 -1996 894 -1976
tri 894 -1996 914 -1976 sw
tri 930 -1990 948 -1972 ne
rect 753 -2066 762 -2032
rect 796 -2005 838 -2004
rect 796 -2039 801 -2005
rect 831 -2039 838 -2005
rect 796 -2048 838 -2039
rect 872 -2005 914 -1996
rect 872 -2039 879 -2005
rect 909 -2039 914 -2005
rect 872 -2044 914 -2039
rect 948 -2032 976 -1972
tri 1021 -1985 1043 -1963 se
rect 1043 -1970 1058 -1962
tri 1043 -1985 1058 -1970 nw
tri 1015 -1991 1021 -1985 se
rect 1021 -1991 1030 -1985
rect 734 -2076 762 -2066
tri 762 -2076 786 -2052 sw
rect 734 -2108 776 -2076
tri 793 -2084 794 -2083 sw
rect 793 -2108 794 -2084
tri 796 -2085 833 -2048 ne
rect 833 -2076 838 -2048
tri 838 -2076 864 -2050 sw
rect 948 -2066 957 -2032
rect 948 -2076 976 -2066
rect 833 -2085 917 -2076
tri 833 -2104 852 -2085 ne
rect 852 -2104 917 -2085
rect 734 -2130 794 -2108
rect 916 -2108 917 -2104
rect 934 -2108 976 -2076
rect 916 -2130 976 -2108
rect 822 -2146 839 -2132
rect 871 -2146 888 -2132
rect 1015 -2146 1030 -1991
tri 1030 -1998 1043 -1985 nw
rect 1116 -2066 1131 -1838
rect 1116 -2146 1131 -2108
rect 1159 1984 1174 2174
tri 1239 2138 1261 2160 se
rect 1261 2153 1276 2174
tri 1261 2138 1276 2153 nw
rect 1595 2153 1610 2174
tri 1233 2132 1239 2138 se
rect 1239 2132 1248 2138
rect 1233 2116 1248 2132
tri 1248 2125 1261 2138 nw
rect 1402 2130 1419 2144
rect 1451 2130 1468 2144
tri 1595 2138 1610 2153 ne
tri 1610 2138 1632 2160 sw
rect 1233 2080 1248 2088
rect 1314 2116 1374 2130
rect 1329 2106 1374 2116
rect 1329 2088 1357 2106
tri 1233 2065 1248 2080 ne
tri 1248 2065 1270 2087 sw
rect 1314 2078 1357 2088
rect 1372 2102 1374 2106
rect 1496 2116 1556 2130
tri 1610 2125 1623 2138 ne
rect 1623 2132 1632 2138
tri 1632 2132 1638 2138 sw
rect 1496 2106 1541 2116
rect 1372 2078 1446 2102
rect 1314 2074 1446 2078
tri 1446 2074 1474 2102 sw
rect 1496 2092 1498 2106
tri 1496 2090 1498 2092 ne
rect 1510 2088 1541 2106
rect 1510 2078 1556 2088
rect 1623 2117 1638 2132
tri 1248 2053 1260 2065 ne
rect 1260 2060 1270 2065
tri 1270 2060 1275 2065 sw
rect 1159 1714 1174 1942
rect 1260 1904 1275 2060
rect 1314 2018 1342 2074
tri 1434 2056 1452 2074 ne
rect 1452 2054 1474 2074
tri 1474 2054 1494 2074 sw
tri 1510 2060 1528 2078 ne
rect 1333 1984 1342 2018
rect 1376 2045 1418 2046
rect 1376 2011 1381 2045
rect 1411 2011 1418 2045
rect 1376 2002 1418 2011
rect 1452 2045 1494 2054
rect 1452 2011 1459 2045
rect 1489 2011 1494 2045
rect 1452 2006 1494 2011
rect 1528 2018 1556 2078
tri 1601 2065 1623 2087 se
rect 1623 2080 1638 2088
tri 1623 2065 1638 2080 nw
tri 1595 2059 1601 2065 se
rect 1601 2059 1610 2065
rect 1314 1974 1342 1984
tri 1342 1974 1366 1998 sw
rect 1314 1942 1356 1974
tri 1373 1966 1374 1967 sw
rect 1373 1942 1374 1966
tri 1376 1965 1413 2002 ne
rect 1413 1974 1418 2002
tri 1418 1974 1444 2000 sw
rect 1528 1984 1537 2018
rect 1528 1974 1556 1984
rect 1413 1965 1497 1974
tri 1413 1946 1432 1965 ne
rect 1432 1946 1497 1965
rect 1314 1920 1374 1942
rect 1496 1942 1497 1946
rect 1514 1942 1556 1974
rect 1496 1920 1556 1942
rect 1402 1904 1419 1918
rect 1451 1904 1468 1918
tri 1239 1868 1261 1890 se
rect 1261 1883 1276 1904
tri 1261 1868 1276 1883 nw
rect 1595 1883 1610 2059
tri 1610 2052 1623 2065 nw
rect 1696 1984 1711 2174
tri 1233 1862 1239 1868 se
rect 1239 1862 1248 1868
rect 1233 1846 1248 1862
tri 1248 1855 1261 1868 nw
rect 1402 1860 1419 1874
rect 1451 1860 1468 1874
tri 1595 1868 1610 1883 ne
tri 1610 1868 1632 1890 sw
rect 1233 1810 1248 1818
rect 1314 1846 1374 1860
rect 1329 1836 1374 1846
rect 1329 1818 1357 1836
tri 1233 1795 1248 1810 ne
tri 1248 1795 1270 1817 sw
rect 1314 1808 1357 1818
rect 1372 1832 1374 1836
rect 1496 1846 1556 1860
tri 1610 1855 1623 1868 ne
rect 1623 1862 1632 1868
tri 1632 1862 1638 1868 sw
rect 1496 1836 1541 1846
rect 1372 1808 1446 1832
rect 1314 1804 1446 1808
tri 1446 1804 1474 1832 sw
rect 1496 1822 1498 1836
tri 1496 1820 1498 1822 ne
rect 1510 1818 1541 1836
rect 1510 1808 1556 1818
rect 1623 1847 1638 1862
tri 1248 1783 1260 1795 ne
rect 1260 1790 1270 1795
tri 1270 1790 1275 1795 sw
rect 1159 1444 1174 1672
rect 1260 1634 1275 1790
rect 1314 1748 1342 1804
tri 1434 1786 1452 1804 ne
rect 1452 1784 1474 1804
tri 1474 1784 1494 1804 sw
tri 1510 1790 1528 1808 ne
rect 1333 1714 1342 1748
rect 1376 1775 1418 1776
rect 1376 1741 1381 1775
rect 1411 1741 1418 1775
rect 1376 1732 1418 1741
rect 1452 1775 1494 1784
rect 1452 1741 1459 1775
rect 1489 1741 1494 1775
rect 1452 1736 1494 1741
rect 1528 1748 1556 1808
tri 1601 1795 1623 1817 se
rect 1623 1810 1638 1818
tri 1623 1795 1638 1810 nw
tri 1595 1789 1601 1795 se
rect 1601 1789 1610 1795
rect 1314 1704 1342 1714
tri 1342 1704 1366 1728 sw
rect 1314 1672 1356 1704
tri 1373 1696 1374 1697 sw
rect 1373 1672 1374 1696
tri 1376 1695 1413 1732 ne
rect 1413 1704 1418 1732
tri 1418 1704 1444 1730 sw
rect 1528 1714 1537 1748
rect 1528 1704 1556 1714
rect 1413 1695 1497 1704
tri 1413 1676 1432 1695 ne
rect 1432 1676 1497 1695
rect 1314 1650 1374 1672
rect 1496 1672 1497 1676
rect 1514 1672 1556 1704
rect 1496 1650 1556 1672
rect 1402 1634 1419 1648
rect 1451 1634 1468 1648
tri 1239 1598 1261 1620 se
rect 1261 1613 1276 1634
tri 1261 1598 1276 1613 nw
rect 1595 1613 1610 1789
tri 1610 1782 1623 1795 nw
rect 1696 1714 1711 1942
tri 1233 1592 1239 1598 se
rect 1239 1592 1248 1598
rect 1233 1576 1248 1592
tri 1248 1585 1261 1598 nw
rect 1402 1590 1419 1604
rect 1451 1590 1468 1604
tri 1595 1598 1610 1613 ne
tri 1610 1598 1632 1620 sw
rect 1233 1540 1248 1548
rect 1314 1576 1374 1590
rect 1329 1566 1374 1576
rect 1329 1548 1357 1566
tri 1233 1525 1248 1540 ne
tri 1248 1525 1270 1547 sw
rect 1314 1538 1357 1548
rect 1372 1562 1374 1566
rect 1496 1576 1556 1590
tri 1610 1585 1623 1598 ne
rect 1623 1592 1632 1598
tri 1632 1592 1638 1598 sw
rect 1496 1566 1541 1576
rect 1372 1538 1446 1562
rect 1314 1534 1446 1538
tri 1446 1534 1474 1562 sw
rect 1496 1552 1498 1566
tri 1496 1550 1498 1552 ne
rect 1510 1548 1541 1566
rect 1510 1538 1556 1548
rect 1623 1577 1638 1592
tri 1248 1513 1260 1525 ne
rect 1260 1520 1270 1525
tri 1270 1520 1275 1525 sw
rect 1159 1174 1174 1402
rect 1260 1364 1275 1520
rect 1314 1478 1342 1534
tri 1434 1516 1452 1534 ne
rect 1452 1514 1474 1534
tri 1474 1514 1494 1534 sw
tri 1510 1520 1528 1538 ne
rect 1333 1444 1342 1478
rect 1376 1505 1418 1506
rect 1376 1471 1381 1505
rect 1411 1471 1418 1505
rect 1376 1462 1418 1471
rect 1452 1505 1494 1514
rect 1452 1471 1459 1505
rect 1489 1471 1494 1505
rect 1452 1466 1494 1471
rect 1528 1478 1556 1538
tri 1601 1525 1623 1547 se
rect 1623 1540 1638 1548
tri 1623 1525 1638 1540 nw
tri 1595 1519 1601 1525 se
rect 1601 1519 1610 1525
rect 1314 1434 1342 1444
tri 1342 1434 1366 1458 sw
rect 1314 1402 1356 1434
tri 1373 1426 1374 1427 sw
rect 1373 1402 1374 1426
tri 1376 1425 1413 1462 ne
rect 1413 1434 1418 1462
tri 1418 1434 1444 1460 sw
rect 1528 1444 1537 1478
rect 1528 1434 1556 1444
rect 1413 1425 1497 1434
tri 1413 1406 1432 1425 ne
rect 1432 1406 1497 1425
rect 1314 1380 1374 1402
rect 1496 1402 1497 1406
rect 1514 1402 1556 1434
rect 1496 1380 1556 1402
rect 1402 1364 1419 1378
rect 1451 1364 1468 1378
tri 1239 1328 1261 1350 se
rect 1261 1343 1276 1364
tri 1261 1328 1276 1343 nw
rect 1595 1343 1610 1519
tri 1610 1512 1623 1525 nw
rect 1696 1444 1711 1672
tri 1233 1322 1239 1328 se
rect 1239 1322 1248 1328
rect 1233 1306 1248 1322
tri 1248 1315 1261 1328 nw
rect 1402 1320 1419 1334
rect 1451 1320 1468 1334
tri 1595 1328 1610 1343 ne
tri 1610 1328 1632 1350 sw
rect 1233 1270 1248 1278
rect 1314 1306 1374 1320
rect 1329 1296 1374 1306
rect 1329 1278 1357 1296
tri 1233 1255 1248 1270 ne
tri 1248 1255 1270 1277 sw
rect 1314 1268 1357 1278
rect 1372 1292 1374 1296
rect 1496 1306 1556 1320
tri 1610 1315 1623 1328 ne
rect 1623 1322 1632 1328
tri 1632 1322 1638 1328 sw
rect 1496 1296 1541 1306
rect 1372 1268 1446 1292
rect 1314 1264 1446 1268
tri 1446 1264 1474 1292 sw
rect 1496 1282 1498 1296
tri 1496 1280 1498 1282 ne
rect 1510 1278 1541 1296
rect 1510 1268 1556 1278
rect 1623 1307 1638 1322
tri 1248 1243 1260 1255 ne
rect 1260 1250 1270 1255
tri 1270 1250 1275 1255 sw
rect 1159 904 1174 1132
rect 1260 1094 1275 1250
rect 1314 1208 1342 1264
tri 1434 1246 1452 1264 ne
rect 1452 1244 1474 1264
tri 1474 1244 1494 1264 sw
tri 1510 1250 1528 1268 ne
rect 1333 1174 1342 1208
rect 1376 1235 1418 1236
rect 1376 1201 1381 1235
rect 1411 1201 1418 1235
rect 1376 1192 1418 1201
rect 1452 1235 1494 1244
rect 1452 1201 1459 1235
rect 1489 1201 1494 1235
rect 1452 1196 1494 1201
rect 1528 1208 1556 1268
tri 1601 1255 1623 1277 se
rect 1623 1270 1638 1278
tri 1623 1255 1638 1270 nw
tri 1595 1249 1601 1255 se
rect 1601 1249 1610 1255
rect 1314 1164 1342 1174
tri 1342 1164 1366 1188 sw
rect 1314 1132 1356 1164
tri 1373 1156 1374 1157 sw
rect 1373 1132 1374 1156
tri 1376 1155 1413 1192 ne
rect 1413 1164 1418 1192
tri 1418 1164 1444 1190 sw
rect 1528 1174 1537 1208
rect 1528 1164 1556 1174
rect 1413 1155 1497 1164
tri 1413 1136 1432 1155 ne
rect 1432 1136 1497 1155
rect 1314 1110 1374 1132
rect 1496 1132 1497 1136
rect 1514 1132 1556 1164
rect 1496 1110 1556 1132
rect 1402 1094 1419 1108
rect 1451 1094 1468 1108
tri 1239 1058 1261 1080 se
rect 1261 1073 1276 1094
tri 1261 1058 1276 1073 nw
rect 1595 1073 1610 1249
tri 1610 1242 1623 1255 nw
rect 1696 1174 1711 1402
tri 1233 1052 1239 1058 se
rect 1239 1052 1248 1058
rect 1233 1036 1248 1052
tri 1248 1045 1261 1058 nw
rect 1402 1050 1419 1064
rect 1451 1050 1468 1064
tri 1595 1058 1610 1073 ne
tri 1610 1058 1632 1080 sw
rect 1233 1000 1248 1008
rect 1314 1036 1374 1050
rect 1329 1026 1374 1036
rect 1329 1008 1357 1026
tri 1233 985 1248 1000 ne
tri 1248 985 1270 1007 sw
rect 1314 998 1357 1008
rect 1372 1022 1374 1026
rect 1496 1036 1556 1050
tri 1610 1045 1623 1058 ne
rect 1623 1052 1632 1058
tri 1632 1052 1638 1058 sw
rect 1496 1026 1541 1036
rect 1372 998 1446 1022
rect 1314 994 1446 998
tri 1446 994 1474 1022 sw
rect 1496 1012 1498 1026
tri 1496 1010 1498 1012 ne
rect 1510 1008 1541 1026
rect 1510 998 1556 1008
rect 1623 1037 1638 1052
tri 1248 973 1260 985 ne
rect 1260 980 1270 985
tri 1270 980 1275 985 sw
rect 1159 634 1174 862
rect 1260 824 1275 980
rect 1314 938 1342 994
tri 1434 976 1452 994 ne
rect 1452 974 1474 994
tri 1474 974 1494 994 sw
tri 1510 980 1528 998 ne
rect 1333 904 1342 938
rect 1376 965 1418 966
rect 1376 931 1381 965
rect 1411 931 1418 965
rect 1376 922 1418 931
rect 1452 965 1494 974
rect 1452 931 1459 965
rect 1489 931 1494 965
rect 1452 926 1494 931
rect 1528 938 1556 998
tri 1601 985 1623 1007 se
rect 1623 1000 1638 1008
tri 1623 985 1638 1000 nw
tri 1595 979 1601 985 se
rect 1601 979 1610 985
rect 1314 894 1342 904
tri 1342 894 1366 918 sw
rect 1314 862 1356 894
tri 1373 886 1374 887 sw
rect 1373 862 1374 886
tri 1376 885 1413 922 ne
rect 1413 894 1418 922
tri 1418 894 1444 920 sw
rect 1528 904 1537 938
rect 1528 894 1556 904
rect 1413 885 1497 894
tri 1413 866 1432 885 ne
rect 1432 866 1497 885
rect 1314 840 1374 862
rect 1496 862 1497 866
rect 1514 862 1556 894
rect 1496 840 1556 862
rect 1402 824 1419 838
rect 1451 824 1468 838
tri 1239 788 1261 810 se
rect 1261 803 1276 824
tri 1261 788 1276 803 nw
rect 1595 803 1610 979
tri 1610 972 1623 985 nw
rect 1696 904 1711 1132
tri 1233 782 1239 788 se
rect 1239 782 1248 788
rect 1233 766 1248 782
tri 1248 775 1261 788 nw
rect 1402 780 1419 794
rect 1451 780 1468 794
tri 1595 788 1610 803 ne
tri 1610 788 1632 810 sw
rect 1233 730 1248 738
rect 1314 766 1374 780
rect 1329 756 1374 766
rect 1329 738 1357 756
tri 1233 715 1248 730 ne
tri 1248 715 1270 737 sw
rect 1314 728 1357 738
rect 1372 752 1374 756
rect 1496 766 1556 780
tri 1610 775 1623 788 ne
rect 1623 782 1632 788
tri 1632 782 1638 788 sw
rect 1496 756 1541 766
rect 1372 728 1446 752
rect 1314 724 1446 728
tri 1446 724 1474 752 sw
rect 1496 742 1498 756
tri 1496 740 1498 742 ne
rect 1510 738 1541 756
rect 1510 728 1556 738
rect 1623 767 1638 782
tri 1248 703 1260 715 ne
rect 1260 710 1270 715
tri 1270 710 1275 715 sw
rect 1159 364 1174 592
rect 1260 554 1275 710
rect 1314 668 1342 724
tri 1434 706 1452 724 ne
rect 1452 704 1474 724
tri 1474 704 1494 724 sw
tri 1510 710 1528 728 ne
rect 1333 634 1342 668
rect 1376 695 1418 696
rect 1376 661 1381 695
rect 1411 661 1418 695
rect 1376 652 1418 661
rect 1452 695 1494 704
rect 1452 661 1459 695
rect 1489 661 1494 695
rect 1452 656 1494 661
rect 1528 668 1556 728
tri 1601 715 1623 737 se
rect 1623 730 1638 738
tri 1623 715 1638 730 nw
tri 1595 709 1601 715 se
rect 1601 709 1610 715
rect 1314 624 1342 634
tri 1342 624 1366 648 sw
rect 1314 592 1356 624
tri 1373 616 1374 617 sw
rect 1373 592 1374 616
tri 1376 615 1413 652 ne
rect 1413 624 1418 652
tri 1418 624 1444 650 sw
rect 1528 634 1537 668
rect 1528 624 1556 634
rect 1413 615 1497 624
tri 1413 596 1432 615 ne
rect 1432 596 1497 615
rect 1314 570 1374 592
rect 1496 592 1497 596
rect 1514 592 1556 624
rect 1496 570 1556 592
rect 1402 554 1419 568
rect 1451 554 1468 568
tri 1239 518 1261 540 se
rect 1261 533 1276 554
tri 1261 518 1276 533 nw
rect 1595 533 1610 709
tri 1610 702 1623 715 nw
rect 1696 634 1711 862
tri 1233 512 1239 518 se
rect 1239 512 1248 518
rect 1233 496 1248 512
tri 1248 505 1261 518 nw
rect 1402 510 1419 524
rect 1451 510 1468 524
tri 1595 518 1610 533 ne
tri 1610 518 1632 540 sw
rect 1233 460 1248 468
rect 1314 496 1374 510
rect 1329 486 1374 496
rect 1329 468 1357 486
tri 1233 445 1248 460 ne
tri 1248 445 1270 467 sw
rect 1314 458 1357 468
rect 1372 482 1374 486
rect 1496 496 1556 510
tri 1610 505 1623 518 ne
rect 1623 512 1632 518
tri 1632 512 1638 518 sw
rect 1496 486 1541 496
rect 1372 458 1446 482
rect 1314 454 1446 458
tri 1446 454 1474 482 sw
rect 1496 472 1498 486
tri 1496 470 1498 472 ne
rect 1510 468 1541 486
rect 1510 458 1556 468
rect 1623 497 1638 512
tri 1248 433 1260 445 ne
rect 1260 440 1270 445
tri 1270 440 1275 445 sw
rect 1159 94 1174 322
rect 1260 284 1275 440
rect 1314 398 1342 454
tri 1434 436 1452 454 ne
rect 1452 434 1474 454
tri 1474 434 1494 454 sw
tri 1510 440 1528 458 ne
rect 1333 364 1342 398
rect 1376 425 1418 426
rect 1376 391 1381 425
rect 1411 391 1418 425
rect 1376 382 1418 391
rect 1452 425 1494 434
rect 1452 391 1459 425
rect 1489 391 1494 425
rect 1452 386 1494 391
rect 1528 398 1556 458
tri 1601 445 1623 467 se
rect 1623 460 1638 468
tri 1623 445 1638 460 nw
tri 1595 439 1601 445 se
rect 1601 439 1610 445
rect 1314 354 1342 364
tri 1342 354 1366 378 sw
rect 1314 322 1356 354
tri 1373 346 1374 347 sw
rect 1373 322 1374 346
tri 1376 345 1413 382 ne
rect 1413 354 1418 382
tri 1418 354 1444 380 sw
rect 1528 364 1537 398
rect 1528 354 1556 364
rect 1413 345 1497 354
tri 1413 326 1432 345 ne
rect 1432 326 1497 345
rect 1314 300 1374 322
rect 1496 322 1497 326
rect 1514 322 1556 354
rect 1496 300 1556 322
rect 1402 284 1419 298
rect 1451 284 1468 298
tri 1239 248 1261 270 se
rect 1261 263 1276 284
tri 1261 248 1276 263 nw
rect 1595 263 1610 439
tri 1610 432 1623 445 nw
rect 1696 364 1711 592
tri 1233 242 1239 248 se
rect 1239 242 1248 248
rect 1233 226 1248 242
tri 1248 235 1261 248 nw
rect 1402 240 1419 254
rect 1451 240 1468 254
tri 1595 248 1610 263 ne
tri 1610 248 1632 270 sw
rect 1233 190 1248 198
rect 1314 226 1374 240
rect 1329 216 1374 226
rect 1329 198 1357 216
tri 1233 175 1248 190 ne
tri 1248 175 1270 197 sw
rect 1314 188 1357 198
rect 1372 212 1374 216
rect 1496 226 1556 240
tri 1610 235 1623 248 ne
rect 1623 242 1632 248
tri 1632 242 1638 248 sw
rect 1496 216 1541 226
rect 1372 188 1446 212
rect 1314 184 1446 188
tri 1446 184 1474 212 sw
rect 1496 202 1498 216
tri 1496 200 1498 202 ne
rect 1510 198 1541 216
rect 1510 188 1556 198
rect 1623 227 1638 242
tri 1248 163 1260 175 ne
rect 1260 170 1270 175
tri 1270 170 1275 175 sw
rect 1159 -176 1174 52
rect 1260 14 1275 170
rect 1314 128 1342 184
tri 1434 166 1452 184 ne
rect 1452 164 1474 184
tri 1474 164 1494 184 sw
tri 1510 170 1528 188 ne
rect 1333 94 1342 128
rect 1376 155 1418 156
rect 1376 121 1381 155
rect 1411 121 1418 155
rect 1376 112 1418 121
rect 1452 155 1494 164
rect 1452 121 1459 155
rect 1489 121 1494 155
rect 1452 116 1494 121
rect 1528 128 1556 188
tri 1601 175 1623 197 se
rect 1623 190 1638 198
tri 1623 175 1638 190 nw
tri 1595 169 1601 175 se
rect 1601 169 1610 175
rect 1314 84 1342 94
tri 1342 84 1366 108 sw
rect 1314 52 1356 84
tri 1373 76 1374 77 sw
rect 1373 52 1374 76
tri 1376 75 1413 112 ne
rect 1413 84 1418 112
tri 1418 84 1444 110 sw
rect 1528 94 1537 128
rect 1528 84 1556 94
rect 1413 75 1497 84
tri 1413 56 1432 75 ne
rect 1432 56 1497 75
rect 1314 30 1374 52
rect 1496 52 1497 56
rect 1514 52 1556 84
rect 1496 30 1556 52
rect 1402 14 1419 28
rect 1451 14 1468 28
tri 1239 -22 1261 0 se
rect 1261 -7 1276 14
tri 1261 -22 1276 -7 nw
rect 1595 -7 1610 169
tri 1610 162 1623 175 nw
rect 1696 94 1711 322
tri 1233 -28 1239 -22 se
rect 1239 -28 1248 -22
rect 1233 -44 1248 -28
tri 1248 -35 1261 -22 nw
rect 1402 -30 1419 -16
rect 1451 -30 1468 -16
tri 1595 -22 1610 -7 ne
tri 1610 -22 1632 0 sw
rect 1233 -80 1248 -72
rect 1314 -44 1374 -30
rect 1329 -54 1374 -44
rect 1329 -72 1357 -54
tri 1233 -95 1248 -80 ne
tri 1248 -95 1270 -73 sw
rect 1314 -82 1357 -72
rect 1372 -58 1374 -54
rect 1496 -44 1556 -30
tri 1610 -35 1623 -22 ne
rect 1623 -28 1632 -22
tri 1632 -28 1638 -22 sw
rect 1496 -54 1541 -44
rect 1372 -82 1446 -58
rect 1314 -86 1446 -82
tri 1446 -86 1474 -58 sw
rect 1496 -68 1498 -54
tri 1496 -70 1498 -68 ne
rect 1510 -72 1541 -54
rect 1510 -82 1556 -72
rect 1623 -43 1638 -28
tri 1248 -107 1260 -95 ne
rect 1260 -100 1270 -95
tri 1270 -100 1275 -95 sw
rect 1159 -446 1174 -218
rect 1260 -256 1275 -100
rect 1314 -142 1342 -86
tri 1434 -104 1452 -86 ne
rect 1452 -106 1474 -86
tri 1474 -106 1494 -86 sw
tri 1510 -100 1528 -82 ne
rect 1333 -176 1342 -142
rect 1376 -115 1418 -114
rect 1376 -149 1381 -115
rect 1411 -149 1418 -115
rect 1376 -158 1418 -149
rect 1452 -115 1494 -106
rect 1452 -149 1459 -115
rect 1489 -149 1494 -115
rect 1452 -154 1494 -149
rect 1528 -142 1556 -82
tri 1601 -95 1623 -73 se
rect 1623 -80 1638 -72
tri 1623 -95 1638 -80 nw
tri 1595 -101 1601 -95 se
rect 1601 -101 1610 -95
rect 1314 -186 1342 -176
tri 1342 -186 1366 -162 sw
rect 1314 -218 1356 -186
tri 1373 -194 1374 -193 sw
rect 1373 -218 1374 -194
tri 1376 -195 1413 -158 ne
rect 1413 -186 1418 -158
tri 1418 -186 1444 -160 sw
rect 1528 -176 1537 -142
rect 1528 -186 1556 -176
rect 1413 -195 1497 -186
tri 1413 -214 1432 -195 ne
rect 1432 -214 1497 -195
rect 1314 -240 1374 -218
rect 1496 -218 1497 -214
rect 1514 -218 1556 -186
rect 1496 -240 1556 -218
rect 1402 -256 1419 -242
rect 1451 -256 1468 -242
tri 1239 -292 1261 -270 se
rect 1261 -277 1276 -256
tri 1261 -292 1276 -277 nw
rect 1595 -277 1610 -101
tri 1610 -108 1623 -95 nw
rect 1696 -176 1711 52
tri 1233 -298 1239 -292 se
rect 1239 -298 1248 -292
rect 1233 -314 1248 -298
tri 1248 -305 1261 -292 nw
rect 1402 -300 1419 -286
rect 1451 -300 1468 -286
tri 1595 -292 1610 -277 ne
tri 1610 -292 1632 -270 sw
rect 1233 -350 1248 -342
rect 1314 -314 1374 -300
rect 1329 -324 1374 -314
rect 1329 -342 1357 -324
tri 1233 -365 1248 -350 ne
tri 1248 -365 1270 -343 sw
rect 1314 -352 1357 -342
rect 1372 -328 1374 -324
rect 1496 -314 1556 -300
tri 1610 -305 1623 -292 ne
rect 1623 -298 1632 -292
tri 1632 -298 1638 -292 sw
rect 1496 -324 1541 -314
rect 1372 -352 1446 -328
rect 1314 -356 1446 -352
tri 1446 -356 1474 -328 sw
rect 1496 -338 1498 -324
tri 1496 -340 1498 -338 ne
rect 1510 -342 1541 -324
rect 1510 -352 1556 -342
rect 1623 -313 1638 -298
tri 1248 -377 1260 -365 ne
rect 1260 -370 1270 -365
tri 1270 -370 1275 -365 sw
rect 1159 -716 1174 -488
rect 1260 -526 1275 -370
rect 1314 -412 1342 -356
tri 1434 -374 1452 -356 ne
rect 1452 -376 1474 -356
tri 1474 -376 1494 -356 sw
tri 1510 -370 1528 -352 ne
rect 1333 -446 1342 -412
rect 1376 -385 1418 -384
rect 1376 -419 1381 -385
rect 1411 -419 1418 -385
rect 1376 -428 1418 -419
rect 1452 -385 1494 -376
rect 1452 -419 1459 -385
rect 1489 -419 1494 -385
rect 1452 -424 1494 -419
rect 1528 -412 1556 -352
tri 1601 -365 1623 -343 se
rect 1623 -350 1638 -342
tri 1623 -365 1638 -350 nw
tri 1595 -371 1601 -365 se
rect 1601 -371 1610 -365
rect 1314 -456 1342 -446
tri 1342 -456 1366 -432 sw
rect 1314 -488 1356 -456
tri 1373 -464 1374 -463 sw
rect 1373 -488 1374 -464
tri 1376 -465 1413 -428 ne
rect 1413 -456 1418 -428
tri 1418 -456 1444 -430 sw
rect 1528 -446 1537 -412
rect 1528 -456 1556 -446
rect 1413 -465 1497 -456
tri 1413 -484 1432 -465 ne
rect 1432 -484 1497 -465
rect 1314 -510 1374 -488
rect 1496 -488 1497 -484
rect 1514 -488 1556 -456
rect 1496 -510 1556 -488
rect 1402 -526 1419 -512
rect 1451 -526 1468 -512
tri 1239 -562 1261 -540 se
rect 1261 -547 1276 -526
tri 1261 -562 1276 -547 nw
rect 1595 -547 1610 -371
tri 1610 -378 1623 -365 nw
rect 1696 -446 1711 -218
tri 1233 -568 1239 -562 se
rect 1239 -568 1248 -562
rect 1233 -584 1248 -568
tri 1248 -575 1261 -562 nw
rect 1402 -570 1419 -556
rect 1451 -570 1468 -556
tri 1595 -562 1610 -547 ne
tri 1610 -562 1632 -540 sw
rect 1233 -620 1248 -612
rect 1314 -584 1374 -570
rect 1329 -594 1374 -584
rect 1329 -612 1357 -594
tri 1233 -635 1248 -620 ne
tri 1248 -635 1270 -613 sw
rect 1314 -622 1357 -612
rect 1372 -598 1374 -594
rect 1496 -584 1556 -570
tri 1610 -575 1623 -562 ne
rect 1623 -568 1632 -562
tri 1632 -568 1638 -562 sw
rect 1496 -594 1541 -584
rect 1372 -622 1446 -598
rect 1314 -626 1446 -622
tri 1446 -626 1474 -598 sw
rect 1496 -608 1498 -594
tri 1496 -610 1498 -608 ne
rect 1510 -612 1541 -594
rect 1510 -622 1556 -612
rect 1623 -583 1638 -568
tri 1248 -647 1260 -635 ne
rect 1260 -640 1270 -635
tri 1270 -640 1275 -635 sw
rect 1159 -986 1174 -758
rect 1260 -796 1275 -640
rect 1314 -682 1342 -626
tri 1434 -644 1452 -626 ne
rect 1452 -646 1474 -626
tri 1474 -646 1494 -626 sw
tri 1510 -640 1528 -622 ne
rect 1333 -716 1342 -682
rect 1376 -655 1418 -654
rect 1376 -689 1381 -655
rect 1411 -689 1418 -655
rect 1376 -698 1418 -689
rect 1452 -655 1494 -646
rect 1452 -689 1459 -655
rect 1489 -689 1494 -655
rect 1452 -694 1494 -689
rect 1528 -682 1556 -622
tri 1601 -635 1623 -613 se
rect 1623 -620 1638 -612
tri 1623 -635 1638 -620 nw
tri 1595 -641 1601 -635 se
rect 1601 -641 1610 -635
rect 1314 -726 1342 -716
tri 1342 -726 1366 -702 sw
rect 1314 -758 1356 -726
tri 1373 -734 1374 -733 sw
rect 1373 -758 1374 -734
tri 1376 -735 1413 -698 ne
rect 1413 -726 1418 -698
tri 1418 -726 1444 -700 sw
rect 1528 -716 1537 -682
rect 1528 -726 1556 -716
rect 1413 -735 1497 -726
tri 1413 -754 1432 -735 ne
rect 1432 -754 1497 -735
rect 1314 -780 1374 -758
rect 1496 -758 1497 -754
rect 1514 -758 1556 -726
rect 1496 -780 1556 -758
rect 1402 -796 1419 -782
rect 1451 -796 1468 -782
tri 1239 -832 1261 -810 se
rect 1261 -817 1276 -796
tri 1261 -832 1276 -817 nw
rect 1595 -817 1610 -641
tri 1610 -648 1623 -635 nw
rect 1696 -716 1711 -488
tri 1233 -838 1239 -832 se
rect 1239 -838 1248 -832
rect 1233 -854 1248 -838
tri 1248 -845 1261 -832 nw
rect 1402 -840 1419 -826
rect 1451 -840 1468 -826
tri 1595 -832 1610 -817 ne
tri 1610 -832 1632 -810 sw
rect 1233 -890 1248 -882
rect 1314 -854 1374 -840
rect 1329 -864 1374 -854
rect 1329 -882 1357 -864
tri 1233 -905 1248 -890 ne
tri 1248 -905 1270 -883 sw
rect 1314 -892 1357 -882
rect 1372 -868 1374 -864
rect 1496 -854 1556 -840
tri 1610 -845 1623 -832 ne
rect 1623 -838 1632 -832
tri 1632 -838 1638 -832 sw
rect 1496 -864 1541 -854
rect 1372 -892 1446 -868
rect 1314 -896 1446 -892
tri 1446 -896 1474 -868 sw
rect 1496 -878 1498 -864
tri 1496 -880 1498 -878 ne
rect 1510 -882 1541 -864
rect 1510 -892 1556 -882
rect 1623 -853 1638 -838
tri 1248 -917 1260 -905 ne
rect 1260 -910 1270 -905
tri 1270 -910 1275 -905 sw
rect 1159 -1256 1174 -1028
rect 1260 -1066 1275 -910
rect 1314 -952 1342 -896
tri 1434 -914 1452 -896 ne
rect 1452 -916 1474 -896
tri 1474 -916 1494 -896 sw
tri 1510 -910 1528 -892 ne
rect 1333 -986 1342 -952
rect 1376 -925 1418 -924
rect 1376 -959 1381 -925
rect 1411 -959 1418 -925
rect 1376 -968 1418 -959
rect 1452 -925 1494 -916
rect 1452 -959 1459 -925
rect 1489 -959 1494 -925
rect 1452 -964 1494 -959
rect 1528 -952 1556 -892
tri 1601 -905 1623 -883 se
rect 1623 -890 1638 -882
tri 1623 -905 1638 -890 nw
tri 1595 -911 1601 -905 se
rect 1601 -911 1610 -905
rect 1314 -996 1342 -986
tri 1342 -996 1366 -972 sw
rect 1314 -1028 1356 -996
tri 1373 -1004 1374 -1003 sw
rect 1373 -1028 1374 -1004
tri 1376 -1005 1413 -968 ne
rect 1413 -996 1418 -968
tri 1418 -996 1444 -970 sw
rect 1528 -986 1537 -952
rect 1528 -996 1556 -986
rect 1413 -1005 1497 -996
tri 1413 -1024 1432 -1005 ne
rect 1432 -1024 1497 -1005
rect 1314 -1050 1374 -1028
rect 1496 -1028 1497 -1024
rect 1514 -1028 1556 -996
rect 1496 -1050 1556 -1028
rect 1402 -1066 1419 -1052
rect 1451 -1066 1468 -1052
tri 1239 -1102 1261 -1080 se
rect 1261 -1087 1276 -1066
tri 1261 -1102 1276 -1087 nw
rect 1595 -1087 1610 -911
tri 1610 -918 1623 -905 nw
rect 1696 -986 1711 -758
tri 1233 -1108 1239 -1102 se
rect 1239 -1108 1248 -1102
rect 1233 -1124 1248 -1108
tri 1248 -1115 1261 -1102 nw
rect 1402 -1110 1419 -1096
rect 1451 -1110 1468 -1096
tri 1595 -1102 1610 -1087 ne
tri 1610 -1102 1632 -1080 sw
rect 1233 -1160 1248 -1152
rect 1314 -1124 1374 -1110
rect 1329 -1134 1374 -1124
rect 1329 -1152 1357 -1134
tri 1233 -1175 1248 -1160 ne
tri 1248 -1175 1270 -1153 sw
rect 1314 -1162 1357 -1152
rect 1372 -1138 1374 -1134
rect 1496 -1124 1556 -1110
tri 1610 -1115 1623 -1102 ne
rect 1623 -1108 1632 -1102
tri 1632 -1108 1638 -1102 sw
rect 1496 -1134 1541 -1124
rect 1372 -1162 1446 -1138
rect 1314 -1166 1446 -1162
tri 1446 -1166 1474 -1138 sw
rect 1496 -1148 1498 -1134
tri 1496 -1150 1498 -1148 ne
rect 1510 -1152 1541 -1134
rect 1510 -1162 1556 -1152
rect 1623 -1123 1638 -1108
tri 1248 -1187 1260 -1175 ne
rect 1260 -1180 1270 -1175
tri 1270 -1180 1275 -1175 sw
rect 1159 -1526 1174 -1298
rect 1260 -1336 1275 -1180
rect 1314 -1222 1342 -1166
tri 1434 -1184 1452 -1166 ne
rect 1452 -1186 1474 -1166
tri 1474 -1186 1494 -1166 sw
tri 1510 -1180 1528 -1162 ne
rect 1333 -1256 1342 -1222
rect 1376 -1195 1418 -1194
rect 1376 -1229 1381 -1195
rect 1411 -1229 1418 -1195
rect 1376 -1238 1418 -1229
rect 1452 -1195 1494 -1186
rect 1452 -1229 1459 -1195
rect 1489 -1229 1494 -1195
rect 1452 -1234 1494 -1229
rect 1528 -1222 1556 -1162
tri 1601 -1175 1623 -1153 se
rect 1623 -1160 1638 -1152
tri 1623 -1175 1638 -1160 nw
tri 1595 -1181 1601 -1175 se
rect 1601 -1181 1610 -1175
rect 1314 -1266 1342 -1256
tri 1342 -1266 1366 -1242 sw
rect 1314 -1298 1356 -1266
tri 1373 -1274 1374 -1273 sw
rect 1373 -1298 1374 -1274
tri 1376 -1275 1413 -1238 ne
rect 1413 -1266 1418 -1238
tri 1418 -1266 1444 -1240 sw
rect 1528 -1256 1537 -1222
rect 1528 -1266 1556 -1256
rect 1413 -1275 1497 -1266
tri 1413 -1294 1432 -1275 ne
rect 1432 -1294 1497 -1275
rect 1314 -1320 1374 -1298
rect 1496 -1298 1497 -1294
rect 1514 -1298 1556 -1266
rect 1496 -1320 1556 -1298
rect 1402 -1336 1419 -1322
rect 1451 -1336 1468 -1322
tri 1239 -1372 1261 -1350 se
rect 1261 -1357 1276 -1336
tri 1261 -1372 1276 -1357 nw
rect 1595 -1357 1610 -1181
tri 1610 -1188 1623 -1175 nw
rect 1696 -1256 1711 -1028
tri 1233 -1378 1239 -1372 se
rect 1239 -1378 1248 -1372
rect 1233 -1394 1248 -1378
tri 1248 -1385 1261 -1372 nw
rect 1402 -1380 1419 -1366
rect 1451 -1380 1468 -1366
tri 1595 -1372 1610 -1357 ne
tri 1610 -1372 1632 -1350 sw
rect 1233 -1430 1248 -1422
rect 1314 -1394 1374 -1380
rect 1329 -1404 1374 -1394
rect 1329 -1422 1357 -1404
tri 1233 -1445 1248 -1430 ne
tri 1248 -1445 1270 -1423 sw
rect 1314 -1432 1357 -1422
rect 1372 -1408 1374 -1404
rect 1496 -1394 1556 -1380
tri 1610 -1385 1623 -1372 ne
rect 1623 -1378 1632 -1372
tri 1632 -1378 1638 -1372 sw
rect 1496 -1404 1541 -1394
rect 1372 -1432 1446 -1408
rect 1314 -1436 1446 -1432
tri 1446 -1436 1474 -1408 sw
rect 1496 -1418 1498 -1404
tri 1496 -1420 1498 -1418 ne
rect 1510 -1422 1541 -1404
rect 1510 -1432 1556 -1422
rect 1623 -1393 1638 -1378
tri 1248 -1457 1260 -1445 ne
rect 1260 -1450 1270 -1445
tri 1270 -1450 1275 -1445 sw
rect 1159 -1796 1174 -1568
rect 1260 -1606 1275 -1450
rect 1314 -1492 1342 -1436
tri 1434 -1454 1452 -1436 ne
rect 1452 -1456 1474 -1436
tri 1474 -1456 1494 -1436 sw
tri 1510 -1450 1528 -1432 ne
rect 1333 -1526 1342 -1492
rect 1376 -1465 1418 -1464
rect 1376 -1499 1381 -1465
rect 1411 -1499 1418 -1465
rect 1376 -1508 1418 -1499
rect 1452 -1465 1494 -1456
rect 1452 -1499 1459 -1465
rect 1489 -1499 1494 -1465
rect 1452 -1504 1494 -1499
rect 1528 -1492 1556 -1432
tri 1601 -1445 1623 -1423 se
rect 1623 -1430 1638 -1422
tri 1623 -1445 1638 -1430 nw
tri 1595 -1451 1601 -1445 se
rect 1601 -1451 1610 -1445
rect 1314 -1536 1342 -1526
tri 1342 -1536 1366 -1512 sw
rect 1314 -1568 1356 -1536
tri 1373 -1544 1374 -1543 sw
rect 1373 -1568 1374 -1544
tri 1376 -1545 1413 -1508 ne
rect 1413 -1536 1418 -1508
tri 1418 -1536 1444 -1510 sw
rect 1528 -1526 1537 -1492
rect 1528 -1536 1556 -1526
rect 1413 -1545 1497 -1536
tri 1413 -1564 1432 -1545 ne
rect 1432 -1564 1497 -1545
rect 1314 -1590 1374 -1568
rect 1496 -1568 1497 -1564
rect 1514 -1568 1556 -1536
rect 1496 -1590 1556 -1568
rect 1402 -1606 1419 -1592
rect 1451 -1606 1468 -1592
tri 1239 -1642 1261 -1620 se
rect 1261 -1627 1276 -1606
tri 1261 -1642 1276 -1627 nw
rect 1595 -1627 1610 -1451
tri 1610 -1458 1623 -1445 nw
rect 1696 -1526 1711 -1298
tri 1233 -1648 1239 -1642 se
rect 1239 -1648 1248 -1642
rect 1233 -1664 1248 -1648
tri 1248 -1655 1261 -1642 nw
rect 1402 -1650 1419 -1636
rect 1451 -1650 1468 -1636
tri 1595 -1642 1610 -1627 ne
tri 1610 -1642 1632 -1620 sw
rect 1233 -1700 1248 -1692
rect 1314 -1664 1374 -1650
rect 1329 -1674 1374 -1664
rect 1329 -1692 1357 -1674
tri 1233 -1715 1248 -1700 ne
tri 1248 -1715 1270 -1693 sw
rect 1314 -1702 1357 -1692
rect 1372 -1678 1374 -1674
rect 1496 -1664 1556 -1650
tri 1610 -1655 1623 -1642 ne
rect 1623 -1648 1632 -1642
tri 1632 -1648 1638 -1642 sw
rect 1496 -1674 1541 -1664
rect 1372 -1702 1446 -1678
rect 1314 -1706 1446 -1702
tri 1446 -1706 1474 -1678 sw
rect 1496 -1688 1498 -1674
tri 1496 -1690 1498 -1688 ne
rect 1510 -1692 1541 -1674
rect 1510 -1702 1556 -1692
rect 1623 -1663 1638 -1648
tri 1248 -1727 1260 -1715 ne
rect 1260 -1720 1270 -1715
tri 1270 -1720 1275 -1715 sw
rect 1159 -2066 1174 -1838
rect 1260 -1876 1275 -1720
rect 1314 -1762 1342 -1706
tri 1434 -1724 1452 -1706 ne
rect 1452 -1726 1474 -1706
tri 1474 -1726 1494 -1706 sw
tri 1510 -1720 1528 -1702 ne
rect 1333 -1796 1342 -1762
rect 1376 -1735 1418 -1734
rect 1376 -1769 1381 -1735
rect 1411 -1769 1418 -1735
rect 1376 -1778 1418 -1769
rect 1452 -1735 1494 -1726
rect 1452 -1769 1459 -1735
rect 1489 -1769 1494 -1735
rect 1452 -1774 1494 -1769
rect 1528 -1762 1556 -1702
tri 1601 -1715 1623 -1693 se
rect 1623 -1700 1638 -1692
tri 1623 -1715 1638 -1700 nw
tri 1595 -1721 1601 -1715 se
rect 1601 -1721 1610 -1715
rect 1314 -1806 1342 -1796
tri 1342 -1806 1366 -1782 sw
rect 1314 -1838 1356 -1806
tri 1373 -1814 1374 -1813 sw
rect 1373 -1838 1374 -1814
tri 1376 -1815 1413 -1778 ne
rect 1413 -1806 1418 -1778
tri 1418 -1806 1444 -1780 sw
rect 1528 -1796 1537 -1762
rect 1528 -1806 1556 -1796
rect 1413 -1815 1497 -1806
tri 1413 -1834 1432 -1815 ne
rect 1432 -1834 1497 -1815
rect 1314 -1860 1374 -1838
rect 1496 -1838 1497 -1834
rect 1514 -1838 1556 -1806
rect 1496 -1860 1556 -1838
rect 1402 -1876 1419 -1862
rect 1451 -1876 1468 -1862
tri 1239 -1912 1261 -1890 se
rect 1261 -1897 1276 -1876
tri 1261 -1912 1276 -1897 nw
rect 1595 -1897 1610 -1721
tri 1610 -1728 1623 -1715 nw
rect 1696 -1796 1711 -1568
tri 1233 -1918 1239 -1912 se
rect 1239 -1918 1248 -1912
rect 1233 -1934 1248 -1918
tri 1248 -1925 1261 -1912 nw
rect 1402 -1920 1419 -1906
rect 1451 -1920 1468 -1906
tri 1595 -1912 1610 -1897 ne
tri 1610 -1912 1632 -1890 sw
rect 1233 -1970 1248 -1962
rect 1314 -1934 1374 -1920
rect 1329 -1944 1374 -1934
rect 1329 -1962 1357 -1944
tri 1233 -1985 1248 -1970 ne
tri 1248 -1985 1270 -1963 sw
rect 1314 -1972 1357 -1962
rect 1372 -1948 1374 -1944
rect 1496 -1934 1556 -1920
tri 1610 -1925 1623 -1912 ne
rect 1623 -1918 1632 -1912
tri 1632 -1918 1638 -1912 sw
rect 1496 -1944 1541 -1934
rect 1372 -1972 1446 -1948
rect 1314 -1976 1446 -1972
tri 1446 -1976 1474 -1948 sw
rect 1496 -1958 1498 -1944
tri 1496 -1960 1498 -1958 ne
rect 1510 -1962 1541 -1944
rect 1510 -1972 1556 -1962
rect 1623 -1933 1638 -1918
tri 1248 -1997 1260 -1985 ne
rect 1260 -1990 1270 -1985
tri 1270 -1990 1275 -1985 sw
rect 1159 -2146 1174 -2108
rect 1260 -2146 1275 -1990
rect 1314 -2032 1342 -1976
tri 1434 -1994 1452 -1976 ne
rect 1452 -1996 1474 -1976
tri 1474 -1996 1494 -1976 sw
tri 1510 -1990 1528 -1972 ne
rect 1333 -2066 1342 -2032
rect 1376 -2005 1418 -2004
rect 1376 -2039 1381 -2005
rect 1411 -2039 1418 -2005
rect 1376 -2048 1418 -2039
rect 1452 -2005 1494 -1996
rect 1452 -2039 1459 -2005
rect 1489 -2039 1494 -2005
rect 1452 -2044 1494 -2039
rect 1528 -2032 1556 -1972
tri 1601 -1985 1623 -1963 se
rect 1623 -1970 1638 -1962
tri 1623 -1985 1638 -1970 nw
tri 1595 -1991 1601 -1985 se
rect 1601 -1991 1610 -1985
rect 1314 -2076 1342 -2066
tri 1342 -2076 1366 -2052 sw
rect 1314 -2108 1356 -2076
tri 1373 -2084 1374 -2083 sw
rect 1373 -2108 1374 -2084
tri 1376 -2085 1413 -2048 ne
rect 1413 -2076 1418 -2048
tri 1418 -2076 1444 -2050 sw
rect 1528 -2066 1537 -2032
rect 1528 -2076 1556 -2066
rect 1413 -2085 1497 -2076
tri 1413 -2104 1432 -2085 ne
rect 1432 -2104 1497 -2085
rect 1314 -2130 1374 -2108
rect 1496 -2108 1497 -2104
rect 1514 -2108 1556 -2076
rect 1496 -2130 1556 -2108
rect 1402 -2146 1419 -2132
rect 1451 -2146 1468 -2132
rect 1595 -2146 1610 -1991
tri 1610 -1998 1623 -1985 nw
rect 1696 -2066 1711 -1838
rect 1696 -2146 1711 -2108
rect 1739 1984 1754 2174
tri 1819 2138 1841 2160 se
rect 1841 2153 1856 2174
tri 1841 2138 1856 2153 nw
rect 2175 2153 2190 2174
tri 1813 2132 1819 2138 se
rect 1819 2132 1828 2138
rect 1813 2116 1828 2132
tri 1828 2125 1841 2138 nw
rect 1982 2130 1999 2144
rect 2031 2130 2048 2144
tri 2175 2138 2190 2153 ne
tri 2190 2138 2212 2160 sw
rect 1813 2080 1828 2088
rect 1894 2116 1954 2130
rect 1909 2106 1954 2116
rect 1909 2088 1937 2106
tri 1813 2065 1828 2080 ne
tri 1828 2065 1850 2087 sw
rect 1894 2078 1937 2088
rect 1952 2102 1954 2106
rect 2076 2116 2136 2130
tri 2190 2125 2203 2138 ne
rect 2203 2132 2212 2138
tri 2212 2132 2218 2138 sw
rect 2076 2106 2121 2116
rect 1952 2078 2026 2102
rect 1894 2074 2026 2078
tri 2026 2074 2054 2102 sw
rect 2076 2092 2078 2106
tri 2076 2090 2078 2092 ne
rect 2090 2088 2121 2106
rect 2090 2078 2136 2088
rect 2203 2117 2218 2132
tri 1828 2053 1840 2065 ne
rect 1840 2060 1850 2065
tri 1850 2060 1855 2065 sw
rect 1739 1714 1754 1942
rect 1840 1904 1855 2060
rect 1894 2018 1922 2074
tri 2014 2056 2032 2074 ne
rect 2032 2054 2054 2074
tri 2054 2054 2074 2074 sw
tri 2090 2060 2108 2078 ne
rect 1913 1984 1922 2018
rect 1956 2045 1998 2046
rect 1956 2011 1961 2045
rect 1991 2011 1998 2045
rect 1956 2002 1998 2011
rect 2032 2045 2074 2054
rect 2032 2011 2039 2045
rect 2069 2011 2074 2045
rect 2032 2006 2074 2011
rect 2108 2018 2136 2078
tri 2181 2065 2203 2087 se
rect 2203 2080 2218 2088
tri 2203 2065 2218 2080 nw
tri 2175 2059 2181 2065 se
rect 2181 2059 2190 2065
rect 1894 1974 1922 1984
tri 1922 1974 1946 1998 sw
rect 1894 1942 1936 1974
tri 1953 1966 1954 1967 sw
rect 1953 1942 1954 1966
tri 1956 1965 1993 2002 ne
rect 1993 1974 1998 2002
tri 1998 1974 2024 2000 sw
rect 2108 1984 2117 2018
rect 2108 1974 2136 1984
rect 1993 1965 2077 1974
tri 1993 1946 2012 1965 ne
rect 2012 1946 2077 1965
rect 1894 1920 1954 1942
rect 2076 1942 2077 1946
rect 2094 1942 2136 1974
rect 2076 1920 2136 1942
rect 1982 1904 1999 1918
rect 2031 1904 2048 1918
tri 1819 1868 1841 1890 se
rect 1841 1883 1856 1904
tri 1841 1868 1856 1883 nw
rect 2175 1883 2190 2059
tri 2190 2052 2203 2065 nw
rect 2276 1984 2291 2174
tri 1813 1862 1819 1868 se
rect 1819 1862 1828 1868
rect 1813 1846 1828 1862
tri 1828 1855 1841 1868 nw
rect 1982 1860 1999 1874
rect 2031 1860 2048 1874
tri 2175 1868 2190 1883 ne
tri 2190 1868 2212 1890 sw
rect 1813 1810 1828 1818
rect 1894 1846 1954 1860
rect 1909 1836 1954 1846
rect 1909 1818 1937 1836
tri 1813 1795 1828 1810 ne
tri 1828 1795 1850 1817 sw
rect 1894 1808 1937 1818
rect 1952 1832 1954 1836
rect 2076 1846 2136 1860
tri 2190 1855 2203 1868 ne
rect 2203 1862 2212 1868
tri 2212 1862 2218 1868 sw
rect 2076 1836 2121 1846
rect 1952 1808 2026 1832
rect 1894 1804 2026 1808
tri 2026 1804 2054 1832 sw
rect 2076 1822 2078 1836
tri 2076 1820 2078 1822 ne
rect 2090 1818 2121 1836
rect 2090 1808 2136 1818
rect 2203 1847 2218 1862
tri 1828 1783 1840 1795 ne
rect 1840 1790 1850 1795
tri 1850 1790 1855 1795 sw
rect 1739 1444 1754 1672
rect 1840 1634 1855 1790
rect 1894 1748 1922 1804
tri 2014 1786 2032 1804 ne
rect 2032 1784 2054 1804
tri 2054 1784 2074 1804 sw
tri 2090 1790 2108 1808 ne
rect 1913 1714 1922 1748
rect 1956 1775 1998 1776
rect 1956 1741 1961 1775
rect 1991 1741 1998 1775
rect 1956 1732 1998 1741
rect 2032 1775 2074 1784
rect 2032 1741 2039 1775
rect 2069 1741 2074 1775
rect 2032 1736 2074 1741
rect 2108 1748 2136 1808
tri 2181 1795 2203 1817 se
rect 2203 1810 2218 1818
tri 2203 1795 2218 1810 nw
tri 2175 1789 2181 1795 se
rect 2181 1789 2190 1795
rect 1894 1704 1922 1714
tri 1922 1704 1946 1728 sw
rect 1894 1672 1936 1704
tri 1953 1696 1954 1697 sw
rect 1953 1672 1954 1696
tri 1956 1695 1993 1732 ne
rect 1993 1704 1998 1732
tri 1998 1704 2024 1730 sw
rect 2108 1714 2117 1748
rect 2108 1704 2136 1714
rect 1993 1695 2077 1704
tri 1993 1676 2012 1695 ne
rect 2012 1676 2077 1695
rect 1894 1650 1954 1672
rect 2076 1672 2077 1676
rect 2094 1672 2136 1704
rect 2076 1650 2136 1672
rect 1982 1634 1999 1648
rect 2031 1634 2048 1648
tri 1819 1598 1841 1620 se
rect 1841 1613 1856 1634
tri 1841 1598 1856 1613 nw
rect 2175 1613 2190 1789
tri 2190 1782 2203 1795 nw
rect 2276 1714 2291 1942
tri 1813 1592 1819 1598 se
rect 1819 1592 1828 1598
rect 1813 1576 1828 1592
tri 1828 1585 1841 1598 nw
rect 1982 1590 1999 1604
rect 2031 1590 2048 1604
tri 2175 1598 2190 1613 ne
tri 2190 1598 2212 1620 sw
rect 1813 1540 1828 1548
rect 1894 1576 1954 1590
rect 1909 1566 1954 1576
rect 1909 1548 1937 1566
tri 1813 1525 1828 1540 ne
tri 1828 1525 1850 1547 sw
rect 1894 1538 1937 1548
rect 1952 1562 1954 1566
rect 2076 1576 2136 1590
tri 2190 1585 2203 1598 ne
rect 2203 1592 2212 1598
tri 2212 1592 2218 1598 sw
rect 2076 1566 2121 1576
rect 1952 1538 2026 1562
rect 1894 1534 2026 1538
tri 2026 1534 2054 1562 sw
rect 2076 1552 2078 1566
tri 2076 1550 2078 1552 ne
rect 2090 1548 2121 1566
rect 2090 1538 2136 1548
rect 2203 1577 2218 1592
tri 1828 1513 1840 1525 ne
rect 1840 1520 1850 1525
tri 1850 1520 1855 1525 sw
rect 1739 1174 1754 1402
rect 1840 1364 1855 1520
rect 1894 1478 1922 1534
tri 2014 1516 2032 1534 ne
rect 2032 1514 2054 1534
tri 2054 1514 2074 1534 sw
tri 2090 1520 2108 1538 ne
rect 1913 1444 1922 1478
rect 1956 1505 1998 1506
rect 1956 1471 1961 1505
rect 1991 1471 1998 1505
rect 1956 1462 1998 1471
rect 2032 1505 2074 1514
rect 2032 1471 2039 1505
rect 2069 1471 2074 1505
rect 2032 1466 2074 1471
rect 2108 1478 2136 1538
tri 2181 1525 2203 1547 se
rect 2203 1540 2218 1548
tri 2203 1525 2218 1540 nw
tri 2175 1519 2181 1525 se
rect 2181 1519 2190 1525
rect 1894 1434 1922 1444
tri 1922 1434 1946 1458 sw
rect 1894 1402 1936 1434
tri 1953 1426 1954 1427 sw
rect 1953 1402 1954 1426
tri 1956 1425 1993 1462 ne
rect 1993 1434 1998 1462
tri 1998 1434 2024 1460 sw
rect 2108 1444 2117 1478
rect 2108 1434 2136 1444
rect 1993 1425 2077 1434
tri 1993 1406 2012 1425 ne
rect 2012 1406 2077 1425
rect 1894 1380 1954 1402
rect 2076 1402 2077 1406
rect 2094 1402 2136 1434
rect 2076 1380 2136 1402
rect 1982 1364 1999 1378
rect 2031 1364 2048 1378
tri 1819 1328 1841 1350 se
rect 1841 1343 1856 1364
tri 1841 1328 1856 1343 nw
rect 2175 1343 2190 1519
tri 2190 1512 2203 1525 nw
rect 2276 1444 2291 1672
tri 1813 1322 1819 1328 se
rect 1819 1322 1828 1328
rect 1813 1306 1828 1322
tri 1828 1315 1841 1328 nw
rect 1982 1320 1999 1334
rect 2031 1320 2048 1334
tri 2175 1328 2190 1343 ne
tri 2190 1328 2212 1350 sw
rect 1813 1270 1828 1278
rect 1894 1306 1954 1320
rect 1909 1296 1954 1306
rect 1909 1278 1937 1296
tri 1813 1255 1828 1270 ne
tri 1828 1255 1850 1277 sw
rect 1894 1268 1937 1278
rect 1952 1292 1954 1296
rect 2076 1306 2136 1320
tri 2190 1315 2203 1328 ne
rect 2203 1322 2212 1328
tri 2212 1322 2218 1328 sw
rect 2076 1296 2121 1306
rect 1952 1268 2026 1292
rect 1894 1264 2026 1268
tri 2026 1264 2054 1292 sw
rect 2076 1282 2078 1296
tri 2076 1280 2078 1282 ne
rect 2090 1278 2121 1296
rect 2090 1268 2136 1278
rect 2203 1307 2218 1322
tri 1828 1243 1840 1255 ne
rect 1840 1250 1850 1255
tri 1850 1250 1855 1255 sw
rect 1739 904 1754 1132
rect 1840 1094 1855 1250
rect 1894 1208 1922 1264
tri 2014 1246 2032 1264 ne
rect 2032 1244 2054 1264
tri 2054 1244 2074 1264 sw
tri 2090 1250 2108 1268 ne
rect 1913 1174 1922 1208
rect 1956 1235 1998 1236
rect 1956 1201 1961 1235
rect 1991 1201 1998 1235
rect 1956 1192 1998 1201
rect 2032 1235 2074 1244
rect 2032 1201 2039 1235
rect 2069 1201 2074 1235
rect 2032 1196 2074 1201
rect 2108 1208 2136 1268
tri 2181 1255 2203 1277 se
rect 2203 1270 2218 1278
tri 2203 1255 2218 1270 nw
tri 2175 1249 2181 1255 se
rect 2181 1249 2190 1255
rect 1894 1164 1922 1174
tri 1922 1164 1946 1188 sw
rect 1894 1132 1936 1164
tri 1953 1156 1954 1157 sw
rect 1953 1132 1954 1156
tri 1956 1155 1993 1192 ne
rect 1993 1164 1998 1192
tri 1998 1164 2024 1190 sw
rect 2108 1174 2117 1208
rect 2108 1164 2136 1174
rect 1993 1155 2077 1164
tri 1993 1136 2012 1155 ne
rect 2012 1136 2077 1155
rect 1894 1110 1954 1132
rect 2076 1132 2077 1136
rect 2094 1132 2136 1164
rect 2076 1110 2136 1132
rect 1982 1094 1999 1108
rect 2031 1094 2048 1108
tri 1819 1058 1841 1080 se
rect 1841 1073 1856 1094
tri 1841 1058 1856 1073 nw
rect 2175 1073 2190 1249
tri 2190 1242 2203 1255 nw
rect 2276 1174 2291 1402
tri 1813 1052 1819 1058 se
rect 1819 1052 1828 1058
rect 1813 1036 1828 1052
tri 1828 1045 1841 1058 nw
rect 1982 1050 1999 1064
rect 2031 1050 2048 1064
tri 2175 1058 2190 1073 ne
tri 2190 1058 2212 1080 sw
rect 1813 1000 1828 1008
rect 1894 1036 1954 1050
rect 1909 1026 1954 1036
rect 1909 1008 1937 1026
tri 1813 985 1828 1000 ne
tri 1828 985 1850 1007 sw
rect 1894 998 1937 1008
rect 1952 1022 1954 1026
rect 2076 1036 2136 1050
tri 2190 1045 2203 1058 ne
rect 2203 1052 2212 1058
tri 2212 1052 2218 1058 sw
rect 2076 1026 2121 1036
rect 1952 998 2026 1022
rect 1894 994 2026 998
tri 2026 994 2054 1022 sw
rect 2076 1012 2078 1026
tri 2076 1010 2078 1012 ne
rect 2090 1008 2121 1026
rect 2090 998 2136 1008
rect 2203 1037 2218 1052
tri 1828 973 1840 985 ne
rect 1840 980 1850 985
tri 1850 980 1855 985 sw
rect 1739 634 1754 862
rect 1840 824 1855 980
rect 1894 938 1922 994
tri 2014 976 2032 994 ne
rect 2032 974 2054 994
tri 2054 974 2074 994 sw
tri 2090 980 2108 998 ne
rect 1913 904 1922 938
rect 1956 965 1998 966
rect 1956 931 1961 965
rect 1991 931 1998 965
rect 1956 922 1998 931
rect 2032 965 2074 974
rect 2032 931 2039 965
rect 2069 931 2074 965
rect 2032 926 2074 931
rect 2108 938 2136 998
tri 2181 985 2203 1007 se
rect 2203 1000 2218 1008
tri 2203 985 2218 1000 nw
tri 2175 979 2181 985 se
rect 2181 979 2190 985
rect 1894 894 1922 904
tri 1922 894 1946 918 sw
rect 1894 862 1936 894
tri 1953 886 1954 887 sw
rect 1953 862 1954 886
tri 1956 885 1993 922 ne
rect 1993 894 1998 922
tri 1998 894 2024 920 sw
rect 2108 904 2117 938
rect 2108 894 2136 904
rect 1993 885 2077 894
tri 1993 866 2012 885 ne
rect 2012 866 2077 885
rect 1894 840 1954 862
rect 2076 862 2077 866
rect 2094 862 2136 894
rect 2076 840 2136 862
rect 1982 824 1999 838
rect 2031 824 2048 838
tri 1819 788 1841 810 se
rect 1841 803 1856 824
tri 1841 788 1856 803 nw
rect 2175 803 2190 979
tri 2190 972 2203 985 nw
rect 2276 904 2291 1132
tri 1813 782 1819 788 se
rect 1819 782 1828 788
rect 1813 766 1828 782
tri 1828 775 1841 788 nw
rect 1982 780 1999 794
rect 2031 780 2048 794
tri 2175 788 2190 803 ne
tri 2190 788 2212 810 sw
rect 1813 730 1828 738
rect 1894 766 1954 780
rect 1909 756 1954 766
rect 1909 738 1937 756
tri 1813 715 1828 730 ne
tri 1828 715 1850 737 sw
rect 1894 728 1937 738
rect 1952 752 1954 756
rect 2076 766 2136 780
tri 2190 775 2203 788 ne
rect 2203 782 2212 788
tri 2212 782 2218 788 sw
rect 2076 756 2121 766
rect 1952 728 2026 752
rect 1894 724 2026 728
tri 2026 724 2054 752 sw
rect 2076 742 2078 756
tri 2076 740 2078 742 ne
rect 2090 738 2121 756
rect 2090 728 2136 738
rect 2203 767 2218 782
tri 1828 703 1840 715 ne
rect 1840 710 1850 715
tri 1850 710 1855 715 sw
rect 1739 364 1754 592
rect 1840 554 1855 710
rect 1894 668 1922 724
tri 2014 706 2032 724 ne
rect 2032 704 2054 724
tri 2054 704 2074 724 sw
tri 2090 710 2108 728 ne
rect 1913 634 1922 668
rect 1956 695 1998 696
rect 1956 661 1961 695
rect 1991 661 1998 695
rect 1956 652 1998 661
rect 2032 695 2074 704
rect 2032 661 2039 695
rect 2069 661 2074 695
rect 2032 656 2074 661
rect 2108 668 2136 728
tri 2181 715 2203 737 se
rect 2203 730 2218 738
tri 2203 715 2218 730 nw
tri 2175 709 2181 715 se
rect 2181 709 2190 715
rect 1894 624 1922 634
tri 1922 624 1946 648 sw
rect 1894 592 1936 624
tri 1953 616 1954 617 sw
rect 1953 592 1954 616
tri 1956 615 1993 652 ne
rect 1993 624 1998 652
tri 1998 624 2024 650 sw
rect 2108 634 2117 668
rect 2108 624 2136 634
rect 1993 615 2077 624
tri 1993 596 2012 615 ne
rect 2012 596 2077 615
rect 1894 570 1954 592
rect 2076 592 2077 596
rect 2094 592 2136 624
rect 2076 570 2136 592
rect 1982 554 1999 568
rect 2031 554 2048 568
tri 1819 518 1841 540 se
rect 1841 533 1856 554
tri 1841 518 1856 533 nw
rect 2175 533 2190 709
tri 2190 702 2203 715 nw
rect 2276 634 2291 862
tri 1813 512 1819 518 se
rect 1819 512 1828 518
rect 1813 496 1828 512
tri 1828 505 1841 518 nw
rect 1982 510 1999 524
rect 2031 510 2048 524
tri 2175 518 2190 533 ne
tri 2190 518 2212 540 sw
rect 1813 460 1828 468
rect 1894 496 1954 510
rect 1909 486 1954 496
rect 1909 468 1937 486
tri 1813 445 1828 460 ne
tri 1828 445 1850 467 sw
rect 1894 458 1937 468
rect 1952 482 1954 486
rect 2076 496 2136 510
tri 2190 505 2203 518 ne
rect 2203 512 2212 518
tri 2212 512 2218 518 sw
rect 2076 486 2121 496
rect 1952 458 2026 482
rect 1894 454 2026 458
tri 2026 454 2054 482 sw
rect 2076 472 2078 486
tri 2076 470 2078 472 ne
rect 2090 468 2121 486
rect 2090 458 2136 468
rect 2203 497 2218 512
tri 1828 433 1840 445 ne
rect 1840 440 1850 445
tri 1850 440 1855 445 sw
rect 1739 94 1754 322
rect 1840 284 1855 440
rect 1894 398 1922 454
tri 2014 436 2032 454 ne
rect 2032 434 2054 454
tri 2054 434 2074 454 sw
tri 2090 440 2108 458 ne
rect 1913 364 1922 398
rect 1956 425 1998 426
rect 1956 391 1961 425
rect 1991 391 1998 425
rect 1956 382 1998 391
rect 2032 425 2074 434
rect 2032 391 2039 425
rect 2069 391 2074 425
rect 2032 386 2074 391
rect 2108 398 2136 458
tri 2181 445 2203 467 se
rect 2203 460 2218 468
tri 2203 445 2218 460 nw
tri 2175 439 2181 445 se
rect 2181 439 2190 445
rect 1894 354 1922 364
tri 1922 354 1946 378 sw
rect 1894 322 1936 354
tri 1953 346 1954 347 sw
rect 1953 322 1954 346
tri 1956 345 1993 382 ne
rect 1993 354 1998 382
tri 1998 354 2024 380 sw
rect 2108 364 2117 398
rect 2108 354 2136 364
rect 1993 345 2077 354
tri 1993 326 2012 345 ne
rect 2012 326 2077 345
rect 1894 300 1954 322
rect 2076 322 2077 326
rect 2094 322 2136 354
rect 2076 300 2136 322
rect 1982 284 1999 298
rect 2031 284 2048 298
tri 1819 248 1841 270 se
rect 1841 263 1856 284
tri 1841 248 1856 263 nw
rect 2175 263 2190 439
tri 2190 432 2203 445 nw
rect 2276 364 2291 592
tri 1813 242 1819 248 se
rect 1819 242 1828 248
rect 1813 226 1828 242
tri 1828 235 1841 248 nw
rect 1982 240 1999 254
rect 2031 240 2048 254
tri 2175 248 2190 263 ne
tri 2190 248 2212 270 sw
rect 1813 190 1828 198
rect 1894 226 1954 240
rect 1909 216 1954 226
rect 1909 198 1937 216
tri 1813 175 1828 190 ne
tri 1828 175 1850 197 sw
rect 1894 188 1937 198
rect 1952 212 1954 216
rect 2076 226 2136 240
tri 2190 235 2203 248 ne
rect 2203 242 2212 248
tri 2212 242 2218 248 sw
rect 2076 216 2121 226
rect 1952 188 2026 212
rect 1894 184 2026 188
tri 2026 184 2054 212 sw
rect 2076 202 2078 216
tri 2076 200 2078 202 ne
rect 2090 198 2121 216
rect 2090 188 2136 198
rect 2203 227 2218 242
tri 1828 163 1840 175 ne
rect 1840 170 1850 175
tri 1850 170 1855 175 sw
rect 1739 -176 1754 52
rect 1840 14 1855 170
rect 1894 128 1922 184
tri 2014 166 2032 184 ne
rect 2032 164 2054 184
tri 2054 164 2074 184 sw
tri 2090 170 2108 188 ne
rect 1913 94 1922 128
rect 1956 155 1998 156
rect 1956 121 1961 155
rect 1991 121 1998 155
rect 1956 112 1998 121
rect 2032 155 2074 164
rect 2032 121 2039 155
rect 2069 121 2074 155
rect 2032 116 2074 121
rect 2108 128 2136 188
tri 2181 175 2203 197 se
rect 2203 190 2218 198
tri 2203 175 2218 190 nw
tri 2175 169 2181 175 se
rect 2181 169 2190 175
rect 1894 84 1922 94
tri 1922 84 1946 108 sw
rect 1894 52 1936 84
tri 1953 76 1954 77 sw
rect 1953 52 1954 76
tri 1956 75 1993 112 ne
rect 1993 84 1998 112
tri 1998 84 2024 110 sw
rect 2108 94 2117 128
rect 2108 84 2136 94
rect 1993 75 2077 84
tri 1993 56 2012 75 ne
rect 2012 56 2077 75
rect 1894 30 1954 52
rect 2076 52 2077 56
rect 2094 52 2136 84
rect 2076 30 2136 52
rect 1982 14 1999 28
rect 2031 14 2048 28
tri 1819 -22 1841 0 se
rect 1841 -7 1856 14
tri 1841 -22 1856 -7 nw
rect 2175 -7 2190 169
tri 2190 162 2203 175 nw
rect 2276 94 2291 322
tri 1813 -28 1819 -22 se
rect 1819 -28 1828 -22
rect 1813 -44 1828 -28
tri 1828 -35 1841 -22 nw
rect 1982 -30 1999 -16
rect 2031 -30 2048 -16
tri 2175 -22 2190 -7 ne
tri 2190 -22 2212 0 sw
rect 1813 -80 1828 -72
rect 1894 -44 1954 -30
rect 1909 -54 1954 -44
rect 1909 -72 1937 -54
tri 1813 -95 1828 -80 ne
tri 1828 -95 1850 -73 sw
rect 1894 -82 1937 -72
rect 1952 -58 1954 -54
rect 2076 -44 2136 -30
tri 2190 -35 2203 -22 ne
rect 2203 -28 2212 -22
tri 2212 -28 2218 -22 sw
rect 2076 -54 2121 -44
rect 1952 -82 2026 -58
rect 1894 -86 2026 -82
tri 2026 -86 2054 -58 sw
rect 2076 -68 2078 -54
tri 2076 -70 2078 -68 ne
rect 2090 -72 2121 -54
rect 2090 -82 2136 -72
rect 2203 -43 2218 -28
tri 1828 -107 1840 -95 ne
rect 1840 -100 1850 -95
tri 1850 -100 1855 -95 sw
rect 1739 -446 1754 -218
rect 1840 -256 1855 -100
rect 1894 -142 1922 -86
tri 2014 -104 2032 -86 ne
rect 2032 -106 2054 -86
tri 2054 -106 2074 -86 sw
tri 2090 -100 2108 -82 ne
rect 1913 -176 1922 -142
rect 1956 -115 1998 -114
rect 1956 -149 1961 -115
rect 1991 -149 1998 -115
rect 1956 -158 1998 -149
rect 2032 -115 2074 -106
rect 2032 -149 2039 -115
rect 2069 -149 2074 -115
rect 2032 -154 2074 -149
rect 2108 -142 2136 -82
tri 2181 -95 2203 -73 se
rect 2203 -80 2218 -72
tri 2203 -95 2218 -80 nw
tri 2175 -101 2181 -95 se
rect 2181 -101 2190 -95
rect 1894 -186 1922 -176
tri 1922 -186 1946 -162 sw
rect 1894 -218 1936 -186
tri 1953 -194 1954 -193 sw
rect 1953 -218 1954 -194
tri 1956 -195 1993 -158 ne
rect 1993 -186 1998 -158
tri 1998 -186 2024 -160 sw
rect 2108 -176 2117 -142
rect 2108 -186 2136 -176
rect 1993 -195 2077 -186
tri 1993 -214 2012 -195 ne
rect 2012 -214 2077 -195
rect 1894 -240 1954 -218
rect 2076 -218 2077 -214
rect 2094 -218 2136 -186
rect 2076 -240 2136 -218
rect 1982 -256 1999 -242
rect 2031 -256 2048 -242
tri 1819 -292 1841 -270 se
rect 1841 -277 1856 -256
tri 1841 -292 1856 -277 nw
rect 2175 -277 2190 -101
tri 2190 -108 2203 -95 nw
rect 2276 -176 2291 52
tri 1813 -298 1819 -292 se
rect 1819 -298 1828 -292
rect 1813 -314 1828 -298
tri 1828 -305 1841 -292 nw
rect 1982 -300 1999 -286
rect 2031 -300 2048 -286
tri 2175 -292 2190 -277 ne
tri 2190 -292 2212 -270 sw
rect 1813 -350 1828 -342
rect 1894 -314 1954 -300
rect 1909 -324 1954 -314
rect 1909 -342 1937 -324
tri 1813 -365 1828 -350 ne
tri 1828 -365 1850 -343 sw
rect 1894 -352 1937 -342
rect 1952 -328 1954 -324
rect 2076 -314 2136 -300
tri 2190 -305 2203 -292 ne
rect 2203 -298 2212 -292
tri 2212 -298 2218 -292 sw
rect 2076 -324 2121 -314
rect 1952 -352 2026 -328
rect 1894 -356 2026 -352
tri 2026 -356 2054 -328 sw
rect 2076 -338 2078 -324
tri 2076 -340 2078 -338 ne
rect 2090 -342 2121 -324
rect 2090 -352 2136 -342
rect 2203 -313 2218 -298
tri 1828 -377 1840 -365 ne
rect 1840 -370 1850 -365
tri 1850 -370 1855 -365 sw
rect 1739 -716 1754 -488
rect 1840 -526 1855 -370
rect 1894 -412 1922 -356
tri 2014 -374 2032 -356 ne
rect 2032 -376 2054 -356
tri 2054 -376 2074 -356 sw
tri 2090 -370 2108 -352 ne
rect 1913 -446 1922 -412
rect 1956 -385 1998 -384
rect 1956 -419 1961 -385
rect 1991 -419 1998 -385
rect 1956 -428 1998 -419
rect 2032 -385 2074 -376
rect 2032 -419 2039 -385
rect 2069 -419 2074 -385
rect 2032 -424 2074 -419
rect 2108 -412 2136 -352
tri 2181 -365 2203 -343 se
rect 2203 -350 2218 -342
tri 2203 -365 2218 -350 nw
tri 2175 -371 2181 -365 se
rect 2181 -371 2190 -365
rect 1894 -456 1922 -446
tri 1922 -456 1946 -432 sw
rect 1894 -488 1936 -456
tri 1953 -464 1954 -463 sw
rect 1953 -488 1954 -464
tri 1956 -465 1993 -428 ne
rect 1993 -456 1998 -428
tri 1998 -456 2024 -430 sw
rect 2108 -446 2117 -412
rect 2108 -456 2136 -446
rect 1993 -465 2077 -456
tri 1993 -484 2012 -465 ne
rect 2012 -484 2077 -465
rect 1894 -510 1954 -488
rect 2076 -488 2077 -484
rect 2094 -488 2136 -456
rect 2076 -510 2136 -488
rect 1982 -526 1999 -512
rect 2031 -526 2048 -512
tri 1819 -562 1841 -540 se
rect 1841 -547 1856 -526
tri 1841 -562 1856 -547 nw
rect 2175 -547 2190 -371
tri 2190 -378 2203 -365 nw
rect 2276 -446 2291 -218
tri 1813 -568 1819 -562 se
rect 1819 -568 1828 -562
rect 1813 -584 1828 -568
tri 1828 -575 1841 -562 nw
rect 1982 -570 1999 -556
rect 2031 -570 2048 -556
tri 2175 -562 2190 -547 ne
tri 2190 -562 2212 -540 sw
rect 1813 -620 1828 -612
rect 1894 -584 1954 -570
rect 1909 -594 1954 -584
rect 1909 -612 1937 -594
tri 1813 -635 1828 -620 ne
tri 1828 -635 1850 -613 sw
rect 1894 -622 1937 -612
rect 1952 -598 1954 -594
rect 2076 -584 2136 -570
tri 2190 -575 2203 -562 ne
rect 2203 -568 2212 -562
tri 2212 -568 2218 -562 sw
rect 2076 -594 2121 -584
rect 1952 -622 2026 -598
rect 1894 -626 2026 -622
tri 2026 -626 2054 -598 sw
rect 2076 -608 2078 -594
tri 2076 -610 2078 -608 ne
rect 2090 -612 2121 -594
rect 2090 -622 2136 -612
rect 2203 -583 2218 -568
tri 1828 -647 1840 -635 ne
rect 1840 -640 1850 -635
tri 1850 -640 1855 -635 sw
rect 1739 -986 1754 -758
rect 1840 -796 1855 -640
rect 1894 -682 1922 -626
tri 2014 -644 2032 -626 ne
rect 2032 -646 2054 -626
tri 2054 -646 2074 -626 sw
tri 2090 -640 2108 -622 ne
rect 1913 -716 1922 -682
rect 1956 -655 1998 -654
rect 1956 -689 1961 -655
rect 1991 -689 1998 -655
rect 1956 -698 1998 -689
rect 2032 -655 2074 -646
rect 2032 -689 2039 -655
rect 2069 -689 2074 -655
rect 2032 -694 2074 -689
rect 2108 -682 2136 -622
tri 2181 -635 2203 -613 se
rect 2203 -620 2218 -612
tri 2203 -635 2218 -620 nw
tri 2175 -641 2181 -635 se
rect 2181 -641 2190 -635
rect 1894 -726 1922 -716
tri 1922 -726 1946 -702 sw
rect 1894 -758 1936 -726
tri 1953 -734 1954 -733 sw
rect 1953 -758 1954 -734
tri 1956 -735 1993 -698 ne
rect 1993 -726 1998 -698
tri 1998 -726 2024 -700 sw
rect 2108 -716 2117 -682
rect 2108 -726 2136 -716
rect 1993 -735 2077 -726
tri 1993 -754 2012 -735 ne
rect 2012 -754 2077 -735
rect 1894 -780 1954 -758
rect 2076 -758 2077 -754
rect 2094 -758 2136 -726
rect 2076 -780 2136 -758
rect 1982 -796 1999 -782
rect 2031 -796 2048 -782
tri 1819 -832 1841 -810 se
rect 1841 -817 1856 -796
tri 1841 -832 1856 -817 nw
rect 2175 -817 2190 -641
tri 2190 -648 2203 -635 nw
rect 2276 -716 2291 -488
tri 1813 -838 1819 -832 se
rect 1819 -838 1828 -832
rect 1813 -854 1828 -838
tri 1828 -845 1841 -832 nw
rect 1982 -840 1999 -826
rect 2031 -840 2048 -826
tri 2175 -832 2190 -817 ne
tri 2190 -832 2212 -810 sw
rect 1813 -890 1828 -882
rect 1894 -854 1954 -840
rect 1909 -864 1954 -854
rect 1909 -882 1937 -864
tri 1813 -905 1828 -890 ne
tri 1828 -905 1850 -883 sw
rect 1894 -892 1937 -882
rect 1952 -868 1954 -864
rect 2076 -854 2136 -840
tri 2190 -845 2203 -832 ne
rect 2203 -838 2212 -832
tri 2212 -838 2218 -832 sw
rect 2076 -864 2121 -854
rect 1952 -892 2026 -868
rect 1894 -896 2026 -892
tri 2026 -896 2054 -868 sw
rect 2076 -878 2078 -864
tri 2076 -880 2078 -878 ne
rect 2090 -882 2121 -864
rect 2090 -892 2136 -882
rect 2203 -853 2218 -838
tri 1828 -917 1840 -905 ne
rect 1840 -910 1850 -905
tri 1850 -910 1855 -905 sw
rect 1739 -1256 1754 -1028
rect 1840 -1066 1855 -910
rect 1894 -952 1922 -896
tri 2014 -914 2032 -896 ne
rect 2032 -916 2054 -896
tri 2054 -916 2074 -896 sw
tri 2090 -910 2108 -892 ne
rect 1913 -986 1922 -952
rect 1956 -925 1998 -924
rect 1956 -959 1961 -925
rect 1991 -959 1998 -925
rect 1956 -968 1998 -959
rect 2032 -925 2074 -916
rect 2032 -959 2039 -925
rect 2069 -959 2074 -925
rect 2032 -964 2074 -959
rect 2108 -952 2136 -892
tri 2181 -905 2203 -883 se
rect 2203 -890 2218 -882
tri 2203 -905 2218 -890 nw
tri 2175 -911 2181 -905 se
rect 2181 -911 2190 -905
rect 1894 -996 1922 -986
tri 1922 -996 1946 -972 sw
rect 1894 -1028 1936 -996
tri 1953 -1004 1954 -1003 sw
rect 1953 -1028 1954 -1004
tri 1956 -1005 1993 -968 ne
rect 1993 -996 1998 -968
tri 1998 -996 2024 -970 sw
rect 2108 -986 2117 -952
rect 2108 -996 2136 -986
rect 1993 -1005 2077 -996
tri 1993 -1024 2012 -1005 ne
rect 2012 -1024 2077 -1005
rect 1894 -1050 1954 -1028
rect 2076 -1028 2077 -1024
rect 2094 -1028 2136 -996
rect 2076 -1050 2136 -1028
rect 1982 -1066 1999 -1052
rect 2031 -1066 2048 -1052
tri 1819 -1102 1841 -1080 se
rect 1841 -1087 1856 -1066
tri 1841 -1102 1856 -1087 nw
rect 2175 -1087 2190 -911
tri 2190 -918 2203 -905 nw
rect 2276 -986 2291 -758
tri 1813 -1108 1819 -1102 se
rect 1819 -1108 1828 -1102
rect 1813 -1124 1828 -1108
tri 1828 -1115 1841 -1102 nw
rect 1982 -1110 1999 -1096
rect 2031 -1110 2048 -1096
tri 2175 -1102 2190 -1087 ne
tri 2190 -1102 2212 -1080 sw
rect 1813 -1160 1828 -1152
rect 1894 -1124 1954 -1110
rect 1909 -1134 1954 -1124
rect 1909 -1152 1937 -1134
tri 1813 -1175 1828 -1160 ne
tri 1828 -1175 1850 -1153 sw
rect 1894 -1162 1937 -1152
rect 1952 -1138 1954 -1134
rect 2076 -1124 2136 -1110
tri 2190 -1115 2203 -1102 ne
rect 2203 -1108 2212 -1102
tri 2212 -1108 2218 -1102 sw
rect 2076 -1134 2121 -1124
rect 1952 -1162 2026 -1138
rect 1894 -1166 2026 -1162
tri 2026 -1166 2054 -1138 sw
rect 2076 -1148 2078 -1134
tri 2076 -1150 2078 -1148 ne
rect 2090 -1152 2121 -1134
rect 2090 -1162 2136 -1152
rect 2203 -1123 2218 -1108
tri 1828 -1187 1840 -1175 ne
rect 1840 -1180 1850 -1175
tri 1850 -1180 1855 -1175 sw
rect 1739 -1526 1754 -1298
rect 1840 -1336 1855 -1180
rect 1894 -1222 1922 -1166
tri 2014 -1184 2032 -1166 ne
rect 2032 -1186 2054 -1166
tri 2054 -1186 2074 -1166 sw
tri 2090 -1180 2108 -1162 ne
rect 1913 -1256 1922 -1222
rect 1956 -1195 1998 -1194
rect 1956 -1229 1961 -1195
rect 1991 -1229 1998 -1195
rect 1956 -1238 1998 -1229
rect 2032 -1195 2074 -1186
rect 2032 -1229 2039 -1195
rect 2069 -1229 2074 -1195
rect 2032 -1234 2074 -1229
rect 2108 -1222 2136 -1162
tri 2181 -1175 2203 -1153 se
rect 2203 -1160 2218 -1152
tri 2203 -1175 2218 -1160 nw
tri 2175 -1181 2181 -1175 se
rect 2181 -1181 2190 -1175
rect 1894 -1266 1922 -1256
tri 1922 -1266 1946 -1242 sw
rect 1894 -1298 1936 -1266
tri 1953 -1274 1954 -1273 sw
rect 1953 -1298 1954 -1274
tri 1956 -1275 1993 -1238 ne
rect 1993 -1266 1998 -1238
tri 1998 -1266 2024 -1240 sw
rect 2108 -1256 2117 -1222
rect 2108 -1266 2136 -1256
rect 1993 -1275 2077 -1266
tri 1993 -1294 2012 -1275 ne
rect 2012 -1294 2077 -1275
rect 1894 -1320 1954 -1298
rect 2076 -1298 2077 -1294
rect 2094 -1298 2136 -1266
rect 2076 -1320 2136 -1298
rect 1982 -1336 1999 -1322
rect 2031 -1336 2048 -1322
tri 1819 -1372 1841 -1350 se
rect 1841 -1357 1856 -1336
tri 1841 -1372 1856 -1357 nw
rect 2175 -1357 2190 -1181
tri 2190 -1188 2203 -1175 nw
rect 2276 -1256 2291 -1028
tri 1813 -1378 1819 -1372 se
rect 1819 -1378 1828 -1372
rect 1813 -1394 1828 -1378
tri 1828 -1385 1841 -1372 nw
rect 1982 -1380 1999 -1366
rect 2031 -1380 2048 -1366
tri 2175 -1372 2190 -1357 ne
tri 2190 -1372 2212 -1350 sw
rect 1813 -1430 1828 -1422
rect 1894 -1394 1954 -1380
rect 1909 -1404 1954 -1394
rect 1909 -1422 1937 -1404
tri 1813 -1445 1828 -1430 ne
tri 1828 -1445 1850 -1423 sw
rect 1894 -1432 1937 -1422
rect 1952 -1408 1954 -1404
rect 2076 -1394 2136 -1380
tri 2190 -1385 2203 -1372 ne
rect 2203 -1378 2212 -1372
tri 2212 -1378 2218 -1372 sw
rect 2076 -1404 2121 -1394
rect 1952 -1432 2026 -1408
rect 1894 -1436 2026 -1432
tri 2026 -1436 2054 -1408 sw
rect 2076 -1418 2078 -1404
tri 2076 -1420 2078 -1418 ne
rect 2090 -1422 2121 -1404
rect 2090 -1432 2136 -1422
rect 2203 -1393 2218 -1378
tri 1828 -1457 1840 -1445 ne
rect 1840 -1450 1850 -1445
tri 1850 -1450 1855 -1445 sw
rect 1739 -1796 1754 -1568
rect 1840 -1606 1855 -1450
rect 1894 -1492 1922 -1436
tri 2014 -1454 2032 -1436 ne
rect 2032 -1456 2054 -1436
tri 2054 -1456 2074 -1436 sw
tri 2090 -1450 2108 -1432 ne
rect 1913 -1526 1922 -1492
rect 1956 -1465 1998 -1464
rect 1956 -1499 1961 -1465
rect 1991 -1499 1998 -1465
rect 1956 -1508 1998 -1499
rect 2032 -1465 2074 -1456
rect 2032 -1499 2039 -1465
rect 2069 -1499 2074 -1465
rect 2032 -1504 2074 -1499
rect 2108 -1492 2136 -1432
tri 2181 -1445 2203 -1423 se
rect 2203 -1430 2218 -1422
tri 2203 -1445 2218 -1430 nw
tri 2175 -1451 2181 -1445 se
rect 2181 -1451 2190 -1445
rect 1894 -1536 1922 -1526
tri 1922 -1536 1946 -1512 sw
rect 1894 -1568 1936 -1536
tri 1953 -1544 1954 -1543 sw
rect 1953 -1568 1954 -1544
tri 1956 -1545 1993 -1508 ne
rect 1993 -1536 1998 -1508
tri 1998 -1536 2024 -1510 sw
rect 2108 -1526 2117 -1492
rect 2108 -1536 2136 -1526
rect 1993 -1545 2077 -1536
tri 1993 -1564 2012 -1545 ne
rect 2012 -1564 2077 -1545
rect 1894 -1590 1954 -1568
rect 2076 -1568 2077 -1564
rect 2094 -1568 2136 -1536
rect 2076 -1590 2136 -1568
rect 1982 -1606 1999 -1592
rect 2031 -1606 2048 -1592
tri 1819 -1642 1841 -1620 se
rect 1841 -1627 1856 -1606
tri 1841 -1642 1856 -1627 nw
rect 2175 -1627 2190 -1451
tri 2190 -1458 2203 -1445 nw
rect 2276 -1526 2291 -1298
tri 1813 -1648 1819 -1642 se
rect 1819 -1648 1828 -1642
rect 1813 -1664 1828 -1648
tri 1828 -1655 1841 -1642 nw
rect 1982 -1650 1999 -1636
rect 2031 -1650 2048 -1636
tri 2175 -1642 2190 -1627 ne
tri 2190 -1642 2212 -1620 sw
rect 1813 -1700 1828 -1692
rect 1894 -1664 1954 -1650
rect 1909 -1674 1954 -1664
rect 1909 -1692 1937 -1674
tri 1813 -1715 1828 -1700 ne
tri 1828 -1715 1850 -1693 sw
rect 1894 -1702 1937 -1692
rect 1952 -1678 1954 -1674
rect 2076 -1664 2136 -1650
tri 2190 -1655 2203 -1642 ne
rect 2203 -1648 2212 -1642
tri 2212 -1648 2218 -1642 sw
rect 2076 -1674 2121 -1664
rect 1952 -1702 2026 -1678
rect 1894 -1706 2026 -1702
tri 2026 -1706 2054 -1678 sw
rect 2076 -1688 2078 -1674
tri 2076 -1690 2078 -1688 ne
rect 2090 -1692 2121 -1674
rect 2090 -1702 2136 -1692
rect 2203 -1663 2218 -1648
tri 1828 -1727 1840 -1715 ne
rect 1840 -1720 1850 -1715
tri 1850 -1720 1855 -1715 sw
rect 1739 -2066 1754 -1838
rect 1840 -1876 1855 -1720
rect 1894 -1762 1922 -1706
tri 2014 -1724 2032 -1706 ne
rect 2032 -1726 2054 -1706
tri 2054 -1726 2074 -1706 sw
tri 2090 -1720 2108 -1702 ne
rect 1913 -1796 1922 -1762
rect 1956 -1735 1998 -1734
rect 1956 -1769 1961 -1735
rect 1991 -1769 1998 -1735
rect 1956 -1778 1998 -1769
rect 2032 -1735 2074 -1726
rect 2032 -1769 2039 -1735
rect 2069 -1769 2074 -1735
rect 2032 -1774 2074 -1769
rect 2108 -1762 2136 -1702
tri 2181 -1715 2203 -1693 se
rect 2203 -1700 2218 -1692
tri 2203 -1715 2218 -1700 nw
tri 2175 -1721 2181 -1715 se
rect 2181 -1721 2190 -1715
rect 1894 -1806 1922 -1796
tri 1922 -1806 1946 -1782 sw
rect 1894 -1838 1936 -1806
tri 1953 -1814 1954 -1813 sw
rect 1953 -1838 1954 -1814
tri 1956 -1815 1993 -1778 ne
rect 1993 -1806 1998 -1778
tri 1998 -1806 2024 -1780 sw
rect 2108 -1796 2117 -1762
rect 2108 -1806 2136 -1796
rect 1993 -1815 2077 -1806
tri 1993 -1834 2012 -1815 ne
rect 2012 -1834 2077 -1815
rect 1894 -1860 1954 -1838
rect 2076 -1838 2077 -1834
rect 2094 -1838 2136 -1806
rect 2076 -1860 2136 -1838
rect 1982 -1876 1999 -1862
rect 2031 -1876 2048 -1862
tri 1819 -1912 1841 -1890 se
rect 1841 -1897 1856 -1876
tri 1841 -1912 1856 -1897 nw
rect 2175 -1897 2190 -1721
tri 2190 -1728 2203 -1715 nw
rect 2276 -1796 2291 -1568
tri 1813 -1918 1819 -1912 se
rect 1819 -1918 1828 -1912
rect 1813 -1934 1828 -1918
tri 1828 -1925 1841 -1912 nw
rect 1982 -1920 1999 -1906
rect 2031 -1920 2048 -1906
tri 2175 -1912 2190 -1897 ne
tri 2190 -1912 2212 -1890 sw
rect 1813 -1970 1828 -1962
rect 1894 -1934 1954 -1920
rect 1909 -1944 1954 -1934
rect 1909 -1962 1937 -1944
tri 1813 -1985 1828 -1970 ne
tri 1828 -1985 1850 -1963 sw
rect 1894 -1972 1937 -1962
rect 1952 -1948 1954 -1944
rect 2076 -1934 2136 -1920
tri 2190 -1925 2203 -1912 ne
rect 2203 -1918 2212 -1912
tri 2212 -1918 2218 -1912 sw
rect 2076 -1944 2121 -1934
rect 1952 -1972 2026 -1948
rect 1894 -1976 2026 -1972
tri 2026 -1976 2054 -1948 sw
rect 2076 -1958 2078 -1944
tri 2076 -1960 2078 -1958 ne
rect 2090 -1962 2121 -1944
rect 2090 -1972 2136 -1962
rect 2203 -1933 2218 -1918
tri 1828 -1997 1840 -1985 ne
rect 1840 -1990 1850 -1985
tri 1850 -1990 1855 -1985 sw
rect 1739 -2146 1754 -2108
rect 1840 -2146 1855 -1990
rect 1894 -2032 1922 -1976
tri 2014 -1994 2032 -1976 ne
rect 2032 -1996 2054 -1976
tri 2054 -1996 2074 -1976 sw
tri 2090 -1990 2108 -1972 ne
rect 1913 -2066 1922 -2032
rect 1956 -2005 1998 -2004
rect 1956 -2039 1961 -2005
rect 1991 -2039 1998 -2005
rect 1956 -2048 1998 -2039
rect 2032 -2005 2074 -1996
rect 2032 -2039 2039 -2005
rect 2069 -2039 2074 -2005
rect 2032 -2044 2074 -2039
rect 2108 -2032 2136 -1972
tri 2181 -1985 2203 -1963 se
rect 2203 -1970 2218 -1962
tri 2203 -1985 2218 -1970 nw
tri 2175 -1991 2181 -1985 se
rect 2181 -1991 2190 -1985
rect 1894 -2076 1922 -2066
tri 1922 -2076 1946 -2052 sw
rect 1894 -2108 1936 -2076
tri 1953 -2084 1954 -2083 sw
rect 1953 -2108 1954 -2084
tri 1956 -2085 1993 -2048 ne
rect 1993 -2076 1998 -2048
tri 1998 -2076 2024 -2050 sw
rect 2108 -2066 2117 -2032
rect 2108 -2076 2136 -2066
rect 1993 -2085 2077 -2076
tri 1993 -2104 2012 -2085 ne
rect 2012 -2104 2077 -2085
rect 1894 -2130 1954 -2108
rect 2076 -2108 2077 -2104
rect 2094 -2108 2136 -2076
rect 2076 -2130 2136 -2108
rect 1982 -2146 1999 -2132
rect 2031 -2146 2048 -2132
rect 2175 -2146 2190 -1991
tri 2190 -1998 2203 -1985 nw
rect 2276 -2066 2291 -1838
rect 2276 -2146 2291 -2108
rect 2319 1984 2334 2174
tri 2399 2138 2421 2160 se
rect 2421 2153 2436 2174
tri 2421 2138 2436 2153 nw
rect 2755 2153 2770 2174
tri 2393 2132 2399 2138 se
rect 2399 2132 2408 2138
rect 2393 2116 2408 2132
tri 2408 2125 2421 2138 nw
rect 2562 2130 2579 2144
rect 2611 2130 2628 2144
tri 2755 2138 2770 2153 ne
tri 2770 2138 2792 2160 sw
rect 2393 2080 2408 2088
rect 2474 2116 2534 2130
rect 2489 2106 2534 2116
rect 2489 2088 2517 2106
tri 2393 2065 2408 2080 ne
tri 2408 2065 2430 2087 sw
rect 2474 2078 2517 2088
rect 2532 2102 2534 2106
rect 2656 2116 2716 2130
tri 2770 2125 2783 2138 ne
rect 2783 2132 2792 2138
tri 2792 2132 2798 2138 sw
rect 2656 2106 2701 2116
rect 2532 2078 2606 2102
rect 2474 2074 2606 2078
tri 2606 2074 2634 2102 sw
rect 2656 2092 2658 2106
tri 2656 2090 2658 2092 ne
rect 2670 2088 2701 2106
rect 2670 2078 2716 2088
rect 2783 2117 2798 2132
tri 2408 2053 2420 2065 ne
rect 2420 2060 2430 2065
tri 2430 2060 2435 2065 sw
rect 2319 1714 2334 1942
rect 2420 1904 2435 2060
rect 2474 2018 2502 2074
tri 2594 2056 2612 2074 ne
rect 2612 2054 2634 2074
tri 2634 2054 2654 2074 sw
tri 2670 2060 2688 2078 ne
rect 2493 1984 2502 2018
rect 2536 2045 2578 2046
rect 2536 2011 2541 2045
rect 2571 2011 2578 2045
rect 2536 2002 2578 2011
rect 2612 2045 2654 2054
rect 2612 2011 2619 2045
rect 2649 2011 2654 2045
rect 2612 2006 2654 2011
rect 2688 2018 2716 2078
tri 2761 2065 2783 2087 se
rect 2783 2080 2798 2088
tri 2783 2065 2798 2080 nw
tri 2755 2059 2761 2065 se
rect 2761 2059 2770 2065
rect 2474 1974 2502 1984
tri 2502 1974 2526 1998 sw
rect 2474 1942 2516 1974
tri 2533 1966 2534 1967 sw
rect 2533 1942 2534 1966
tri 2536 1965 2573 2002 ne
rect 2573 1974 2578 2002
tri 2578 1974 2604 2000 sw
rect 2688 1984 2697 2018
rect 2688 1974 2716 1984
rect 2573 1965 2657 1974
tri 2573 1946 2592 1965 ne
rect 2592 1946 2657 1965
rect 2474 1920 2534 1942
rect 2656 1942 2657 1946
rect 2674 1942 2716 1974
rect 2656 1920 2716 1942
rect 2562 1904 2579 1918
rect 2611 1904 2628 1918
tri 2399 1868 2421 1890 se
rect 2421 1883 2436 1904
tri 2421 1868 2436 1883 nw
rect 2755 1883 2770 2059
tri 2770 2052 2783 2065 nw
rect 2856 1984 2871 2174
tri 2393 1862 2399 1868 se
rect 2399 1862 2408 1868
rect 2393 1846 2408 1862
tri 2408 1855 2421 1868 nw
rect 2562 1860 2579 1874
rect 2611 1860 2628 1874
tri 2755 1868 2770 1883 ne
tri 2770 1868 2792 1890 sw
rect 2393 1810 2408 1818
rect 2474 1846 2534 1860
rect 2489 1836 2534 1846
rect 2489 1818 2517 1836
tri 2393 1795 2408 1810 ne
tri 2408 1795 2430 1817 sw
rect 2474 1808 2517 1818
rect 2532 1832 2534 1836
rect 2656 1846 2716 1860
tri 2770 1855 2783 1868 ne
rect 2783 1862 2792 1868
tri 2792 1862 2798 1868 sw
rect 2656 1836 2701 1846
rect 2532 1808 2606 1832
rect 2474 1804 2606 1808
tri 2606 1804 2634 1832 sw
rect 2656 1822 2658 1836
tri 2656 1820 2658 1822 ne
rect 2670 1818 2701 1836
rect 2670 1808 2716 1818
rect 2783 1847 2798 1862
tri 2408 1783 2420 1795 ne
rect 2420 1790 2430 1795
tri 2430 1790 2435 1795 sw
rect 2319 1444 2334 1672
rect 2420 1634 2435 1790
rect 2474 1748 2502 1804
tri 2594 1786 2612 1804 ne
rect 2612 1784 2634 1804
tri 2634 1784 2654 1804 sw
tri 2670 1790 2688 1808 ne
rect 2493 1714 2502 1748
rect 2536 1775 2578 1776
rect 2536 1741 2541 1775
rect 2571 1741 2578 1775
rect 2536 1732 2578 1741
rect 2612 1775 2654 1784
rect 2612 1741 2619 1775
rect 2649 1741 2654 1775
rect 2612 1736 2654 1741
rect 2688 1748 2716 1808
tri 2761 1795 2783 1817 se
rect 2783 1810 2798 1818
tri 2783 1795 2798 1810 nw
tri 2755 1789 2761 1795 se
rect 2761 1789 2770 1795
rect 2474 1704 2502 1714
tri 2502 1704 2526 1728 sw
rect 2474 1672 2516 1704
tri 2533 1696 2534 1697 sw
rect 2533 1672 2534 1696
tri 2536 1695 2573 1732 ne
rect 2573 1704 2578 1732
tri 2578 1704 2604 1730 sw
rect 2688 1714 2697 1748
rect 2688 1704 2716 1714
rect 2573 1695 2657 1704
tri 2573 1676 2592 1695 ne
rect 2592 1676 2657 1695
rect 2474 1650 2534 1672
rect 2656 1672 2657 1676
rect 2674 1672 2716 1704
rect 2656 1650 2716 1672
rect 2562 1634 2579 1648
rect 2611 1634 2628 1648
tri 2399 1598 2421 1620 se
rect 2421 1613 2436 1634
tri 2421 1598 2436 1613 nw
rect 2755 1613 2770 1789
tri 2770 1782 2783 1795 nw
rect 2856 1714 2871 1942
tri 2393 1592 2399 1598 se
rect 2399 1592 2408 1598
rect 2393 1576 2408 1592
tri 2408 1585 2421 1598 nw
rect 2562 1590 2579 1604
rect 2611 1590 2628 1604
tri 2755 1598 2770 1613 ne
tri 2770 1598 2792 1620 sw
rect 2393 1540 2408 1548
rect 2474 1576 2534 1590
rect 2489 1566 2534 1576
rect 2489 1548 2517 1566
tri 2393 1525 2408 1540 ne
tri 2408 1525 2430 1547 sw
rect 2474 1538 2517 1548
rect 2532 1562 2534 1566
rect 2656 1576 2716 1590
tri 2770 1585 2783 1598 ne
rect 2783 1592 2792 1598
tri 2792 1592 2798 1598 sw
rect 2656 1566 2701 1576
rect 2532 1538 2606 1562
rect 2474 1534 2606 1538
tri 2606 1534 2634 1562 sw
rect 2656 1552 2658 1566
tri 2656 1550 2658 1552 ne
rect 2670 1548 2701 1566
rect 2670 1538 2716 1548
rect 2783 1577 2798 1592
tri 2408 1513 2420 1525 ne
rect 2420 1520 2430 1525
tri 2430 1520 2435 1525 sw
rect 2319 1174 2334 1402
rect 2420 1364 2435 1520
rect 2474 1478 2502 1534
tri 2594 1516 2612 1534 ne
rect 2612 1514 2634 1534
tri 2634 1514 2654 1534 sw
tri 2670 1520 2688 1538 ne
rect 2493 1444 2502 1478
rect 2536 1505 2578 1506
rect 2536 1471 2541 1505
rect 2571 1471 2578 1505
rect 2536 1462 2578 1471
rect 2612 1505 2654 1514
rect 2612 1471 2619 1505
rect 2649 1471 2654 1505
rect 2612 1466 2654 1471
rect 2688 1478 2716 1538
tri 2761 1525 2783 1547 se
rect 2783 1540 2798 1548
tri 2783 1525 2798 1540 nw
tri 2755 1519 2761 1525 se
rect 2761 1519 2770 1525
rect 2474 1434 2502 1444
tri 2502 1434 2526 1458 sw
rect 2474 1402 2516 1434
tri 2533 1426 2534 1427 sw
rect 2533 1402 2534 1426
tri 2536 1425 2573 1462 ne
rect 2573 1434 2578 1462
tri 2578 1434 2604 1460 sw
rect 2688 1444 2697 1478
rect 2688 1434 2716 1444
rect 2573 1425 2657 1434
tri 2573 1406 2592 1425 ne
rect 2592 1406 2657 1425
rect 2474 1380 2534 1402
rect 2656 1402 2657 1406
rect 2674 1402 2716 1434
rect 2656 1380 2716 1402
rect 2562 1364 2579 1378
rect 2611 1364 2628 1378
tri 2399 1328 2421 1350 se
rect 2421 1343 2436 1364
tri 2421 1328 2436 1343 nw
rect 2755 1343 2770 1519
tri 2770 1512 2783 1525 nw
rect 2856 1444 2871 1672
tri 2393 1322 2399 1328 se
rect 2399 1322 2408 1328
rect 2393 1306 2408 1322
tri 2408 1315 2421 1328 nw
rect 2562 1320 2579 1334
rect 2611 1320 2628 1334
tri 2755 1328 2770 1343 ne
tri 2770 1328 2792 1350 sw
rect 2393 1270 2408 1278
rect 2474 1306 2534 1320
rect 2489 1296 2534 1306
rect 2489 1278 2517 1296
tri 2393 1255 2408 1270 ne
tri 2408 1255 2430 1277 sw
rect 2474 1268 2517 1278
rect 2532 1292 2534 1296
rect 2656 1306 2716 1320
tri 2770 1315 2783 1328 ne
rect 2783 1322 2792 1328
tri 2792 1322 2798 1328 sw
rect 2656 1296 2701 1306
rect 2532 1268 2606 1292
rect 2474 1264 2606 1268
tri 2606 1264 2634 1292 sw
rect 2656 1282 2658 1296
tri 2656 1280 2658 1282 ne
rect 2670 1278 2701 1296
rect 2670 1268 2716 1278
rect 2783 1307 2798 1322
tri 2408 1243 2420 1255 ne
rect 2420 1250 2430 1255
tri 2430 1250 2435 1255 sw
rect 2319 904 2334 1132
rect 2420 1094 2435 1250
rect 2474 1208 2502 1264
tri 2594 1246 2612 1264 ne
rect 2612 1244 2634 1264
tri 2634 1244 2654 1264 sw
tri 2670 1250 2688 1268 ne
rect 2493 1174 2502 1208
rect 2536 1235 2578 1236
rect 2536 1201 2541 1235
rect 2571 1201 2578 1235
rect 2536 1192 2578 1201
rect 2612 1235 2654 1244
rect 2612 1201 2619 1235
rect 2649 1201 2654 1235
rect 2612 1196 2654 1201
rect 2688 1208 2716 1268
tri 2761 1255 2783 1277 se
rect 2783 1270 2798 1278
tri 2783 1255 2798 1270 nw
tri 2755 1249 2761 1255 se
rect 2761 1249 2770 1255
rect 2474 1164 2502 1174
tri 2502 1164 2526 1188 sw
rect 2474 1132 2516 1164
tri 2533 1156 2534 1157 sw
rect 2533 1132 2534 1156
tri 2536 1155 2573 1192 ne
rect 2573 1164 2578 1192
tri 2578 1164 2604 1190 sw
rect 2688 1174 2697 1208
rect 2688 1164 2716 1174
rect 2573 1155 2657 1164
tri 2573 1136 2592 1155 ne
rect 2592 1136 2657 1155
rect 2474 1110 2534 1132
rect 2656 1132 2657 1136
rect 2674 1132 2716 1164
rect 2656 1110 2716 1132
rect 2562 1094 2579 1108
rect 2611 1094 2628 1108
tri 2399 1058 2421 1080 se
rect 2421 1073 2436 1094
tri 2421 1058 2436 1073 nw
rect 2755 1073 2770 1249
tri 2770 1242 2783 1255 nw
rect 2856 1174 2871 1402
tri 2393 1052 2399 1058 se
rect 2399 1052 2408 1058
rect 2393 1036 2408 1052
tri 2408 1045 2421 1058 nw
rect 2562 1050 2579 1064
rect 2611 1050 2628 1064
tri 2755 1058 2770 1073 ne
tri 2770 1058 2792 1080 sw
rect 2393 1000 2408 1008
rect 2474 1036 2534 1050
rect 2489 1026 2534 1036
rect 2489 1008 2517 1026
tri 2393 985 2408 1000 ne
tri 2408 985 2430 1007 sw
rect 2474 998 2517 1008
rect 2532 1022 2534 1026
rect 2656 1036 2716 1050
tri 2770 1045 2783 1058 ne
rect 2783 1052 2792 1058
tri 2792 1052 2798 1058 sw
rect 2656 1026 2701 1036
rect 2532 998 2606 1022
rect 2474 994 2606 998
tri 2606 994 2634 1022 sw
rect 2656 1012 2658 1026
tri 2656 1010 2658 1012 ne
rect 2670 1008 2701 1026
rect 2670 998 2716 1008
rect 2783 1037 2798 1052
tri 2408 973 2420 985 ne
rect 2420 980 2430 985
tri 2430 980 2435 985 sw
rect 2319 634 2334 862
rect 2420 824 2435 980
rect 2474 938 2502 994
tri 2594 976 2612 994 ne
rect 2612 974 2634 994
tri 2634 974 2654 994 sw
tri 2670 980 2688 998 ne
rect 2493 904 2502 938
rect 2536 965 2578 966
rect 2536 931 2541 965
rect 2571 931 2578 965
rect 2536 922 2578 931
rect 2612 965 2654 974
rect 2612 931 2619 965
rect 2649 931 2654 965
rect 2612 926 2654 931
rect 2688 938 2716 998
tri 2761 985 2783 1007 se
rect 2783 1000 2798 1008
tri 2783 985 2798 1000 nw
tri 2755 979 2761 985 se
rect 2761 979 2770 985
rect 2474 894 2502 904
tri 2502 894 2526 918 sw
rect 2474 862 2516 894
tri 2533 886 2534 887 sw
rect 2533 862 2534 886
tri 2536 885 2573 922 ne
rect 2573 894 2578 922
tri 2578 894 2604 920 sw
rect 2688 904 2697 938
rect 2688 894 2716 904
rect 2573 885 2657 894
tri 2573 866 2592 885 ne
rect 2592 866 2657 885
rect 2474 840 2534 862
rect 2656 862 2657 866
rect 2674 862 2716 894
rect 2656 840 2716 862
rect 2562 824 2579 838
rect 2611 824 2628 838
tri 2399 788 2421 810 se
rect 2421 803 2436 824
tri 2421 788 2436 803 nw
rect 2755 803 2770 979
tri 2770 972 2783 985 nw
rect 2856 904 2871 1132
tri 2393 782 2399 788 se
rect 2399 782 2408 788
rect 2393 766 2408 782
tri 2408 775 2421 788 nw
rect 2562 780 2579 794
rect 2611 780 2628 794
tri 2755 788 2770 803 ne
tri 2770 788 2792 810 sw
rect 2393 730 2408 738
rect 2474 766 2534 780
rect 2489 756 2534 766
rect 2489 738 2517 756
tri 2393 715 2408 730 ne
tri 2408 715 2430 737 sw
rect 2474 728 2517 738
rect 2532 752 2534 756
rect 2656 766 2716 780
tri 2770 775 2783 788 ne
rect 2783 782 2792 788
tri 2792 782 2798 788 sw
rect 2656 756 2701 766
rect 2532 728 2606 752
rect 2474 724 2606 728
tri 2606 724 2634 752 sw
rect 2656 742 2658 756
tri 2656 740 2658 742 ne
rect 2670 738 2701 756
rect 2670 728 2716 738
rect 2783 767 2798 782
tri 2408 703 2420 715 ne
rect 2420 710 2430 715
tri 2430 710 2435 715 sw
rect 2319 364 2334 592
rect 2420 554 2435 710
rect 2474 668 2502 724
tri 2594 706 2612 724 ne
rect 2612 704 2634 724
tri 2634 704 2654 724 sw
tri 2670 710 2688 728 ne
rect 2493 634 2502 668
rect 2536 695 2578 696
rect 2536 661 2541 695
rect 2571 661 2578 695
rect 2536 652 2578 661
rect 2612 695 2654 704
rect 2612 661 2619 695
rect 2649 661 2654 695
rect 2612 656 2654 661
rect 2688 668 2716 728
tri 2761 715 2783 737 se
rect 2783 730 2798 738
tri 2783 715 2798 730 nw
tri 2755 709 2761 715 se
rect 2761 709 2770 715
rect 2474 624 2502 634
tri 2502 624 2526 648 sw
rect 2474 592 2516 624
tri 2533 616 2534 617 sw
rect 2533 592 2534 616
tri 2536 615 2573 652 ne
rect 2573 624 2578 652
tri 2578 624 2604 650 sw
rect 2688 634 2697 668
rect 2688 624 2716 634
rect 2573 615 2657 624
tri 2573 596 2592 615 ne
rect 2592 596 2657 615
rect 2474 570 2534 592
rect 2656 592 2657 596
rect 2674 592 2716 624
rect 2656 570 2716 592
rect 2562 554 2579 568
rect 2611 554 2628 568
tri 2399 518 2421 540 se
rect 2421 533 2436 554
tri 2421 518 2436 533 nw
rect 2755 533 2770 709
tri 2770 702 2783 715 nw
rect 2856 634 2871 862
tri 2393 512 2399 518 se
rect 2399 512 2408 518
rect 2393 496 2408 512
tri 2408 505 2421 518 nw
rect 2562 510 2579 524
rect 2611 510 2628 524
tri 2755 518 2770 533 ne
tri 2770 518 2792 540 sw
rect 2393 460 2408 468
rect 2474 496 2534 510
rect 2489 486 2534 496
rect 2489 468 2517 486
tri 2393 445 2408 460 ne
tri 2408 445 2430 467 sw
rect 2474 458 2517 468
rect 2532 482 2534 486
rect 2656 496 2716 510
tri 2770 505 2783 518 ne
rect 2783 512 2792 518
tri 2792 512 2798 518 sw
rect 2656 486 2701 496
rect 2532 458 2606 482
rect 2474 454 2606 458
tri 2606 454 2634 482 sw
rect 2656 472 2658 486
tri 2656 470 2658 472 ne
rect 2670 468 2701 486
rect 2670 458 2716 468
rect 2783 497 2798 512
tri 2408 433 2420 445 ne
rect 2420 440 2430 445
tri 2430 440 2435 445 sw
rect 2319 94 2334 322
rect 2420 284 2435 440
rect 2474 398 2502 454
tri 2594 436 2612 454 ne
rect 2612 434 2634 454
tri 2634 434 2654 454 sw
tri 2670 440 2688 458 ne
rect 2493 364 2502 398
rect 2536 425 2578 426
rect 2536 391 2541 425
rect 2571 391 2578 425
rect 2536 382 2578 391
rect 2612 425 2654 434
rect 2612 391 2619 425
rect 2649 391 2654 425
rect 2612 386 2654 391
rect 2688 398 2716 458
tri 2761 445 2783 467 se
rect 2783 460 2798 468
tri 2783 445 2798 460 nw
tri 2755 439 2761 445 se
rect 2761 439 2770 445
rect 2474 354 2502 364
tri 2502 354 2526 378 sw
rect 2474 322 2516 354
tri 2533 346 2534 347 sw
rect 2533 322 2534 346
tri 2536 345 2573 382 ne
rect 2573 354 2578 382
tri 2578 354 2604 380 sw
rect 2688 364 2697 398
rect 2688 354 2716 364
rect 2573 345 2657 354
tri 2573 326 2592 345 ne
rect 2592 326 2657 345
rect 2474 300 2534 322
rect 2656 322 2657 326
rect 2674 322 2716 354
rect 2656 300 2716 322
rect 2562 284 2579 298
rect 2611 284 2628 298
tri 2399 248 2421 270 se
rect 2421 263 2436 284
tri 2421 248 2436 263 nw
rect 2755 263 2770 439
tri 2770 432 2783 445 nw
rect 2856 364 2871 592
tri 2393 242 2399 248 se
rect 2399 242 2408 248
rect 2393 226 2408 242
tri 2408 235 2421 248 nw
rect 2562 240 2579 254
rect 2611 240 2628 254
tri 2755 248 2770 263 ne
tri 2770 248 2792 270 sw
rect 2393 190 2408 198
rect 2474 226 2534 240
rect 2489 216 2534 226
rect 2489 198 2517 216
tri 2393 175 2408 190 ne
tri 2408 175 2430 197 sw
rect 2474 188 2517 198
rect 2532 212 2534 216
rect 2656 226 2716 240
tri 2770 235 2783 248 ne
rect 2783 242 2792 248
tri 2792 242 2798 248 sw
rect 2656 216 2701 226
rect 2532 188 2606 212
rect 2474 184 2606 188
tri 2606 184 2634 212 sw
rect 2656 202 2658 216
tri 2656 200 2658 202 ne
rect 2670 198 2701 216
rect 2670 188 2716 198
rect 2783 227 2798 242
tri 2408 163 2420 175 ne
rect 2420 170 2430 175
tri 2430 170 2435 175 sw
rect 2319 -176 2334 52
rect 2420 14 2435 170
rect 2474 128 2502 184
tri 2594 166 2612 184 ne
rect 2612 164 2634 184
tri 2634 164 2654 184 sw
tri 2670 170 2688 188 ne
rect 2493 94 2502 128
rect 2536 155 2578 156
rect 2536 121 2541 155
rect 2571 121 2578 155
rect 2536 112 2578 121
rect 2612 155 2654 164
rect 2612 121 2619 155
rect 2649 121 2654 155
rect 2612 116 2654 121
rect 2688 128 2716 188
tri 2761 175 2783 197 se
rect 2783 190 2798 198
tri 2783 175 2798 190 nw
tri 2755 169 2761 175 se
rect 2761 169 2770 175
rect 2474 84 2502 94
tri 2502 84 2526 108 sw
rect 2474 52 2516 84
tri 2533 76 2534 77 sw
rect 2533 52 2534 76
tri 2536 75 2573 112 ne
rect 2573 84 2578 112
tri 2578 84 2604 110 sw
rect 2688 94 2697 128
rect 2688 84 2716 94
rect 2573 75 2657 84
tri 2573 56 2592 75 ne
rect 2592 56 2657 75
rect 2474 30 2534 52
rect 2656 52 2657 56
rect 2674 52 2716 84
rect 2656 30 2716 52
rect 2562 14 2579 28
rect 2611 14 2628 28
tri 2399 -22 2421 0 se
rect 2421 -7 2436 14
tri 2421 -22 2436 -7 nw
rect 2755 -7 2770 169
tri 2770 162 2783 175 nw
rect 2856 94 2871 322
tri 2393 -28 2399 -22 se
rect 2399 -28 2408 -22
rect 2393 -44 2408 -28
tri 2408 -35 2421 -22 nw
rect 2562 -30 2579 -16
rect 2611 -30 2628 -16
tri 2755 -22 2770 -7 ne
tri 2770 -22 2792 0 sw
rect 2393 -80 2408 -72
rect 2474 -44 2534 -30
rect 2489 -54 2534 -44
rect 2489 -72 2517 -54
tri 2393 -95 2408 -80 ne
tri 2408 -95 2430 -73 sw
rect 2474 -82 2517 -72
rect 2532 -58 2534 -54
rect 2656 -44 2716 -30
tri 2770 -35 2783 -22 ne
rect 2783 -28 2792 -22
tri 2792 -28 2798 -22 sw
rect 2656 -54 2701 -44
rect 2532 -82 2606 -58
rect 2474 -86 2606 -82
tri 2606 -86 2634 -58 sw
rect 2656 -68 2658 -54
tri 2656 -70 2658 -68 ne
rect 2670 -72 2701 -54
rect 2670 -82 2716 -72
rect 2783 -43 2798 -28
tri 2408 -107 2420 -95 ne
rect 2420 -100 2430 -95
tri 2430 -100 2435 -95 sw
rect 2319 -446 2334 -218
rect 2420 -256 2435 -100
rect 2474 -142 2502 -86
tri 2594 -104 2612 -86 ne
rect 2612 -106 2634 -86
tri 2634 -106 2654 -86 sw
tri 2670 -100 2688 -82 ne
rect 2493 -176 2502 -142
rect 2536 -115 2578 -114
rect 2536 -149 2541 -115
rect 2571 -149 2578 -115
rect 2536 -158 2578 -149
rect 2612 -115 2654 -106
rect 2612 -149 2619 -115
rect 2649 -149 2654 -115
rect 2612 -154 2654 -149
rect 2688 -142 2716 -82
tri 2761 -95 2783 -73 se
rect 2783 -80 2798 -72
tri 2783 -95 2798 -80 nw
tri 2755 -101 2761 -95 se
rect 2761 -101 2770 -95
rect 2474 -186 2502 -176
tri 2502 -186 2526 -162 sw
rect 2474 -218 2516 -186
tri 2533 -194 2534 -193 sw
rect 2533 -218 2534 -194
tri 2536 -195 2573 -158 ne
rect 2573 -186 2578 -158
tri 2578 -186 2604 -160 sw
rect 2688 -176 2697 -142
rect 2688 -186 2716 -176
rect 2573 -195 2657 -186
tri 2573 -214 2592 -195 ne
rect 2592 -214 2657 -195
rect 2474 -240 2534 -218
rect 2656 -218 2657 -214
rect 2674 -218 2716 -186
rect 2656 -240 2716 -218
rect 2562 -256 2579 -242
rect 2611 -256 2628 -242
tri 2399 -292 2421 -270 se
rect 2421 -277 2436 -256
tri 2421 -292 2436 -277 nw
rect 2755 -277 2770 -101
tri 2770 -108 2783 -95 nw
rect 2856 -176 2871 52
tri 2393 -298 2399 -292 se
rect 2399 -298 2408 -292
rect 2393 -314 2408 -298
tri 2408 -305 2421 -292 nw
rect 2562 -300 2579 -286
rect 2611 -300 2628 -286
tri 2755 -292 2770 -277 ne
tri 2770 -292 2792 -270 sw
rect 2393 -350 2408 -342
rect 2474 -314 2534 -300
rect 2489 -324 2534 -314
rect 2489 -342 2517 -324
tri 2393 -365 2408 -350 ne
tri 2408 -365 2430 -343 sw
rect 2474 -352 2517 -342
rect 2532 -328 2534 -324
rect 2656 -314 2716 -300
tri 2770 -305 2783 -292 ne
rect 2783 -298 2792 -292
tri 2792 -298 2798 -292 sw
rect 2656 -324 2701 -314
rect 2532 -352 2606 -328
rect 2474 -356 2606 -352
tri 2606 -356 2634 -328 sw
rect 2656 -338 2658 -324
tri 2656 -340 2658 -338 ne
rect 2670 -342 2701 -324
rect 2670 -352 2716 -342
rect 2783 -313 2798 -298
tri 2408 -377 2420 -365 ne
rect 2420 -370 2430 -365
tri 2430 -370 2435 -365 sw
rect 2319 -716 2334 -488
rect 2420 -526 2435 -370
rect 2474 -412 2502 -356
tri 2594 -374 2612 -356 ne
rect 2612 -376 2634 -356
tri 2634 -376 2654 -356 sw
tri 2670 -370 2688 -352 ne
rect 2493 -446 2502 -412
rect 2536 -385 2578 -384
rect 2536 -419 2541 -385
rect 2571 -419 2578 -385
rect 2536 -428 2578 -419
rect 2612 -385 2654 -376
rect 2612 -419 2619 -385
rect 2649 -419 2654 -385
rect 2612 -424 2654 -419
rect 2688 -412 2716 -352
tri 2761 -365 2783 -343 se
rect 2783 -350 2798 -342
tri 2783 -365 2798 -350 nw
tri 2755 -371 2761 -365 se
rect 2761 -371 2770 -365
rect 2474 -456 2502 -446
tri 2502 -456 2526 -432 sw
rect 2474 -488 2516 -456
tri 2533 -464 2534 -463 sw
rect 2533 -488 2534 -464
tri 2536 -465 2573 -428 ne
rect 2573 -456 2578 -428
tri 2578 -456 2604 -430 sw
rect 2688 -446 2697 -412
rect 2688 -456 2716 -446
rect 2573 -465 2657 -456
tri 2573 -484 2592 -465 ne
rect 2592 -484 2657 -465
rect 2474 -510 2534 -488
rect 2656 -488 2657 -484
rect 2674 -488 2716 -456
rect 2656 -510 2716 -488
rect 2562 -526 2579 -512
rect 2611 -526 2628 -512
tri 2399 -562 2421 -540 se
rect 2421 -547 2436 -526
tri 2421 -562 2436 -547 nw
rect 2755 -547 2770 -371
tri 2770 -378 2783 -365 nw
rect 2856 -446 2871 -218
tri 2393 -568 2399 -562 se
rect 2399 -568 2408 -562
rect 2393 -584 2408 -568
tri 2408 -575 2421 -562 nw
rect 2562 -570 2579 -556
rect 2611 -570 2628 -556
tri 2755 -562 2770 -547 ne
tri 2770 -562 2792 -540 sw
rect 2393 -620 2408 -612
rect 2474 -584 2534 -570
rect 2489 -594 2534 -584
rect 2489 -612 2517 -594
tri 2393 -635 2408 -620 ne
tri 2408 -635 2430 -613 sw
rect 2474 -622 2517 -612
rect 2532 -598 2534 -594
rect 2656 -584 2716 -570
tri 2770 -575 2783 -562 ne
rect 2783 -568 2792 -562
tri 2792 -568 2798 -562 sw
rect 2656 -594 2701 -584
rect 2532 -622 2606 -598
rect 2474 -626 2606 -622
tri 2606 -626 2634 -598 sw
rect 2656 -608 2658 -594
tri 2656 -610 2658 -608 ne
rect 2670 -612 2701 -594
rect 2670 -622 2716 -612
rect 2783 -583 2798 -568
tri 2408 -647 2420 -635 ne
rect 2420 -640 2430 -635
tri 2430 -640 2435 -635 sw
rect 2319 -986 2334 -758
rect 2420 -796 2435 -640
rect 2474 -682 2502 -626
tri 2594 -644 2612 -626 ne
rect 2612 -646 2634 -626
tri 2634 -646 2654 -626 sw
tri 2670 -640 2688 -622 ne
rect 2493 -716 2502 -682
rect 2536 -655 2578 -654
rect 2536 -689 2541 -655
rect 2571 -689 2578 -655
rect 2536 -698 2578 -689
rect 2612 -655 2654 -646
rect 2612 -689 2619 -655
rect 2649 -689 2654 -655
rect 2612 -694 2654 -689
rect 2688 -682 2716 -622
tri 2761 -635 2783 -613 se
rect 2783 -620 2798 -612
tri 2783 -635 2798 -620 nw
tri 2755 -641 2761 -635 se
rect 2761 -641 2770 -635
rect 2474 -726 2502 -716
tri 2502 -726 2526 -702 sw
rect 2474 -758 2516 -726
tri 2533 -734 2534 -733 sw
rect 2533 -758 2534 -734
tri 2536 -735 2573 -698 ne
rect 2573 -726 2578 -698
tri 2578 -726 2604 -700 sw
rect 2688 -716 2697 -682
rect 2688 -726 2716 -716
rect 2573 -735 2657 -726
tri 2573 -754 2592 -735 ne
rect 2592 -754 2657 -735
rect 2474 -780 2534 -758
rect 2656 -758 2657 -754
rect 2674 -758 2716 -726
rect 2656 -780 2716 -758
rect 2562 -796 2579 -782
rect 2611 -796 2628 -782
tri 2399 -832 2421 -810 se
rect 2421 -817 2436 -796
tri 2421 -832 2436 -817 nw
rect 2755 -817 2770 -641
tri 2770 -648 2783 -635 nw
rect 2856 -716 2871 -488
tri 2393 -838 2399 -832 se
rect 2399 -838 2408 -832
rect 2393 -854 2408 -838
tri 2408 -845 2421 -832 nw
rect 2562 -840 2579 -826
rect 2611 -840 2628 -826
tri 2755 -832 2770 -817 ne
tri 2770 -832 2792 -810 sw
rect 2393 -890 2408 -882
rect 2474 -854 2534 -840
rect 2489 -864 2534 -854
rect 2489 -882 2517 -864
tri 2393 -905 2408 -890 ne
tri 2408 -905 2430 -883 sw
rect 2474 -892 2517 -882
rect 2532 -868 2534 -864
rect 2656 -854 2716 -840
tri 2770 -845 2783 -832 ne
rect 2783 -838 2792 -832
tri 2792 -838 2798 -832 sw
rect 2656 -864 2701 -854
rect 2532 -892 2606 -868
rect 2474 -896 2606 -892
tri 2606 -896 2634 -868 sw
rect 2656 -878 2658 -864
tri 2656 -880 2658 -878 ne
rect 2670 -882 2701 -864
rect 2670 -892 2716 -882
rect 2783 -853 2798 -838
tri 2408 -917 2420 -905 ne
rect 2420 -910 2430 -905
tri 2430 -910 2435 -905 sw
rect 2319 -1256 2334 -1028
rect 2420 -1066 2435 -910
rect 2474 -952 2502 -896
tri 2594 -914 2612 -896 ne
rect 2612 -916 2634 -896
tri 2634 -916 2654 -896 sw
tri 2670 -910 2688 -892 ne
rect 2493 -986 2502 -952
rect 2536 -925 2578 -924
rect 2536 -959 2541 -925
rect 2571 -959 2578 -925
rect 2536 -968 2578 -959
rect 2612 -925 2654 -916
rect 2612 -959 2619 -925
rect 2649 -959 2654 -925
rect 2612 -964 2654 -959
rect 2688 -952 2716 -892
tri 2761 -905 2783 -883 se
rect 2783 -890 2798 -882
tri 2783 -905 2798 -890 nw
tri 2755 -911 2761 -905 se
rect 2761 -911 2770 -905
rect 2474 -996 2502 -986
tri 2502 -996 2526 -972 sw
rect 2474 -1028 2516 -996
tri 2533 -1004 2534 -1003 sw
rect 2533 -1028 2534 -1004
tri 2536 -1005 2573 -968 ne
rect 2573 -996 2578 -968
tri 2578 -996 2604 -970 sw
rect 2688 -986 2697 -952
rect 2688 -996 2716 -986
rect 2573 -1005 2657 -996
tri 2573 -1024 2592 -1005 ne
rect 2592 -1024 2657 -1005
rect 2474 -1050 2534 -1028
rect 2656 -1028 2657 -1024
rect 2674 -1028 2716 -996
rect 2656 -1050 2716 -1028
rect 2562 -1066 2579 -1052
rect 2611 -1066 2628 -1052
tri 2399 -1102 2421 -1080 se
rect 2421 -1087 2436 -1066
tri 2421 -1102 2436 -1087 nw
rect 2755 -1087 2770 -911
tri 2770 -918 2783 -905 nw
rect 2856 -986 2871 -758
tri 2393 -1108 2399 -1102 se
rect 2399 -1108 2408 -1102
rect 2393 -1124 2408 -1108
tri 2408 -1115 2421 -1102 nw
rect 2562 -1110 2579 -1096
rect 2611 -1110 2628 -1096
tri 2755 -1102 2770 -1087 ne
tri 2770 -1102 2792 -1080 sw
rect 2393 -1160 2408 -1152
rect 2474 -1124 2534 -1110
rect 2489 -1134 2534 -1124
rect 2489 -1152 2517 -1134
tri 2393 -1175 2408 -1160 ne
tri 2408 -1175 2430 -1153 sw
rect 2474 -1162 2517 -1152
rect 2532 -1138 2534 -1134
rect 2656 -1124 2716 -1110
tri 2770 -1115 2783 -1102 ne
rect 2783 -1108 2792 -1102
tri 2792 -1108 2798 -1102 sw
rect 2656 -1134 2701 -1124
rect 2532 -1162 2606 -1138
rect 2474 -1166 2606 -1162
tri 2606 -1166 2634 -1138 sw
rect 2656 -1148 2658 -1134
tri 2656 -1150 2658 -1148 ne
rect 2670 -1152 2701 -1134
rect 2670 -1162 2716 -1152
rect 2783 -1123 2798 -1108
tri 2408 -1187 2420 -1175 ne
rect 2420 -1180 2430 -1175
tri 2430 -1180 2435 -1175 sw
rect 2319 -1526 2334 -1298
rect 2420 -1336 2435 -1180
rect 2474 -1222 2502 -1166
tri 2594 -1184 2612 -1166 ne
rect 2612 -1186 2634 -1166
tri 2634 -1186 2654 -1166 sw
tri 2670 -1180 2688 -1162 ne
rect 2493 -1256 2502 -1222
rect 2536 -1195 2578 -1194
rect 2536 -1229 2541 -1195
rect 2571 -1229 2578 -1195
rect 2536 -1238 2578 -1229
rect 2612 -1195 2654 -1186
rect 2612 -1229 2619 -1195
rect 2649 -1229 2654 -1195
rect 2612 -1234 2654 -1229
rect 2688 -1222 2716 -1162
tri 2761 -1175 2783 -1153 se
rect 2783 -1160 2798 -1152
tri 2783 -1175 2798 -1160 nw
tri 2755 -1181 2761 -1175 se
rect 2761 -1181 2770 -1175
rect 2474 -1266 2502 -1256
tri 2502 -1266 2526 -1242 sw
rect 2474 -1298 2516 -1266
tri 2533 -1274 2534 -1273 sw
rect 2533 -1298 2534 -1274
tri 2536 -1275 2573 -1238 ne
rect 2573 -1266 2578 -1238
tri 2578 -1266 2604 -1240 sw
rect 2688 -1256 2697 -1222
rect 2688 -1266 2716 -1256
rect 2573 -1275 2657 -1266
tri 2573 -1294 2592 -1275 ne
rect 2592 -1294 2657 -1275
rect 2474 -1320 2534 -1298
rect 2656 -1298 2657 -1294
rect 2674 -1298 2716 -1266
rect 2656 -1320 2716 -1298
rect 2562 -1336 2579 -1322
rect 2611 -1336 2628 -1322
tri 2399 -1372 2421 -1350 se
rect 2421 -1357 2436 -1336
tri 2421 -1372 2436 -1357 nw
rect 2755 -1357 2770 -1181
tri 2770 -1188 2783 -1175 nw
rect 2856 -1256 2871 -1028
tri 2393 -1378 2399 -1372 se
rect 2399 -1378 2408 -1372
rect 2393 -1394 2408 -1378
tri 2408 -1385 2421 -1372 nw
rect 2562 -1380 2579 -1366
rect 2611 -1380 2628 -1366
tri 2755 -1372 2770 -1357 ne
tri 2770 -1372 2792 -1350 sw
rect 2393 -1430 2408 -1422
rect 2474 -1394 2534 -1380
rect 2489 -1404 2534 -1394
rect 2489 -1422 2517 -1404
tri 2393 -1445 2408 -1430 ne
tri 2408 -1445 2430 -1423 sw
rect 2474 -1432 2517 -1422
rect 2532 -1408 2534 -1404
rect 2656 -1394 2716 -1380
tri 2770 -1385 2783 -1372 ne
rect 2783 -1378 2792 -1372
tri 2792 -1378 2798 -1372 sw
rect 2656 -1404 2701 -1394
rect 2532 -1432 2606 -1408
rect 2474 -1436 2606 -1432
tri 2606 -1436 2634 -1408 sw
rect 2656 -1418 2658 -1404
tri 2656 -1420 2658 -1418 ne
rect 2670 -1422 2701 -1404
rect 2670 -1432 2716 -1422
rect 2783 -1393 2798 -1378
tri 2408 -1457 2420 -1445 ne
rect 2420 -1450 2430 -1445
tri 2430 -1450 2435 -1445 sw
rect 2319 -1796 2334 -1568
rect 2420 -1606 2435 -1450
rect 2474 -1492 2502 -1436
tri 2594 -1454 2612 -1436 ne
rect 2612 -1456 2634 -1436
tri 2634 -1456 2654 -1436 sw
tri 2670 -1450 2688 -1432 ne
rect 2493 -1526 2502 -1492
rect 2536 -1465 2578 -1464
rect 2536 -1499 2541 -1465
rect 2571 -1499 2578 -1465
rect 2536 -1508 2578 -1499
rect 2612 -1465 2654 -1456
rect 2612 -1499 2619 -1465
rect 2649 -1499 2654 -1465
rect 2612 -1504 2654 -1499
rect 2688 -1492 2716 -1432
tri 2761 -1445 2783 -1423 se
rect 2783 -1430 2798 -1422
tri 2783 -1445 2798 -1430 nw
tri 2755 -1451 2761 -1445 se
rect 2761 -1451 2770 -1445
rect 2474 -1536 2502 -1526
tri 2502 -1536 2526 -1512 sw
rect 2474 -1568 2516 -1536
tri 2533 -1544 2534 -1543 sw
rect 2533 -1568 2534 -1544
tri 2536 -1545 2573 -1508 ne
rect 2573 -1536 2578 -1508
tri 2578 -1536 2604 -1510 sw
rect 2688 -1526 2697 -1492
rect 2688 -1536 2716 -1526
rect 2573 -1545 2657 -1536
tri 2573 -1564 2592 -1545 ne
rect 2592 -1564 2657 -1545
rect 2474 -1590 2534 -1568
rect 2656 -1568 2657 -1564
rect 2674 -1568 2716 -1536
rect 2656 -1590 2716 -1568
rect 2562 -1606 2579 -1592
rect 2611 -1606 2628 -1592
tri 2399 -1642 2421 -1620 se
rect 2421 -1627 2436 -1606
tri 2421 -1642 2436 -1627 nw
rect 2755 -1627 2770 -1451
tri 2770 -1458 2783 -1445 nw
rect 2856 -1526 2871 -1298
tri 2393 -1648 2399 -1642 se
rect 2399 -1648 2408 -1642
rect 2393 -1664 2408 -1648
tri 2408 -1655 2421 -1642 nw
rect 2562 -1650 2579 -1636
rect 2611 -1650 2628 -1636
tri 2755 -1642 2770 -1627 ne
tri 2770 -1642 2792 -1620 sw
rect 2393 -1700 2408 -1692
rect 2474 -1664 2534 -1650
rect 2489 -1674 2534 -1664
rect 2489 -1692 2517 -1674
tri 2393 -1715 2408 -1700 ne
tri 2408 -1715 2430 -1693 sw
rect 2474 -1702 2517 -1692
rect 2532 -1678 2534 -1674
rect 2656 -1664 2716 -1650
tri 2770 -1655 2783 -1642 ne
rect 2783 -1648 2792 -1642
tri 2792 -1648 2798 -1642 sw
rect 2656 -1674 2701 -1664
rect 2532 -1702 2606 -1678
rect 2474 -1706 2606 -1702
tri 2606 -1706 2634 -1678 sw
rect 2656 -1688 2658 -1674
tri 2656 -1690 2658 -1688 ne
rect 2670 -1692 2701 -1674
rect 2670 -1702 2716 -1692
rect 2783 -1663 2798 -1648
tri 2408 -1727 2420 -1715 ne
rect 2420 -1720 2430 -1715
tri 2430 -1720 2435 -1715 sw
rect 2319 -2066 2334 -1838
rect 2420 -1876 2435 -1720
rect 2474 -1762 2502 -1706
tri 2594 -1724 2612 -1706 ne
rect 2612 -1726 2634 -1706
tri 2634 -1726 2654 -1706 sw
tri 2670 -1720 2688 -1702 ne
rect 2493 -1796 2502 -1762
rect 2536 -1735 2578 -1734
rect 2536 -1769 2541 -1735
rect 2571 -1769 2578 -1735
rect 2536 -1778 2578 -1769
rect 2612 -1735 2654 -1726
rect 2612 -1769 2619 -1735
rect 2649 -1769 2654 -1735
rect 2612 -1774 2654 -1769
rect 2688 -1762 2716 -1702
tri 2761 -1715 2783 -1693 se
rect 2783 -1700 2798 -1692
tri 2783 -1715 2798 -1700 nw
tri 2755 -1721 2761 -1715 se
rect 2761 -1721 2770 -1715
rect 2474 -1806 2502 -1796
tri 2502 -1806 2526 -1782 sw
rect 2474 -1838 2516 -1806
tri 2533 -1814 2534 -1813 sw
rect 2533 -1838 2534 -1814
tri 2536 -1815 2573 -1778 ne
rect 2573 -1806 2578 -1778
tri 2578 -1806 2604 -1780 sw
rect 2688 -1796 2697 -1762
rect 2688 -1806 2716 -1796
rect 2573 -1815 2657 -1806
tri 2573 -1834 2592 -1815 ne
rect 2592 -1834 2657 -1815
rect 2474 -1860 2534 -1838
rect 2656 -1838 2657 -1834
rect 2674 -1838 2716 -1806
rect 2656 -1860 2716 -1838
rect 2562 -1876 2579 -1862
rect 2611 -1876 2628 -1862
tri 2399 -1912 2421 -1890 se
rect 2421 -1897 2436 -1876
tri 2421 -1912 2436 -1897 nw
rect 2755 -1897 2770 -1721
tri 2770 -1728 2783 -1715 nw
rect 2856 -1796 2871 -1568
tri 2393 -1918 2399 -1912 se
rect 2399 -1918 2408 -1912
rect 2393 -1934 2408 -1918
tri 2408 -1925 2421 -1912 nw
rect 2562 -1920 2579 -1906
rect 2611 -1920 2628 -1906
tri 2755 -1912 2770 -1897 ne
tri 2770 -1912 2792 -1890 sw
rect 2393 -1970 2408 -1962
rect 2474 -1934 2534 -1920
rect 2489 -1944 2534 -1934
rect 2489 -1962 2517 -1944
tri 2393 -1985 2408 -1970 ne
tri 2408 -1985 2430 -1963 sw
rect 2474 -1972 2517 -1962
rect 2532 -1948 2534 -1944
rect 2656 -1934 2716 -1920
tri 2770 -1925 2783 -1912 ne
rect 2783 -1918 2792 -1912
tri 2792 -1918 2798 -1912 sw
rect 2656 -1944 2701 -1934
rect 2532 -1972 2606 -1948
rect 2474 -1976 2606 -1972
tri 2606 -1976 2634 -1948 sw
rect 2656 -1958 2658 -1944
tri 2656 -1960 2658 -1958 ne
rect 2670 -1962 2701 -1944
rect 2670 -1972 2716 -1962
rect 2783 -1933 2798 -1918
tri 2408 -1997 2420 -1985 ne
rect 2420 -1990 2430 -1985
tri 2430 -1990 2435 -1985 sw
rect 2319 -2146 2334 -2108
rect 2420 -2146 2435 -1990
rect 2474 -2032 2502 -1976
tri 2594 -1994 2612 -1976 ne
rect 2612 -1996 2634 -1976
tri 2634 -1996 2654 -1976 sw
tri 2670 -1990 2688 -1972 ne
rect 2493 -2066 2502 -2032
rect 2536 -2005 2578 -2004
rect 2536 -2039 2541 -2005
rect 2571 -2039 2578 -2005
rect 2536 -2048 2578 -2039
rect 2612 -2005 2654 -1996
rect 2612 -2039 2619 -2005
rect 2649 -2039 2654 -2005
rect 2612 -2044 2654 -2039
rect 2688 -2032 2716 -1972
tri 2761 -1985 2783 -1963 se
rect 2783 -1970 2798 -1962
tri 2783 -1985 2798 -1970 nw
tri 2755 -1991 2761 -1985 se
rect 2761 -1991 2770 -1985
rect 2474 -2076 2502 -2066
tri 2502 -2076 2526 -2052 sw
rect 2474 -2108 2516 -2076
tri 2533 -2084 2534 -2083 sw
rect 2533 -2108 2534 -2084
tri 2536 -2085 2573 -2048 ne
rect 2573 -2076 2578 -2048
tri 2578 -2076 2604 -2050 sw
rect 2688 -2066 2697 -2032
rect 2688 -2076 2716 -2066
rect 2573 -2085 2657 -2076
tri 2573 -2104 2592 -2085 ne
rect 2592 -2104 2657 -2085
rect 2474 -2130 2534 -2108
rect 2656 -2108 2657 -2104
rect 2674 -2108 2716 -2076
rect 2656 -2130 2716 -2108
rect 2562 -2146 2579 -2132
rect 2611 -2146 2628 -2132
rect 2755 -2146 2770 -1991
tri 2770 -1998 2783 -1985 nw
rect 2856 -2066 2871 -1838
rect 2856 -2146 2871 -2108
rect 2899 1984 2914 2174
tri 2979 2138 3001 2160 se
rect 3001 2153 3016 2174
tri 3001 2138 3016 2153 nw
rect 3335 2153 3350 2174
tri 2973 2132 2979 2138 se
rect 2979 2132 2988 2138
rect 2973 2116 2988 2132
tri 2988 2125 3001 2138 nw
rect 3142 2130 3159 2144
rect 3191 2130 3208 2144
tri 3335 2138 3350 2153 ne
tri 3350 2138 3372 2160 sw
rect 2973 2080 2988 2088
rect 3054 2116 3114 2130
rect 3069 2106 3114 2116
rect 3069 2088 3097 2106
tri 2973 2065 2988 2080 ne
tri 2988 2065 3010 2087 sw
rect 3054 2078 3097 2088
rect 3112 2102 3114 2106
rect 3236 2116 3296 2130
tri 3350 2125 3363 2138 ne
rect 3363 2132 3372 2138
tri 3372 2132 3378 2138 sw
rect 3236 2106 3281 2116
rect 3112 2078 3186 2102
rect 3054 2074 3186 2078
tri 3186 2074 3214 2102 sw
rect 3236 2092 3238 2106
tri 3236 2090 3238 2092 ne
rect 3250 2088 3281 2106
rect 3250 2078 3296 2088
rect 3363 2117 3378 2132
tri 2988 2053 3000 2065 ne
rect 3000 2060 3010 2065
tri 3010 2060 3015 2065 sw
rect 2899 1714 2914 1942
rect 3000 1904 3015 2060
rect 3054 2018 3082 2074
tri 3174 2056 3192 2074 ne
rect 3192 2054 3214 2074
tri 3214 2054 3234 2074 sw
tri 3250 2060 3268 2078 ne
rect 3073 1984 3082 2018
rect 3116 2045 3158 2046
rect 3116 2011 3121 2045
rect 3151 2011 3158 2045
rect 3116 2002 3158 2011
rect 3192 2045 3234 2054
rect 3192 2011 3199 2045
rect 3229 2011 3234 2045
rect 3192 2006 3234 2011
rect 3268 2018 3296 2078
tri 3341 2065 3363 2087 se
rect 3363 2080 3378 2088
tri 3363 2065 3378 2080 nw
tri 3335 2059 3341 2065 se
rect 3341 2059 3350 2065
rect 3054 1974 3082 1984
tri 3082 1974 3106 1998 sw
rect 3054 1942 3096 1974
tri 3113 1966 3114 1967 sw
rect 3113 1942 3114 1966
tri 3116 1965 3153 2002 ne
rect 3153 1974 3158 2002
tri 3158 1974 3184 2000 sw
rect 3268 1984 3277 2018
rect 3268 1974 3296 1984
rect 3153 1965 3237 1974
tri 3153 1946 3172 1965 ne
rect 3172 1946 3237 1965
rect 3054 1920 3114 1942
rect 3236 1942 3237 1946
rect 3254 1942 3296 1974
rect 3236 1920 3296 1942
rect 3142 1904 3159 1918
rect 3191 1904 3208 1918
tri 2979 1868 3001 1890 se
rect 3001 1883 3016 1904
tri 3001 1868 3016 1883 nw
rect 3335 1883 3350 2059
tri 3350 2052 3363 2065 nw
rect 3436 1984 3451 2174
tri 2973 1862 2979 1868 se
rect 2979 1862 2988 1868
rect 2973 1846 2988 1862
tri 2988 1855 3001 1868 nw
rect 3142 1860 3159 1874
rect 3191 1860 3208 1874
tri 3335 1868 3350 1883 ne
tri 3350 1868 3372 1890 sw
rect 2973 1810 2988 1818
rect 3054 1846 3114 1860
rect 3069 1836 3114 1846
rect 3069 1818 3097 1836
tri 2973 1795 2988 1810 ne
tri 2988 1795 3010 1817 sw
rect 3054 1808 3097 1818
rect 3112 1832 3114 1836
rect 3236 1846 3296 1860
tri 3350 1855 3363 1868 ne
rect 3363 1862 3372 1868
tri 3372 1862 3378 1868 sw
rect 3236 1836 3281 1846
rect 3112 1808 3186 1832
rect 3054 1804 3186 1808
tri 3186 1804 3214 1832 sw
rect 3236 1822 3238 1836
tri 3236 1820 3238 1822 ne
rect 3250 1818 3281 1836
rect 3250 1808 3296 1818
rect 3363 1847 3378 1862
tri 2988 1783 3000 1795 ne
rect 3000 1790 3010 1795
tri 3010 1790 3015 1795 sw
rect 2899 1444 2914 1672
rect 3000 1634 3015 1790
rect 3054 1748 3082 1804
tri 3174 1786 3192 1804 ne
rect 3192 1784 3214 1804
tri 3214 1784 3234 1804 sw
tri 3250 1790 3268 1808 ne
rect 3073 1714 3082 1748
rect 3116 1775 3158 1776
rect 3116 1741 3121 1775
rect 3151 1741 3158 1775
rect 3116 1732 3158 1741
rect 3192 1775 3234 1784
rect 3192 1741 3199 1775
rect 3229 1741 3234 1775
rect 3192 1736 3234 1741
rect 3268 1748 3296 1808
tri 3341 1795 3363 1817 se
rect 3363 1810 3378 1818
tri 3363 1795 3378 1810 nw
tri 3335 1789 3341 1795 se
rect 3341 1789 3350 1795
rect 3054 1704 3082 1714
tri 3082 1704 3106 1728 sw
rect 3054 1672 3096 1704
tri 3113 1696 3114 1697 sw
rect 3113 1672 3114 1696
tri 3116 1695 3153 1732 ne
rect 3153 1704 3158 1732
tri 3158 1704 3184 1730 sw
rect 3268 1714 3277 1748
rect 3268 1704 3296 1714
rect 3153 1695 3237 1704
tri 3153 1676 3172 1695 ne
rect 3172 1676 3237 1695
rect 3054 1650 3114 1672
rect 3236 1672 3237 1676
rect 3254 1672 3296 1704
rect 3236 1650 3296 1672
rect 3142 1634 3159 1648
rect 3191 1634 3208 1648
tri 2979 1598 3001 1620 se
rect 3001 1613 3016 1634
tri 3001 1598 3016 1613 nw
rect 3335 1613 3350 1789
tri 3350 1782 3363 1795 nw
rect 3436 1714 3451 1942
tri 2973 1592 2979 1598 se
rect 2979 1592 2988 1598
rect 2973 1576 2988 1592
tri 2988 1585 3001 1598 nw
rect 3142 1590 3159 1604
rect 3191 1590 3208 1604
tri 3335 1598 3350 1613 ne
tri 3350 1598 3372 1620 sw
rect 2973 1540 2988 1548
rect 3054 1576 3114 1590
rect 3069 1566 3114 1576
rect 3069 1548 3097 1566
tri 2973 1525 2988 1540 ne
tri 2988 1525 3010 1547 sw
rect 3054 1538 3097 1548
rect 3112 1562 3114 1566
rect 3236 1576 3296 1590
tri 3350 1585 3363 1598 ne
rect 3363 1592 3372 1598
tri 3372 1592 3378 1598 sw
rect 3236 1566 3281 1576
rect 3112 1538 3186 1562
rect 3054 1534 3186 1538
tri 3186 1534 3214 1562 sw
rect 3236 1552 3238 1566
tri 3236 1550 3238 1552 ne
rect 3250 1548 3281 1566
rect 3250 1538 3296 1548
rect 3363 1577 3378 1592
tri 2988 1513 3000 1525 ne
rect 3000 1520 3010 1525
tri 3010 1520 3015 1525 sw
rect 2899 1174 2914 1402
rect 3000 1364 3015 1520
rect 3054 1478 3082 1534
tri 3174 1516 3192 1534 ne
rect 3192 1514 3214 1534
tri 3214 1514 3234 1534 sw
tri 3250 1520 3268 1538 ne
rect 3073 1444 3082 1478
rect 3116 1505 3158 1506
rect 3116 1471 3121 1505
rect 3151 1471 3158 1505
rect 3116 1462 3158 1471
rect 3192 1505 3234 1514
rect 3192 1471 3199 1505
rect 3229 1471 3234 1505
rect 3192 1466 3234 1471
rect 3268 1478 3296 1538
tri 3341 1525 3363 1547 se
rect 3363 1540 3378 1548
tri 3363 1525 3378 1540 nw
tri 3335 1519 3341 1525 se
rect 3341 1519 3350 1525
rect 3054 1434 3082 1444
tri 3082 1434 3106 1458 sw
rect 3054 1402 3096 1434
tri 3113 1426 3114 1427 sw
rect 3113 1402 3114 1426
tri 3116 1425 3153 1462 ne
rect 3153 1434 3158 1462
tri 3158 1434 3184 1460 sw
rect 3268 1444 3277 1478
rect 3268 1434 3296 1444
rect 3153 1425 3237 1434
tri 3153 1406 3172 1425 ne
rect 3172 1406 3237 1425
rect 3054 1380 3114 1402
rect 3236 1402 3237 1406
rect 3254 1402 3296 1434
rect 3236 1380 3296 1402
rect 3142 1364 3159 1378
rect 3191 1364 3208 1378
tri 2979 1328 3001 1350 se
rect 3001 1343 3016 1364
tri 3001 1328 3016 1343 nw
rect 3335 1343 3350 1519
tri 3350 1512 3363 1525 nw
rect 3436 1444 3451 1672
tri 2973 1322 2979 1328 se
rect 2979 1322 2988 1328
rect 2973 1306 2988 1322
tri 2988 1315 3001 1328 nw
rect 3142 1320 3159 1334
rect 3191 1320 3208 1334
tri 3335 1328 3350 1343 ne
tri 3350 1328 3372 1350 sw
rect 2973 1270 2988 1278
rect 3054 1306 3114 1320
rect 3069 1296 3114 1306
rect 3069 1278 3097 1296
tri 2973 1255 2988 1270 ne
tri 2988 1255 3010 1277 sw
rect 3054 1268 3097 1278
rect 3112 1292 3114 1296
rect 3236 1306 3296 1320
tri 3350 1315 3363 1328 ne
rect 3363 1322 3372 1328
tri 3372 1322 3378 1328 sw
rect 3236 1296 3281 1306
rect 3112 1268 3186 1292
rect 3054 1264 3186 1268
tri 3186 1264 3214 1292 sw
rect 3236 1282 3238 1296
tri 3236 1280 3238 1282 ne
rect 3250 1278 3281 1296
rect 3250 1268 3296 1278
rect 3363 1307 3378 1322
tri 2988 1243 3000 1255 ne
rect 3000 1250 3010 1255
tri 3010 1250 3015 1255 sw
rect 2899 904 2914 1132
rect 3000 1094 3015 1250
rect 3054 1208 3082 1264
tri 3174 1246 3192 1264 ne
rect 3192 1244 3214 1264
tri 3214 1244 3234 1264 sw
tri 3250 1250 3268 1268 ne
rect 3073 1174 3082 1208
rect 3116 1235 3158 1236
rect 3116 1201 3121 1235
rect 3151 1201 3158 1235
rect 3116 1192 3158 1201
rect 3192 1235 3234 1244
rect 3192 1201 3199 1235
rect 3229 1201 3234 1235
rect 3192 1196 3234 1201
rect 3268 1208 3296 1268
tri 3341 1255 3363 1277 se
rect 3363 1270 3378 1278
tri 3363 1255 3378 1270 nw
tri 3335 1249 3341 1255 se
rect 3341 1249 3350 1255
rect 3054 1164 3082 1174
tri 3082 1164 3106 1188 sw
rect 3054 1132 3096 1164
tri 3113 1156 3114 1157 sw
rect 3113 1132 3114 1156
tri 3116 1155 3153 1192 ne
rect 3153 1164 3158 1192
tri 3158 1164 3184 1190 sw
rect 3268 1174 3277 1208
rect 3268 1164 3296 1174
rect 3153 1155 3237 1164
tri 3153 1136 3172 1155 ne
rect 3172 1136 3237 1155
rect 3054 1110 3114 1132
rect 3236 1132 3237 1136
rect 3254 1132 3296 1164
rect 3236 1110 3296 1132
rect 3142 1094 3159 1108
rect 3191 1094 3208 1108
tri 2979 1058 3001 1080 se
rect 3001 1073 3016 1094
tri 3001 1058 3016 1073 nw
rect 3335 1073 3350 1249
tri 3350 1242 3363 1255 nw
rect 3436 1174 3451 1402
tri 2973 1052 2979 1058 se
rect 2979 1052 2988 1058
rect 2973 1036 2988 1052
tri 2988 1045 3001 1058 nw
rect 3142 1050 3159 1064
rect 3191 1050 3208 1064
tri 3335 1058 3350 1073 ne
tri 3350 1058 3372 1080 sw
rect 2973 1000 2988 1008
rect 3054 1036 3114 1050
rect 3069 1026 3114 1036
rect 3069 1008 3097 1026
tri 2973 985 2988 1000 ne
tri 2988 985 3010 1007 sw
rect 3054 998 3097 1008
rect 3112 1022 3114 1026
rect 3236 1036 3296 1050
tri 3350 1045 3363 1058 ne
rect 3363 1052 3372 1058
tri 3372 1052 3378 1058 sw
rect 3236 1026 3281 1036
rect 3112 998 3186 1022
rect 3054 994 3186 998
tri 3186 994 3214 1022 sw
rect 3236 1012 3238 1026
tri 3236 1010 3238 1012 ne
rect 3250 1008 3281 1026
rect 3250 998 3296 1008
rect 3363 1037 3378 1052
tri 2988 973 3000 985 ne
rect 3000 980 3010 985
tri 3010 980 3015 985 sw
rect 2899 634 2914 862
rect 3000 824 3015 980
rect 3054 938 3082 994
tri 3174 976 3192 994 ne
rect 3192 974 3214 994
tri 3214 974 3234 994 sw
tri 3250 980 3268 998 ne
rect 3073 904 3082 938
rect 3116 965 3158 966
rect 3116 931 3121 965
rect 3151 931 3158 965
rect 3116 922 3158 931
rect 3192 965 3234 974
rect 3192 931 3199 965
rect 3229 931 3234 965
rect 3192 926 3234 931
rect 3268 938 3296 998
tri 3341 985 3363 1007 se
rect 3363 1000 3378 1008
tri 3363 985 3378 1000 nw
tri 3335 979 3341 985 se
rect 3341 979 3350 985
rect 3054 894 3082 904
tri 3082 894 3106 918 sw
rect 3054 862 3096 894
tri 3113 886 3114 887 sw
rect 3113 862 3114 886
tri 3116 885 3153 922 ne
rect 3153 894 3158 922
tri 3158 894 3184 920 sw
rect 3268 904 3277 938
rect 3268 894 3296 904
rect 3153 885 3237 894
tri 3153 866 3172 885 ne
rect 3172 866 3237 885
rect 3054 840 3114 862
rect 3236 862 3237 866
rect 3254 862 3296 894
rect 3236 840 3296 862
rect 3142 824 3159 838
rect 3191 824 3208 838
tri 2979 788 3001 810 se
rect 3001 803 3016 824
tri 3001 788 3016 803 nw
rect 3335 803 3350 979
tri 3350 972 3363 985 nw
rect 3436 904 3451 1132
tri 2973 782 2979 788 se
rect 2979 782 2988 788
rect 2973 766 2988 782
tri 2988 775 3001 788 nw
rect 3142 780 3159 794
rect 3191 780 3208 794
tri 3335 788 3350 803 ne
tri 3350 788 3372 810 sw
rect 2973 730 2988 738
rect 3054 766 3114 780
rect 3069 756 3114 766
rect 3069 738 3097 756
tri 2973 715 2988 730 ne
tri 2988 715 3010 737 sw
rect 3054 728 3097 738
rect 3112 752 3114 756
rect 3236 766 3296 780
tri 3350 775 3363 788 ne
rect 3363 782 3372 788
tri 3372 782 3378 788 sw
rect 3236 756 3281 766
rect 3112 728 3186 752
rect 3054 724 3186 728
tri 3186 724 3214 752 sw
rect 3236 742 3238 756
tri 3236 740 3238 742 ne
rect 3250 738 3281 756
rect 3250 728 3296 738
rect 3363 767 3378 782
tri 2988 703 3000 715 ne
rect 3000 710 3010 715
tri 3010 710 3015 715 sw
rect 2899 364 2914 592
rect 3000 554 3015 710
rect 3054 668 3082 724
tri 3174 706 3192 724 ne
rect 3192 704 3214 724
tri 3214 704 3234 724 sw
tri 3250 710 3268 728 ne
rect 3073 634 3082 668
rect 3116 695 3158 696
rect 3116 661 3121 695
rect 3151 661 3158 695
rect 3116 652 3158 661
rect 3192 695 3234 704
rect 3192 661 3199 695
rect 3229 661 3234 695
rect 3192 656 3234 661
rect 3268 668 3296 728
tri 3341 715 3363 737 se
rect 3363 730 3378 738
tri 3363 715 3378 730 nw
tri 3335 709 3341 715 se
rect 3341 709 3350 715
rect 3054 624 3082 634
tri 3082 624 3106 648 sw
rect 3054 592 3096 624
tri 3113 616 3114 617 sw
rect 3113 592 3114 616
tri 3116 615 3153 652 ne
rect 3153 624 3158 652
tri 3158 624 3184 650 sw
rect 3268 634 3277 668
rect 3268 624 3296 634
rect 3153 615 3237 624
tri 3153 596 3172 615 ne
rect 3172 596 3237 615
rect 3054 570 3114 592
rect 3236 592 3237 596
rect 3254 592 3296 624
rect 3236 570 3296 592
rect 3142 554 3159 568
rect 3191 554 3208 568
tri 2979 518 3001 540 se
rect 3001 533 3016 554
tri 3001 518 3016 533 nw
rect 3335 533 3350 709
tri 3350 702 3363 715 nw
rect 3436 634 3451 862
tri 2973 512 2979 518 se
rect 2979 512 2988 518
rect 2973 496 2988 512
tri 2988 505 3001 518 nw
rect 3142 510 3159 524
rect 3191 510 3208 524
tri 3335 518 3350 533 ne
tri 3350 518 3372 540 sw
rect 2973 460 2988 468
rect 3054 496 3114 510
rect 3069 486 3114 496
rect 3069 468 3097 486
tri 2973 445 2988 460 ne
tri 2988 445 3010 467 sw
rect 3054 458 3097 468
rect 3112 482 3114 486
rect 3236 496 3296 510
tri 3350 505 3363 518 ne
rect 3363 512 3372 518
tri 3372 512 3378 518 sw
rect 3236 486 3281 496
rect 3112 458 3186 482
rect 3054 454 3186 458
tri 3186 454 3214 482 sw
rect 3236 472 3238 486
tri 3236 470 3238 472 ne
rect 3250 468 3281 486
rect 3250 458 3296 468
rect 3363 497 3378 512
tri 2988 433 3000 445 ne
rect 3000 440 3010 445
tri 3010 440 3015 445 sw
rect 2899 94 2914 322
rect 3000 284 3015 440
rect 3054 398 3082 454
tri 3174 436 3192 454 ne
rect 3192 434 3214 454
tri 3214 434 3234 454 sw
tri 3250 440 3268 458 ne
rect 3073 364 3082 398
rect 3116 425 3158 426
rect 3116 391 3121 425
rect 3151 391 3158 425
rect 3116 382 3158 391
rect 3192 425 3234 434
rect 3192 391 3199 425
rect 3229 391 3234 425
rect 3192 386 3234 391
rect 3268 398 3296 458
tri 3341 445 3363 467 se
rect 3363 460 3378 468
tri 3363 445 3378 460 nw
tri 3335 439 3341 445 se
rect 3341 439 3350 445
rect 3054 354 3082 364
tri 3082 354 3106 378 sw
rect 3054 322 3096 354
tri 3113 346 3114 347 sw
rect 3113 322 3114 346
tri 3116 345 3153 382 ne
rect 3153 354 3158 382
tri 3158 354 3184 380 sw
rect 3268 364 3277 398
rect 3268 354 3296 364
rect 3153 345 3237 354
tri 3153 326 3172 345 ne
rect 3172 326 3237 345
rect 3054 300 3114 322
rect 3236 322 3237 326
rect 3254 322 3296 354
rect 3236 300 3296 322
rect 3142 284 3159 298
rect 3191 284 3208 298
tri 2979 248 3001 270 se
rect 3001 263 3016 284
tri 3001 248 3016 263 nw
rect 3335 263 3350 439
tri 3350 432 3363 445 nw
rect 3436 364 3451 592
tri 2973 242 2979 248 se
rect 2979 242 2988 248
rect 2973 226 2988 242
tri 2988 235 3001 248 nw
rect 3142 240 3159 254
rect 3191 240 3208 254
tri 3335 248 3350 263 ne
tri 3350 248 3372 270 sw
rect 2973 190 2988 198
rect 3054 226 3114 240
rect 3069 216 3114 226
rect 3069 198 3097 216
tri 2973 175 2988 190 ne
tri 2988 175 3010 197 sw
rect 3054 188 3097 198
rect 3112 212 3114 216
rect 3236 226 3296 240
tri 3350 235 3363 248 ne
rect 3363 242 3372 248
tri 3372 242 3378 248 sw
rect 3236 216 3281 226
rect 3112 188 3186 212
rect 3054 184 3186 188
tri 3186 184 3214 212 sw
rect 3236 202 3238 216
tri 3236 200 3238 202 ne
rect 3250 198 3281 216
rect 3250 188 3296 198
rect 3363 227 3378 242
tri 2988 163 3000 175 ne
rect 3000 170 3010 175
tri 3010 170 3015 175 sw
rect 2899 -176 2914 52
rect 3000 14 3015 170
rect 3054 128 3082 184
tri 3174 166 3192 184 ne
rect 3192 164 3214 184
tri 3214 164 3234 184 sw
tri 3250 170 3268 188 ne
rect 3073 94 3082 128
rect 3116 155 3158 156
rect 3116 121 3121 155
rect 3151 121 3158 155
rect 3116 112 3158 121
rect 3192 155 3234 164
rect 3192 121 3199 155
rect 3229 121 3234 155
rect 3192 116 3234 121
rect 3268 128 3296 188
tri 3341 175 3363 197 se
rect 3363 190 3378 198
tri 3363 175 3378 190 nw
tri 3335 169 3341 175 se
rect 3341 169 3350 175
rect 3054 84 3082 94
tri 3082 84 3106 108 sw
rect 3054 52 3096 84
tri 3113 76 3114 77 sw
rect 3113 52 3114 76
tri 3116 75 3153 112 ne
rect 3153 84 3158 112
tri 3158 84 3184 110 sw
rect 3268 94 3277 128
rect 3268 84 3296 94
rect 3153 75 3237 84
tri 3153 56 3172 75 ne
rect 3172 56 3237 75
rect 3054 30 3114 52
rect 3236 52 3237 56
rect 3254 52 3296 84
rect 3236 30 3296 52
rect 3142 14 3159 28
rect 3191 14 3208 28
tri 2979 -22 3001 0 se
rect 3001 -7 3016 14
tri 3001 -22 3016 -7 nw
rect 3335 -7 3350 169
tri 3350 162 3363 175 nw
rect 3436 94 3451 322
tri 2973 -28 2979 -22 se
rect 2979 -28 2988 -22
rect 2973 -44 2988 -28
tri 2988 -35 3001 -22 nw
rect 3142 -30 3159 -16
rect 3191 -30 3208 -16
tri 3335 -22 3350 -7 ne
tri 3350 -22 3372 0 sw
rect 2973 -80 2988 -72
rect 3054 -44 3114 -30
rect 3069 -54 3114 -44
rect 3069 -72 3097 -54
tri 2973 -95 2988 -80 ne
tri 2988 -95 3010 -73 sw
rect 3054 -82 3097 -72
rect 3112 -58 3114 -54
rect 3236 -44 3296 -30
tri 3350 -35 3363 -22 ne
rect 3363 -28 3372 -22
tri 3372 -28 3378 -22 sw
rect 3236 -54 3281 -44
rect 3112 -82 3186 -58
rect 3054 -86 3186 -82
tri 3186 -86 3214 -58 sw
rect 3236 -68 3238 -54
tri 3236 -70 3238 -68 ne
rect 3250 -72 3281 -54
rect 3250 -82 3296 -72
rect 3363 -43 3378 -28
tri 2988 -107 3000 -95 ne
rect 3000 -100 3010 -95
tri 3010 -100 3015 -95 sw
rect 2899 -446 2914 -218
rect 3000 -256 3015 -100
rect 3054 -142 3082 -86
tri 3174 -104 3192 -86 ne
rect 3192 -106 3214 -86
tri 3214 -106 3234 -86 sw
tri 3250 -100 3268 -82 ne
rect 3073 -176 3082 -142
rect 3116 -115 3158 -114
rect 3116 -149 3121 -115
rect 3151 -149 3158 -115
rect 3116 -158 3158 -149
rect 3192 -115 3234 -106
rect 3192 -149 3199 -115
rect 3229 -149 3234 -115
rect 3192 -154 3234 -149
rect 3268 -142 3296 -82
tri 3341 -95 3363 -73 se
rect 3363 -80 3378 -72
tri 3363 -95 3378 -80 nw
tri 3335 -101 3341 -95 se
rect 3341 -101 3350 -95
rect 3054 -186 3082 -176
tri 3082 -186 3106 -162 sw
rect 3054 -218 3096 -186
tri 3113 -194 3114 -193 sw
rect 3113 -218 3114 -194
tri 3116 -195 3153 -158 ne
rect 3153 -186 3158 -158
tri 3158 -186 3184 -160 sw
rect 3268 -176 3277 -142
rect 3268 -186 3296 -176
rect 3153 -195 3237 -186
tri 3153 -214 3172 -195 ne
rect 3172 -214 3237 -195
rect 3054 -240 3114 -218
rect 3236 -218 3237 -214
rect 3254 -218 3296 -186
rect 3236 -240 3296 -218
rect 3142 -256 3159 -242
rect 3191 -256 3208 -242
tri 2979 -292 3001 -270 se
rect 3001 -277 3016 -256
tri 3001 -292 3016 -277 nw
rect 3335 -277 3350 -101
tri 3350 -108 3363 -95 nw
rect 3436 -176 3451 52
tri 2973 -298 2979 -292 se
rect 2979 -298 2988 -292
rect 2973 -314 2988 -298
tri 2988 -305 3001 -292 nw
rect 3142 -300 3159 -286
rect 3191 -300 3208 -286
tri 3335 -292 3350 -277 ne
tri 3350 -292 3372 -270 sw
rect 2973 -350 2988 -342
rect 3054 -314 3114 -300
rect 3069 -324 3114 -314
rect 3069 -342 3097 -324
tri 2973 -365 2988 -350 ne
tri 2988 -365 3010 -343 sw
rect 3054 -352 3097 -342
rect 3112 -328 3114 -324
rect 3236 -314 3296 -300
tri 3350 -305 3363 -292 ne
rect 3363 -298 3372 -292
tri 3372 -298 3378 -292 sw
rect 3236 -324 3281 -314
rect 3112 -352 3186 -328
rect 3054 -356 3186 -352
tri 3186 -356 3214 -328 sw
rect 3236 -338 3238 -324
tri 3236 -340 3238 -338 ne
rect 3250 -342 3281 -324
rect 3250 -352 3296 -342
rect 3363 -313 3378 -298
tri 2988 -377 3000 -365 ne
rect 3000 -370 3010 -365
tri 3010 -370 3015 -365 sw
rect 2899 -716 2914 -488
rect 3000 -526 3015 -370
rect 3054 -412 3082 -356
tri 3174 -374 3192 -356 ne
rect 3192 -376 3214 -356
tri 3214 -376 3234 -356 sw
tri 3250 -370 3268 -352 ne
rect 3073 -446 3082 -412
rect 3116 -385 3158 -384
rect 3116 -419 3121 -385
rect 3151 -419 3158 -385
rect 3116 -428 3158 -419
rect 3192 -385 3234 -376
rect 3192 -419 3199 -385
rect 3229 -419 3234 -385
rect 3192 -424 3234 -419
rect 3268 -412 3296 -352
tri 3341 -365 3363 -343 se
rect 3363 -350 3378 -342
tri 3363 -365 3378 -350 nw
tri 3335 -371 3341 -365 se
rect 3341 -371 3350 -365
rect 3054 -456 3082 -446
tri 3082 -456 3106 -432 sw
rect 3054 -488 3096 -456
tri 3113 -464 3114 -463 sw
rect 3113 -488 3114 -464
tri 3116 -465 3153 -428 ne
rect 3153 -456 3158 -428
tri 3158 -456 3184 -430 sw
rect 3268 -446 3277 -412
rect 3268 -456 3296 -446
rect 3153 -465 3237 -456
tri 3153 -484 3172 -465 ne
rect 3172 -484 3237 -465
rect 3054 -510 3114 -488
rect 3236 -488 3237 -484
rect 3254 -488 3296 -456
rect 3236 -510 3296 -488
rect 3142 -526 3159 -512
rect 3191 -526 3208 -512
tri 2979 -562 3001 -540 se
rect 3001 -547 3016 -526
tri 3001 -562 3016 -547 nw
rect 3335 -547 3350 -371
tri 3350 -378 3363 -365 nw
rect 3436 -446 3451 -218
tri 2973 -568 2979 -562 se
rect 2979 -568 2988 -562
rect 2973 -584 2988 -568
tri 2988 -575 3001 -562 nw
rect 3142 -570 3159 -556
rect 3191 -570 3208 -556
tri 3335 -562 3350 -547 ne
tri 3350 -562 3372 -540 sw
rect 2973 -620 2988 -612
rect 3054 -584 3114 -570
rect 3069 -594 3114 -584
rect 3069 -612 3097 -594
tri 2973 -635 2988 -620 ne
tri 2988 -635 3010 -613 sw
rect 3054 -622 3097 -612
rect 3112 -598 3114 -594
rect 3236 -584 3296 -570
tri 3350 -575 3363 -562 ne
rect 3363 -568 3372 -562
tri 3372 -568 3378 -562 sw
rect 3236 -594 3281 -584
rect 3112 -622 3186 -598
rect 3054 -626 3186 -622
tri 3186 -626 3214 -598 sw
rect 3236 -608 3238 -594
tri 3236 -610 3238 -608 ne
rect 3250 -612 3281 -594
rect 3250 -622 3296 -612
rect 3363 -583 3378 -568
tri 2988 -647 3000 -635 ne
rect 3000 -640 3010 -635
tri 3010 -640 3015 -635 sw
rect 2899 -986 2914 -758
rect 3000 -796 3015 -640
rect 3054 -682 3082 -626
tri 3174 -644 3192 -626 ne
rect 3192 -646 3214 -626
tri 3214 -646 3234 -626 sw
tri 3250 -640 3268 -622 ne
rect 3073 -716 3082 -682
rect 3116 -655 3158 -654
rect 3116 -689 3121 -655
rect 3151 -689 3158 -655
rect 3116 -698 3158 -689
rect 3192 -655 3234 -646
rect 3192 -689 3199 -655
rect 3229 -689 3234 -655
rect 3192 -694 3234 -689
rect 3268 -682 3296 -622
tri 3341 -635 3363 -613 se
rect 3363 -620 3378 -612
tri 3363 -635 3378 -620 nw
tri 3335 -641 3341 -635 se
rect 3341 -641 3350 -635
rect 3054 -726 3082 -716
tri 3082 -726 3106 -702 sw
rect 3054 -758 3096 -726
tri 3113 -734 3114 -733 sw
rect 3113 -758 3114 -734
tri 3116 -735 3153 -698 ne
rect 3153 -726 3158 -698
tri 3158 -726 3184 -700 sw
rect 3268 -716 3277 -682
rect 3268 -726 3296 -716
rect 3153 -735 3237 -726
tri 3153 -754 3172 -735 ne
rect 3172 -754 3237 -735
rect 3054 -780 3114 -758
rect 3236 -758 3237 -754
rect 3254 -758 3296 -726
rect 3236 -780 3296 -758
rect 3142 -796 3159 -782
rect 3191 -796 3208 -782
tri 2979 -832 3001 -810 se
rect 3001 -817 3016 -796
tri 3001 -832 3016 -817 nw
rect 3335 -817 3350 -641
tri 3350 -648 3363 -635 nw
rect 3436 -716 3451 -488
tri 2973 -838 2979 -832 se
rect 2979 -838 2988 -832
rect 2973 -854 2988 -838
tri 2988 -845 3001 -832 nw
rect 3142 -840 3159 -826
rect 3191 -840 3208 -826
tri 3335 -832 3350 -817 ne
tri 3350 -832 3372 -810 sw
rect 2973 -890 2988 -882
rect 3054 -854 3114 -840
rect 3069 -864 3114 -854
rect 3069 -882 3097 -864
tri 2973 -905 2988 -890 ne
tri 2988 -905 3010 -883 sw
rect 3054 -892 3097 -882
rect 3112 -868 3114 -864
rect 3236 -854 3296 -840
tri 3350 -845 3363 -832 ne
rect 3363 -838 3372 -832
tri 3372 -838 3378 -832 sw
rect 3236 -864 3281 -854
rect 3112 -892 3186 -868
rect 3054 -896 3186 -892
tri 3186 -896 3214 -868 sw
rect 3236 -878 3238 -864
tri 3236 -880 3238 -878 ne
rect 3250 -882 3281 -864
rect 3250 -892 3296 -882
rect 3363 -853 3378 -838
tri 2988 -917 3000 -905 ne
rect 3000 -910 3010 -905
tri 3010 -910 3015 -905 sw
rect 2899 -1256 2914 -1028
rect 3000 -1066 3015 -910
rect 3054 -952 3082 -896
tri 3174 -914 3192 -896 ne
rect 3192 -916 3214 -896
tri 3214 -916 3234 -896 sw
tri 3250 -910 3268 -892 ne
rect 3073 -986 3082 -952
rect 3116 -925 3158 -924
rect 3116 -959 3121 -925
rect 3151 -959 3158 -925
rect 3116 -968 3158 -959
rect 3192 -925 3234 -916
rect 3192 -959 3199 -925
rect 3229 -959 3234 -925
rect 3192 -964 3234 -959
rect 3268 -952 3296 -892
tri 3341 -905 3363 -883 se
rect 3363 -890 3378 -882
tri 3363 -905 3378 -890 nw
tri 3335 -911 3341 -905 se
rect 3341 -911 3350 -905
rect 3054 -996 3082 -986
tri 3082 -996 3106 -972 sw
rect 3054 -1028 3096 -996
tri 3113 -1004 3114 -1003 sw
rect 3113 -1028 3114 -1004
tri 3116 -1005 3153 -968 ne
rect 3153 -996 3158 -968
tri 3158 -996 3184 -970 sw
rect 3268 -986 3277 -952
rect 3268 -996 3296 -986
rect 3153 -1005 3237 -996
tri 3153 -1024 3172 -1005 ne
rect 3172 -1024 3237 -1005
rect 3054 -1050 3114 -1028
rect 3236 -1028 3237 -1024
rect 3254 -1028 3296 -996
rect 3236 -1050 3296 -1028
rect 3142 -1066 3159 -1052
rect 3191 -1066 3208 -1052
tri 2979 -1102 3001 -1080 se
rect 3001 -1087 3016 -1066
tri 3001 -1102 3016 -1087 nw
rect 3335 -1087 3350 -911
tri 3350 -918 3363 -905 nw
rect 3436 -986 3451 -758
tri 2973 -1108 2979 -1102 se
rect 2979 -1108 2988 -1102
rect 2973 -1124 2988 -1108
tri 2988 -1115 3001 -1102 nw
rect 3142 -1110 3159 -1096
rect 3191 -1110 3208 -1096
tri 3335 -1102 3350 -1087 ne
tri 3350 -1102 3372 -1080 sw
rect 2973 -1160 2988 -1152
rect 3054 -1124 3114 -1110
rect 3069 -1134 3114 -1124
rect 3069 -1152 3097 -1134
tri 2973 -1175 2988 -1160 ne
tri 2988 -1175 3010 -1153 sw
rect 3054 -1162 3097 -1152
rect 3112 -1138 3114 -1134
rect 3236 -1124 3296 -1110
tri 3350 -1115 3363 -1102 ne
rect 3363 -1108 3372 -1102
tri 3372 -1108 3378 -1102 sw
rect 3236 -1134 3281 -1124
rect 3112 -1162 3186 -1138
rect 3054 -1166 3186 -1162
tri 3186 -1166 3214 -1138 sw
rect 3236 -1148 3238 -1134
tri 3236 -1150 3238 -1148 ne
rect 3250 -1152 3281 -1134
rect 3250 -1162 3296 -1152
rect 3363 -1123 3378 -1108
tri 2988 -1187 3000 -1175 ne
rect 3000 -1180 3010 -1175
tri 3010 -1180 3015 -1175 sw
rect 2899 -1526 2914 -1298
rect 3000 -1336 3015 -1180
rect 3054 -1222 3082 -1166
tri 3174 -1184 3192 -1166 ne
rect 3192 -1186 3214 -1166
tri 3214 -1186 3234 -1166 sw
tri 3250 -1180 3268 -1162 ne
rect 3073 -1256 3082 -1222
rect 3116 -1195 3158 -1194
rect 3116 -1229 3121 -1195
rect 3151 -1229 3158 -1195
rect 3116 -1238 3158 -1229
rect 3192 -1195 3234 -1186
rect 3192 -1229 3199 -1195
rect 3229 -1229 3234 -1195
rect 3192 -1234 3234 -1229
rect 3268 -1222 3296 -1162
tri 3341 -1175 3363 -1153 se
rect 3363 -1160 3378 -1152
tri 3363 -1175 3378 -1160 nw
tri 3335 -1181 3341 -1175 se
rect 3341 -1181 3350 -1175
rect 3054 -1266 3082 -1256
tri 3082 -1266 3106 -1242 sw
rect 3054 -1298 3096 -1266
tri 3113 -1274 3114 -1273 sw
rect 3113 -1298 3114 -1274
tri 3116 -1275 3153 -1238 ne
rect 3153 -1266 3158 -1238
tri 3158 -1266 3184 -1240 sw
rect 3268 -1256 3277 -1222
rect 3268 -1266 3296 -1256
rect 3153 -1275 3237 -1266
tri 3153 -1294 3172 -1275 ne
rect 3172 -1294 3237 -1275
rect 3054 -1320 3114 -1298
rect 3236 -1298 3237 -1294
rect 3254 -1298 3296 -1266
rect 3236 -1320 3296 -1298
rect 3142 -1336 3159 -1322
rect 3191 -1336 3208 -1322
tri 2979 -1372 3001 -1350 se
rect 3001 -1357 3016 -1336
tri 3001 -1372 3016 -1357 nw
rect 3335 -1357 3350 -1181
tri 3350 -1188 3363 -1175 nw
rect 3436 -1256 3451 -1028
tri 2973 -1378 2979 -1372 se
rect 2979 -1378 2988 -1372
rect 2973 -1394 2988 -1378
tri 2988 -1385 3001 -1372 nw
rect 3142 -1380 3159 -1366
rect 3191 -1380 3208 -1366
tri 3335 -1372 3350 -1357 ne
tri 3350 -1372 3372 -1350 sw
rect 2973 -1430 2988 -1422
rect 3054 -1394 3114 -1380
rect 3069 -1404 3114 -1394
rect 3069 -1422 3097 -1404
tri 2973 -1445 2988 -1430 ne
tri 2988 -1445 3010 -1423 sw
rect 3054 -1432 3097 -1422
rect 3112 -1408 3114 -1404
rect 3236 -1394 3296 -1380
tri 3350 -1385 3363 -1372 ne
rect 3363 -1378 3372 -1372
tri 3372 -1378 3378 -1372 sw
rect 3236 -1404 3281 -1394
rect 3112 -1432 3186 -1408
rect 3054 -1436 3186 -1432
tri 3186 -1436 3214 -1408 sw
rect 3236 -1418 3238 -1404
tri 3236 -1420 3238 -1418 ne
rect 3250 -1422 3281 -1404
rect 3250 -1432 3296 -1422
rect 3363 -1393 3378 -1378
tri 2988 -1457 3000 -1445 ne
rect 3000 -1450 3010 -1445
tri 3010 -1450 3015 -1445 sw
rect 2899 -1796 2914 -1568
rect 3000 -1606 3015 -1450
rect 3054 -1492 3082 -1436
tri 3174 -1454 3192 -1436 ne
rect 3192 -1456 3214 -1436
tri 3214 -1456 3234 -1436 sw
tri 3250 -1450 3268 -1432 ne
rect 3073 -1526 3082 -1492
rect 3116 -1465 3158 -1464
rect 3116 -1499 3121 -1465
rect 3151 -1499 3158 -1465
rect 3116 -1508 3158 -1499
rect 3192 -1465 3234 -1456
rect 3192 -1499 3199 -1465
rect 3229 -1499 3234 -1465
rect 3192 -1504 3234 -1499
rect 3268 -1492 3296 -1432
tri 3341 -1445 3363 -1423 se
rect 3363 -1430 3378 -1422
tri 3363 -1445 3378 -1430 nw
tri 3335 -1451 3341 -1445 se
rect 3341 -1451 3350 -1445
rect 3054 -1536 3082 -1526
tri 3082 -1536 3106 -1512 sw
rect 3054 -1568 3096 -1536
tri 3113 -1544 3114 -1543 sw
rect 3113 -1568 3114 -1544
tri 3116 -1545 3153 -1508 ne
rect 3153 -1536 3158 -1508
tri 3158 -1536 3184 -1510 sw
rect 3268 -1526 3277 -1492
rect 3268 -1536 3296 -1526
rect 3153 -1545 3237 -1536
tri 3153 -1564 3172 -1545 ne
rect 3172 -1564 3237 -1545
rect 3054 -1590 3114 -1568
rect 3236 -1568 3237 -1564
rect 3254 -1568 3296 -1536
rect 3236 -1590 3296 -1568
rect 3142 -1606 3159 -1592
rect 3191 -1606 3208 -1592
tri 2979 -1642 3001 -1620 se
rect 3001 -1627 3016 -1606
tri 3001 -1642 3016 -1627 nw
rect 3335 -1627 3350 -1451
tri 3350 -1458 3363 -1445 nw
rect 3436 -1526 3451 -1298
tri 2973 -1648 2979 -1642 se
rect 2979 -1648 2988 -1642
rect 2973 -1664 2988 -1648
tri 2988 -1655 3001 -1642 nw
rect 3142 -1650 3159 -1636
rect 3191 -1650 3208 -1636
tri 3335 -1642 3350 -1627 ne
tri 3350 -1642 3372 -1620 sw
rect 2973 -1700 2988 -1692
rect 3054 -1664 3114 -1650
rect 3069 -1674 3114 -1664
rect 3069 -1692 3097 -1674
tri 2973 -1715 2988 -1700 ne
tri 2988 -1715 3010 -1693 sw
rect 3054 -1702 3097 -1692
rect 3112 -1678 3114 -1674
rect 3236 -1664 3296 -1650
tri 3350 -1655 3363 -1642 ne
rect 3363 -1648 3372 -1642
tri 3372 -1648 3378 -1642 sw
rect 3236 -1674 3281 -1664
rect 3112 -1702 3186 -1678
rect 3054 -1706 3186 -1702
tri 3186 -1706 3214 -1678 sw
rect 3236 -1688 3238 -1674
tri 3236 -1690 3238 -1688 ne
rect 3250 -1692 3281 -1674
rect 3250 -1702 3296 -1692
rect 3363 -1663 3378 -1648
tri 2988 -1727 3000 -1715 ne
rect 3000 -1720 3010 -1715
tri 3010 -1720 3015 -1715 sw
rect 2899 -2066 2914 -1838
rect 3000 -1876 3015 -1720
rect 3054 -1762 3082 -1706
tri 3174 -1724 3192 -1706 ne
rect 3192 -1726 3214 -1706
tri 3214 -1726 3234 -1706 sw
tri 3250 -1720 3268 -1702 ne
rect 3073 -1796 3082 -1762
rect 3116 -1735 3158 -1734
rect 3116 -1769 3121 -1735
rect 3151 -1769 3158 -1735
rect 3116 -1778 3158 -1769
rect 3192 -1735 3234 -1726
rect 3192 -1769 3199 -1735
rect 3229 -1769 3234 -1735
rect 3192 -1774 3234 -1769
rect 3268 -1762 3296 -1702
tri 3341 -1715 3363 -1693 se
rect 3363 -1700 3378 -1692
tri 3363 -1715 3378 -1700 nw
tri 3335 -1721 3341 -1715 se
rect 3341 -1721 3350 -1715
rect 3054 -1806 3082 -1796
tri 3082 -1806 3106 -1782 sw
rect 3054 -1838 3096 -1806
tri 3113 -1814 3114 -1813 sw
rect 3113 -1838 3114 -1814
tri 3116 -1815 3153 -1778 ne
rect 3153 -1806 3158 -1778
tri 3158 -1806 3184 -1780 sw
rect 3268 -1796 3277 -1762
rect 3268 -1806 3296 -1796
rect 3153 -1815 3237 -1806
tri 3153 -1834 3172 -1815 ne
rect 3172 -1834 3237 -1815
rect 3054 -1860 3114 -1838
rect 3236 -1838 3237 -1834
rect 3254 -1838 3296 -1806
rect 3236 -1860 3296 -1838
rect 3142 -1876 3159 -1862
rect 3191 -1876 3208 -1862
tri 2979 -1912 3001 -1890 se
rect 3001 -1897 3016 -1876
tri 3001 -1912 3016 -1897 nw
rect 3335 -1897 3350 -1721
tri 3350 -1728 3363 -1715 nw
rect 3436 -1796 3451 -1568
tri 2973 -1918 2979 -1912 se
rect 2979 -1918 2988 -1912
rect 2973 -1934 2988 -1918
tri 2988 -1925 3001 -1912 nw
rect 3142 -1920 3159 -1906
rect 3191 -1920 3208 -1906
tri 3335 -1912 3350 -1897 ne
tri 3350 -1912 3372 -1890 sw
rect 2973 -1970 2988 -1962
rect 3054 -1934 3114 -1920
rect 3069 -1944 3114 -1934
rect 3069 -1962 3097 -1944
tri 2973 -1985 2988 -1970 ne
tri 2988 -1985 3010 -1963 sw
rect 3054 -1972 3097 -1962
rect 3112 -1948 3114 -1944
rect 3236 -1934 3296 -1920
tri 3350 -1925 3363 -1912 ne
rect 3363 -1918 3372 -1912
tri 3372 -1918 3378 -1912 sw
rect 3236 -1944 3281 -1934
rect 3112 -1972 3186 -1948
rect 3054 -1976 3186 -1972
tri 3186 -1976 3214 -1948 sw
rect 3236 -1958 3238 -1944
tri 3236 -1960 3238 -1958 ne
rect 3250 -1962 3281 -1944
rect 3250 -1972 3296 -1962
rect 3363 -1933 3378 -1918
tri 2988 -1997 3000 -1985 ne
rect 3000 -1990 3010 -1985
tri 3010 -1990 3015 -1985 sw
rect 2899 -2146 2914 -2108
rect 3000 -2146 3015 -1990
rect 3054 -2032 3082 -1976
tri 3174 -1994 3192 -1976 ne
rect 3192 -1996 3214 -1976
tri 3214 -1996 3234 -1976 sw
tri 3250 -1990 3268 -1972 ne
rect 3073 -2066 3082 -2032
rect 3116 -2005 3158 -2004
rect 3116 -2039 3121 -2005
rect 3151 -2039 3158 -2005
rect 3116 -2048 3158 -2039
rect 3192 -2005 3234 -1996
rect 3192 -2039 3199 -2005
rect 3229 -2039 3234 -2005
rect 3192 -2044 3234 -2039
rect 3268 -2032 3296 -1972
tri 3341 -1985 3363 -1963 se
rect 3363 -1970 3378 -1962
tri 3363 -1985 3378 -1970 nw
tri 3335 -1991 3341 -1985 se
rect 3341 -1991 3350 -1985
rect 3054 -2076 3082 -2066
tri 3082 -2076 3106 -2052 sw
rect 3054 -2108 3096 -2076
tri 3113 -2084 3114 -2083 sw
rect 3113 -2108 3114 -2084
tri 3116 -2085 3153 -2048 ne
rect 3153 -2076 3158 -2048
tri 3158 -2076 3184 -2050 sw
rect 3268 -2066 3277 -2032
rect 3268 -2076 3296 -2066
rect 3153 -2085 3237 -2076
tri 3153 -2104 3172 -2085 ne
rect 3172 -2104 3237 -2085
rect 3054 -2130 3114 -2108
rect 3236 -2108 3237 -2104
rect 3254 -2108 3296 -2076
rect 3236 -2130 3296 -2108
rect 3142 -2146 3159 -2132
rect 3191 -2146 3208 -2132
rect 3335 -2146 3350 -1991
tri 3350 -1998 3363 -1985 nw
rect 3436 -2066 3451 -1838
rect 3436 -2146 3451 -2108
rect 3479 1984 3494 2174
tri 3559 2138 3581 2160 se
rect 3581 2153 3596 2174
tri 3581 2138 3596 2153 nw
rect 3915 2153 3930 2174
tri 3553 2132 3559 2138 se
rect 3559 2132 3568 2138
rect 3553 2116 3568 2132
tri 3568 2125 3581 2138 nw
rect 3722 2130 3739 2144
rect 3771 2130 3788 2144
tri 3915 2138 3930 2153 ne
tri 3930 2138 3952 2160 sw
rect 3553 2080 3568 2088
rect 3634 2116 3694 2130
rect 3649 2106 3694 2116
rect 3649 2088 3677 2106
tri 3553 2065 3568 2080 ne
tri 3568 2065 3590 2087 sw
rect 3634 2078 3677 2088
rect 3692 2102 3694 2106
rect 3816 2116 3876 2130
tri 3930 2125 3943 2138 ne
rect 3943 2132 3952 2138
tri 3952 2132 3958 2138 sw
rect 3816 2106 3861 2116
rect 3692 2078 3766 2102
rect 3634 2074 3766 2078
tri 3766 2074 3794 2102 sw
rect 3816 2092 3818 2106
tri 3816 2090 3818 2092 ne
rect 3830 2088 3861 2106
rect 3830 2078 3876 2088
rect 3943 2117 3958 2132
tri 3568 2053 3580 2065 ne
rect 3580 2060 3590 2065
tri 3590 2060 3595 2065 sw
rect 3479 1714 3494 1942
rect 3580 1904 3595 2060
rect 3634 2018 3662 2074
tri 3754 2056 3772 2074 ne
rect 3772 2054 3794 2074
tri 3794 2054 3814 2074 sw
tri 3830 2060 3848 2078 ne
rect 3653 1984 3662 2018
rect 3696 2045 3738 2046
rect 3696 2011 3701 2045
rect 3731 2011 3738 2045
rect 3696 2002 3738 2011
rect 3772 2045 3814 2054
rect 3772 2011 3779 2045
rect 3809 2011 3814 2045
rect 3772 2006 3814 2011
rect 3848 2018 3876 2078
tri 3921 2065 3943 2087 se
rect 3943 2080 3958 2088
tri 3943 2065 3958 2080 nw
tri 3915 2059 3921 2065 se
rect 3921 2059 3930 2065
rect 3634 1974 3662 1984
tri 3662 1974 3686 1998 sw
rect 3634 1942 3676 1974
tri 3693 1966 3694 1967 sw
rect 3693 1942 3694 1966
tri 3696 1965 3733 2002 ne
rect 3733 1974 3738 2002
tri 3738 1974 3764 2000 sw
rect 3848 1984 3857 2018
rect 3848 1974 3876 1984
rect 3733 1965 3817 1974
tri 3733 1946 3752 1965 ne
rect 3752 1946 3817 1965
rect 3634 1920 3694 1942
rect 3816 1942 3817 1946
rect 3834 1942 3876 1974
rect 3816 1920 3876 1942
rect 3722 1904 3739 1918
rect 3771 1904 3788 1918
tri 3559 1868 3581 1890 se
rect 3581 1883 3596 1904
tri 3581 1868 3596 1883 nw
rect 3915 1883 3930 2059
tri 3930 2052 3943 2065 nw
rect 4016 1984 4031 2174
tri 3553 1862 3559 1868 se
rect 3559 1862 3568 1868
rect 3553 1846 3568 1862
tri 3568 1855 3581 1868 nw
rect 3722 1860 3739 1874
rect 3771 1860 3788 1874
tri 3915 1868 3930 1883 ne
tri 3930 1868 3952 1890 sw
rect 3553 1810 3568 1818
rect 3634 1846 3694 1860
rect 3649 1836 3694 1846
rect 3649 1818 3677 1836
tri 3553 1795 3568 1810 ne
tri 3568 1795 3590 1817 sw
rect 3634 1808 3677 1818
rect 3692 1832 3694 1836
rect 3816 1846 3876 1860
tri 3930 1855 3943 1868 ne
rect 3943 1862 3952 1868
tri 3952 1862 3958 1868 sw
rect 3816 1836 3861 1846
rect 3692 1808 3766 1832
rect 3634 1804 3766 1808
tri 3766 1804 3794 1832 sw
rect 3816 1822 3818 1836
tri 3816 1820 3818 1822 ne
rect 3830 1818 3861 1836
rect 3830 1808 3876 1818
rect 3943 1847 3958 1862
tri 3568 1783 3580 1795 ne
rect 3580 1790 3590 1795
tri 3590 1790 3595 1795 sw
rect 3479 1444 3494 1672
rect 3580 1634 3595 1790
rect 3634 1748 3662 1804
tri 3754 1786 3772 1804 ne
rect 3772 1784 3794 1804
tri 3794 1784 3814 1804 sw
tri 3830 1790 3848 1808 ne
rect 3653 1714 3662 1748
rect 3696 1775 3738 1776
rect 3696 1741 3701 1775
rect 3731 1741 3738 1775
rect 3696 1732 3738 1741
rect 3772 1775 3814 1784
rect 3772 1741 3779 1775
rect 3809 1741 3814 1775
rect 3772 1736 3814 1741
rect 3848 1748 3876 1808
tri 3921 1795 3943 1817 se
rect 3943 1810 3958 1818
tri 3943 1795 3958 1810 nw
tri 3915 1789 3921 1795 se
rect 3921 1789 3930 1795
rect 3634 1704 3662 1714
tri 3662 1704 3686 1728 sw
rect 3634 1672 3676 1704
tri 3693 1696 3694 1697 sw
rect 3693 1672 3694 1696
tri 3696 1695 3733 1732 ne
rect 3733 1704 3738 1732
tri 3738 1704 3764 1730 sw
rect 3848 1714 3857 1748
rect 3848 1704 3876 1714
rect 3733 1695 3817 1704
tri 3733 1676 3752 1695 ne
rect 3752 1676 3817 1695
rect 3634 1650 3694 1672
rect 3816 1672 3817 1676
rect 3834 1672 3876 1704
rect 3816 1650 3876 1672
rect 3722 1634 3739 1648
rect 3771 1634 3788 1648
tri 3559 1598 3581 1620 se
rect 3581 1613 3596 1634
tri 3581 1598 3596 1613 nw
rect 3915 1613 3930 1789
tri 3930 1782 3943 1795 nw
rect 4016 1714 4031 1942
tri 3553 1592 3559 1598 se
rect 3559 1592 3568 1598
rect 3553 1576 3568 1592
tri 3568 1585 3581 1598 nw
rect 3722 1590 3739 1604
rect 3771 1590 3788 1604
tri 3915 1598 3930 1613 ne
tri 3930 1598 3952 1620 sw
rect 3553 1540 3568 1548
rect 3634 1576 3694 1590
rect 3649 1566 3694 1576
rect 3649 1548 3677 1566
tri 3553 1525 3568 1540 ne
tri 3568 1525 3590 1547 sw
rect 3634 1538 3677 1548
rect 3692 1562 3694 1566
rect 3816 1576 3876 1590
tri 3930 1585 3943 1598 ne
rect 3943 1592 3952 1598
tri 3952 1592 3958 1598 sw
rect 3816 1566 3861 1576
rect 3692 1538 3766 1562
rect 3634 1534 3766 1538
tri 3766 1534 3794 1562 sw
rect 3816 1552 3818 1566
tri 3816 1550 3818 1552 ne
rect 3830 1548 3861 1566
rect 3830 1538 3876 1548
rect 3943 1577 3958 1592
tri 3568 1513 3580 1525 ne
rect 3580 1520 3590 1525
tri 3590 1520 3595 1525 sw
rect 3479 1174 3494 1402
rect 3580 1364 3595 1520
rect 3634 1478 3662 1534
tri 3754 1516 3772 1534 ne
rect 3772 1514 3794 1534
tri 3794 1514 3814 1534 sw
tri 3830 1520 3848 1538 ne
rect 3653 1444 3662 1478
rect 3696 1505 3738 1506
rect 3696 1471 3701 1505
rect 3731 1471 3738 1505
rect 3696 1462 3738 1471
rect 3772 1505 3814 1514
rect 3772 1471 3779 1505
rect 3809 1471 3814 1505
rect 3772 1466 3814 1471
rect 3848 1478 3876 1538
tri 3921 1525 3943 1547 se
rect 3943 1540 3958 1548
tri 3943 1525 3958 1540 nw
tri 3915 1519 3921 1525 se
rect 3921 1519 3930 1525
rect 3634 1434 3662 1444
tri 3662 1434 3686 1458 sw
rect 3634 1402 3676 1434
tri 3693 1426 3694 1427 sw
rect 3693 1402 3694 1426
tri 3696 1425 3733 1462 ne
rect 3733 1434 3738 1462
tri 3738 1434 3764 1460 sw
rect 3848 1444 3857 1478
rect 3848 1434 3876 1444
rect 3733 1425 3817 1434
tri 3733 1406 3752 1425 ne
rect 3752 1406 3817 1425
rect 3634 1380 3694 1402
rect 3816 1402 3817 1406
rect 3834 1402 3876 1434
rect 3816 1380 3876 1402
rect 3722 1364 3739 1378
rect 3771 1364 3788 1378
tri 3559 1328 3581 1350 se
rect 3581 1343 3596 1364
tri 3581 1328 3596 1343 nw
rect 3915 1343 3930 1519
tri 3930 1512 3943 1525 nw
rect 4016 1444 4031 1672
tri 3553 1322 3559 1328 se
rect 3559 1322 3568 1328
rect 3553 1306 3568 1322
tri 3568 1315 3581 1328 nw
rect 3722 1320 3739 1334
rect 3771 1320 3788 1334
tri 3915 1328 3930 1343 ne
tri 3930 1328 3952 1350 sw
rect 3553 1270 3568 1278
rect 3634 1306 3694 1320
rect 3649 1296 3694 1306
rect 3649 1278 3677 1296
tri 3553 1255 3568 1270 ne
tri 3568 1255 3590 1277 sw
rect 3634 1268 3677 1278
rect 3692 1292 3694 1296
rect 3816 1306 3876 1320
tri 3930 1315 3943 1328 ne
rect 3943 1322 3952 1328
tri 3952 1322 3958 1328 sw
rect 3816 1296 3861 1306
rect 3692 1268 3766 1292
rect 3634 1264 3766 1268
tri 3766 1264 3794 1292 sw
rect 3816 1282 3818 1296
tri 3816 1280 3818 1282 ne
rect 3830 1278 3861 1296
rect 3830 1268 3876 1278
rect 3943 1307 3958 1322
tri 3568 1243 3580 1255 ne
rect 3580 1250 3590 1255
tri 3590 1250 3595 1255 sw
rect 3479 904 3494 1132
rect 3580 1094 3595 1250
rect 3634 1208 3662 1264
tri 3754 1246 3772 1264 ne
rect 3772 1244 3794 1264
tri 3794 1244 3814 1264 sw
tri 3830 1250 3848 1268 ne
rect 3653 1174 3662 1208
rect 3696 1235 3738 1236
rect 3696 1201 3701 1235
rect 3731 1201 3738 1235
rect 3696 1192 3738 1201
rect 3772 1235 3814 1244
rect 3772 1201 3779 1235
rect 3809 1201 3814 1235
rect 3772 1196 3814 1201
rect 3848 1208 3876 1268
tri 3921 1255 3943 1277 se
rect 3943 1270 3958 1278
tri 3943 1255 3958 1270 nw
tri 3915 1249 3921 1255 se
rect 3921 1249 3930 1255
rect 3634 1164 3662 1174
tri 3662 1164 3686 1188 sw
rect 3634 1132 3676 1164
tri 3693 1156 3694 1157 sw
rect 3693 1132 3694 1156
tri 3696 1155 3733 1192 ne
rect 3733 1164 3738 1192
tri 3738 1164 3764 1190 sw
rect 3848 1174 3857 1208
rect 3848 1164 3876 1174
rect 3733 1155 3817 1164
tri 3733 1136 3752 1155 ne
rect 3752 1136 3817 1155
rect 3634 1110 3694 1132
rect 3816 1132 3817 1136
rect 3834 1132 3876 1164
rect 3816 1110 3876 1132
rect 3722 1094 3739 1108
rect 3771 1094 3788 1108
tri 3559 1058 3581 1080 se
rect 3581 1073 3596 1094
tri 3581 1058 3596 1073 nw
rect 3915 1073 3930 1249
tri 3930 1242 3943 1255 nw
rect 4016 1174 4031 1402
tri 3553 1052 3559 1058 se
rect 3559 1052 3568 1058
rect 3553 1036 3568 1052
tri 3568 1045 3581 1058 nw
rect 3722 1050 3739 1064
rect 3771 1050 3788 1064
tri 3915 1058 3930 1073 ne
tri 3930 1058 3952 1080 sw
rect 3553 1000 3568 1008
rect 3634 1036 3694 1050
rect 3649 1026 3694 1036
rect 3649 1008 3677 1026
tri 3553 985 3568 1000 ne
tri 3568 985 3590 1007 sw
rect 3634 998 3677 1008
rect 3692 1022 3694 1026
rect 3816 1036 3876 1050
tri 3930 1045 3943 1058 ne
rect 3943 1052 3952 1058
tri 3952 1052 3958 1058 sw
rect 3816 1026 3861 1036
rect 3692 998 3766 1022
rect 3634 994 3766 998
tri 3766 994 3794 1022 sw
rect 3816 1012 3818 1026
tri 3816 1010 3818 1012 ne
rect 3830 1008 3861 1026
rect 3830 998 3876 1008
rect 3943 1037 3958 1052
tri 3568 973 3580 985 ne
rect 3580 980 3590 985
tri 3590 980 3595 985 sw
rect 3479 634 3494 862
rect 3580 824 3595 980
rect 3634 938 3662 994
tri 3754 976 3772 994 ne
rect 3772 974 3794 994
tri 3794 974 3814 994 sw
tri 3830 980 3848 998 ne
rect 3653 904 3662 938
rect 3696 965 3738 966
rect 3696 931 3701 965
rect 3731 931 3738 965
rect 3696 922 3738 931
rect 3772 965 3814 974
rect 3772 931 3779 965
rect 3809 931 3814 965
rect 3772 926 3814 931
rect 3848 938 3876 998
tri 3921 985 3943 1007 se
rect 3943 1000 3958 1008
tri 3943 985 3958 1000 nw
tri 3915 979 3921 985 se
rect 3921 979 3930 985
rect 3634 894 3662 904
tri 3662 894 3686 918 sw
rect 3634 862 3676 894
tri 3693 886 3694 887 sw
rect 3693 862 3694 886
tri 3696 885 3733 922 ne
rect 3733 894 3738 922
tri 3738 894 3764 920 sw
rect 3848 904 3857 938
rect 3848 894 3876 904
rect 3733 885 3817 894
tri 3733 866 3752 885 ne
rect 3752 866 3817 885
rect 3634 840 3694 862
rect 3816 862 3817 866
rect 3834 862 3876 894
rect 3816 840 3876 862
rect 3722 824 3739 838
rect 3771 824 3788 838
tri 3559 788 3581 810 se
rect 3581 803 3596 824
tri 3581 788 3596 803 nw
rect 3915 803 3930 979
tri 3930 972 3943 985 nw
rect 4016 904 4031 1132
tri 3553 782 3559 788 se
rect 3559 782 3568 788
rect 3553 766 3568 782
tri 3568 775 3581 788 nw
rect 3722 780 3739 794
rect 3771 780 3788 794
tri 3915 788 3930 803 ne
tri 3930 788 3952 810 sw
rect 3553 730 3568 738
rect 3634 766 3694 780
rect 3649 756 3694 766
rect 3649 738 3677 756
tri 3553 715 3568 730 ne
tri 3568 715 3590 737 sw
rect 3634 728 3677 738
rect 3692 752 3694 756
rect 3816 766 3876 780
tri 3930 775 3943 788 ne
rect 3943 782 3952 788
tri 3952 782 3958 788 sw
rect 3816 756 3861 766
rect 3692 728 3766 752
rect 3634 724 3766 728
tri 3766 724 3794 752 sw
rect 3816 742 3818 756
tri 3816 740 3818 742 ne
rect 3830 738 3861 756
rect 3830 728 3876 738
rect 3943 767 3958 782
tri 3568 703 3580 715 ne
rect 3580 710 3590 715
tri 3590 710 3595 715 sw
rect 3479 364 3494 592
rect 3580 554 3595 710
rect 3634 668 3662 724
tri 3754 706 3772 724 ne
rect 3772 704 3794 724
tri 3794 704 3814 724 sw
tri 3830 710 3848 728 ne
rect 3653 634 3662 668
rect 3696 695 3738 696
rect 3696 661 3701 695
rect 3731 661 3738 695
rect 3696 652 3738 661
rect 3772 695 3814 704
rect 3772 661 3779 695
rect 3809 661 3814 695
rect 3772 656 3814 661
rect 3848 668 3876 728
tri 3921 715 3943 737 se
rect 3943 730 3958 738
tri 3943 715 3958 730 nw
tri 3915 709 3921 715 se
rect 3921 709 3930 715
rect 3634 624 3662 634
tri 3662 624 3686 648 sw
rect 3634 592 3676 624
tri 3693 616 3694 617 sw
rect 3693 592 3694 616
tri 3696 615 3733 652 ne
rect 3733 624 3738 652
tri 3738 624 3764 650 sw
rect 3848 634 3857 668
rect 3848 624 3876 634
rect 3733 615 3817 624
tri 3733 596 3752 615 ne
rect 3752 596 3817 615
rect 3634 570 3694 592
rect 3816 592 3817 596
rect 3834 592 3876 624
rect 3816 570 3876 592
rect 3722 554 3739 568
rect 3771 554 3788 568
tri 3559 518 3581 540 se
rect 3581 533 3596 554
tri 3581 518 3596 533 nw
rect 3915 533 3930 709
tri 3930 702 3943 715 nw
rect 4016 634 4031 862
tri 3553 512 3559 518 se
rect 3559 512 3568 518
rect 3553 496 3568 512
tri 3568 505 3581 518 nw
rect 3722 510 3739 524
rect 3771 510 3788 524
tri 3915 518 3930 533 ne
tri 3930 518 3952 540 sw
rect 3553 460 3568 468
rect 3634 496 3694 510
rect 3649 486 3694 496
rect 3649 468 3677 486
tri 3553 445 3568 460 ne
tri 3568 445 3590 467 sw
rect 3634 458 3677 468
rect 3692 482 3694 486
rect 3816 496 3876 510
tri 3930 505 3943 518 ne
rect 3943 512 3952 518
tri 3952 512 3958 518 sw
rect 3816 486 3861 496
rect 3692 458 3766 482
rect 3634 454 3766 458
tri 3766 454 3794 482 sw
rect 3816 472 3818 486
tri 3816 470 3818 472 ne
rect 3830 468 3861 486
rect 3830 458 3876 468
rect 3943 497 3958 512
tri 3568 433 3580 445 ne
rect 3580 440 3590 445
tri 3590 440 3595 445 sw
rect 3479 94 3494 322
rect 3580 284 3595 440
rect 3634 398 3662 454
tri 3754 436 3772 454 ne
rect 3772 434 3794 454
tri 3794 434 3814 454 sw
tri 3830 440 3848 458 ne
rect 3653 364 3662 398
rect 3696 425 3738 426
rect 3696 391 3701 425
rect 3731 391 3738 425
rect 3696 382 3738 391
rect 3772 425 3814 434
rect 3772 391 3779 425
rect 3809 391 3814 425
rect 3772 386 3814 391
rect 3848 398 3876 458
tri 3921 445 3943 467 se
rect 3943 460 3958 468
tri 3943 445 3958 460 nw
tri 3915 439 3921 445 se
rect 3921 439 3930 445
rect 3634 354 3662 364
tri 3662 354 3686 378 sw
rect 3634 322 3676 354
tri 3693 346 3694 347 sw
rect 3693 322 3694 346
tri 3696 345 3733 382 ne
rect 3733 354 3738 382
tri 3738 354 3764 380 sw
rect 3848 364 3857 398
rect 3848 354 3876 364
rect 3733 345 3817 354
tri 3733 326 3752 345 ne
rect 3752 326 3817 345
rect 3634 300 3694 322
rect 3816 322 3817 326
rect 3834 322 3876 354
rect 3816 300 3876 322
rect 3722 284 3739 298
rect 3771 284 3788 298
tri 3559 248 3581 270 se
rect 3581 263 3596 284
tri 3581 248 3596 263 nw
rect 3915 263 3930 439
tri 3930 432 3943 445 nw
rect 4016 364 4031 592
tri 3553 242 3559 248 se
rect 3559 242 3568 248
rect 3553 226 3568 242
tri 3568 235 3581 248 nw
rect 3722 240 3739 254
rect 3771 240 3788 254
tri 3915 248 3930 263 ne
tri 3930 248 3952 270 sw
rect 3553 190 3568 198
rect 3634 226 3694 240
rect 3649 216 3694 226
rect 3649 198 3677 216
tri 3553 175 3568 190 ne
tri 3568 175 3590 197 sw
rect 3634 188 3677 198
rect 3692 212 3694 216
rect 3816 226 3876 240
tri 3930 235 3943 248 ne
rect 3943 242 3952 248
tri 3952 242 3958 248 sw
rect 3816 216 3861 226
rect 3692 188 3766 212
rect 3634 184 3766 188
tri 3766 184 3794 212 sw
rect 3816 202 3818 216
tri 3816 200 3818 202 ne
rect 3830 198 3861 216
rect 3830 188 3876 198
rect 3943 227 3958 242
tri 3568 163 3580 175 ne
rect 3580 170 3590 175
tri 3590 170 3595 175 sw
rect 3479 -176 3494 52
rect 3580 14 3595 170
rect 3634 128 3662 184
tri 3754 166 3772 184 ne
rect 3772 164 3794 184
tri 3794 164 3814 184 sw
tri 3830 170 3848 188 ne
rect 3653 94 3662 128
rect 3696 155 3738 156
rect 3696 121 3701 155
rect 3731 121 3738 155
rect 3696 112 3738 121
rect 3772 155 3814 164
rect 3772 121 3779 155
rect 3809 121 3814 155
rect 3772 116 3814 121
rect 3848 128 3876 188
tri 3921 175 3943 197 se
rect 3943 190 3958 198
tri 3943 175 3958 190 nw
tri 3915 169 3921 175 se
rect 3921 169 3930 175
rect 3634 84 3662 94
tri 3662 84 3686 108 sw
rect 3634 52 3676 84
tri 3693 76 3694 77 sw
rect 3693 52 3694 76
tri 3696 75 3733 112 ne
rect 3733 84 3738 112
tri 3738 84 3764 110 sw
rect 3848 94 3857 128
rect 3848 84 3876 94
rect 3733 75 3817 84
tri 3733 56 3752 75 ne
rect 3752 56 3817 75
rect 3634 30 3694 52
rect 3816 52 3817 56
rect 3834 52 3876 84
rect 3816 30 3876 52
rect 3722 14 3739 28
rect 3771 14 3788 28
tri 3559 -22 3581 0 se
rect 3581 -7 3596 14
tri 3581 -22 3596 -7 nw
rect 3915 -7 3930 169
tri 3930 162 3943 175 nw
rect 4016 94 4031 322
tri 3553 -28 3559 -22 se
rect 3559 -28 3568 -22
rect 3553 -44 3568 -28
tri 3568 -35 3581 -22 nw
rect 3722 -30 3739 -16
rect 3771 -30 3788 -16
tri 3915 -22 3930 -7 ne
tri 3930 -22 3952 0 sw
rect 3553 -80 3568 -72
rect 3634 -44 3694 -30
rect 3649 -54 3694 -44
rect 3649 -72 3677 -54
tri 3553 -95 3568 -80 ne
tri 3568 -95 3590 -73 sw
rect 3634 -82 3677 -72
rect 3692 -58 3694 -54
rect 3816 -44 3876 -30
tri 3930 -35 3943 -22 ne
rect 3943 -28 3952 -22
tri 3952 -28 3958 -22 sw
rect 3816 -54 3861 -44
rect 3692 -82 3766 -58
rect 3634 -86 3766 -82
tri 3766 -86 3794 -58 sw
rect 3816 -68 3818 -54
tri 3816 -70 3818 -68 ne
rect 3830 -72 3861 -54
rect 3830 -82 3876 -72
rect 3943 -43 3958 -28
tri 3568 -107 3580 -95 ne
rect 3580 -100 3590 -95
tri 3590 -100 3595 -95 sw
rect 3479 -446 3494 -218
rect 3580 -256 3595 -100
rect 3634 -142 3662 -86
tri 3754 -104 3772 -86 ne
rect 3772 -106 3794 -86
tri 3794 -106 3814 -86 sw
tri 3830 -100 3848 -82 ne
rect 3653 -176 3662 -142
rect 3696 -115 3738 -114
rect 3696 -149 3701 -115
rect 3731 -149 3738 -115
rect 3696 -158 3738 -149
rect 3772 -115 3814 -106
rect 3772 -149 3779 -115
rect 3809 -149 3814 -115
rect 3772 -154 3814 -149
rect 3848 -142 3876 -82
tri 3921 -95 3943 -73 se
rect 3943 -80 3958 -72
tri 3943 -95 3958 -80 nw
tri 3915 -101 3921 -95 se
rect 3921 -101 3930 -95
rect 3634 -186 3662 -176
tri 3662 -186 3686 -162 sw
rect 3634 -218 3676 -186
tri 3693 -194 3694 -193 sw
rect 3693 -218 3694 -194
tri 3696 -195 3733 -158 ne
rect 3733 -186 3738 -158
tri 3738 -186 3764 -160 sw
rect 3848 -176 3857 -142
rect 3848 -186 3876 -176
rect 3733 -195 3817 -186
tri 3733 -214 3752 -195 ne
rect 3752 -214 3817 -195
rect 3634 -240 3694 -218
rect 3816 -218 3817 -214
rect 3834 -218 3876 -186
rect 3816 -240 3876 -218
rect 3722 -256 3739 -242
rect 3771 -256 3788 -242
tri 3559 -292 3581 -270 se
rect 3581 -277 3596 -256
tri 3581 -292 3596 -277 nw
rect 3915 -277 3930 -101
tri 3930 -108 3943 -95 nw
rect 4016 -176 4031 52
tri 3553 -298 3559 -292 se
rect 3559 -298 3568 -292
rect 3553 -314 3568 -298
tri 3568 -305 3581 -292 nw
rect 3722 -300 3739 -286
rect 3771 -300 3788 -286
tri 3915 -292 3930 -277 ne
tri 3930 -292 3952 -270 sw
rect 3553 -350 3568 -342
rect 3634 -314 3694 -300
rect 3649 -324 3694 -314
rect 3649 -342 3677 -324
tri 3553 -365 3568 -350 ne
tri 3568 -365 3590 -343 sw
rect 3634 -352 3677 -342
rect 3692 -328 3694 -324
rect 3816 -314 3876 -300
tri 3930 -305 3943 -292 ne
rect 3943 -298 3952 -292
tri 3952 -298 3958 -292 sw
rect 3816 -324 3861 -314
rect 3692 -352 3766 -328
rect 3634 -356 3766 -352
tri 3766 -356 3794 -328 sw
rect 3816 -338 3818 -324
tri 3816 -340 3818 -338 ne
rect 3830 -342 3861 -324
rect 3830 -352 3876 -342
rect 3943 -313 3958 -298
tri 3568 -377 3580 -365 ne
rect 3580 -370 3590 -365
tri 3590 -370 3595 -365 sw
rect 3479 -716 3494 -488
rect 3580 -526 3595 -370
rect 3634 -412 3662 -356
tri 3754 -374 3772 -356 ne
rect 3772 -376 3794 -356
tri 3794 -376 3814 -356 sw
tri 3830 -370 3848 -352 ne
rect 3653 -446 3662 -412
rect 3696 -385 3738 -384
rect 3696 -419 3701 -385
rect 3731 -419 3738 -385
rect 3696 -428 3738 -419
rect 3772 -385 3814 -376
rect 3772 -419 3779 -385
rect 3809 -419 3814 -385
rect 3772 -424 3814 -419
rect 3848 -412 3876 -352
tri 3921 -365 3943 -343 se
rect 3943 -350 3958 -342
tri 3943 -365 3958 -350 nw
tri 3915 -371 3921 -365 se
rect 3921 -371 3930 -365
rect 3634 -456 3662 -446
tri 3662 -456 3686 -432 sw
rect 3634 -488 3676 -456
tri 3693 -464 3694 -463 sw
rect 3693 -488 3694 -464
tri 3696 -465 3733 -428 ne
rect 3733 -456 3738 -428
tri 3738 -456 3764 -430 sw
rect 3848 -446 3857 -412
rect 3848 -456 3876 -446
rect 3733 -465 3817 -456
tri 3733 -484 3752 -465 ne
rect 3752 -484 3817 -465
rect 3634 -510 3694 -488
rect 3816 -488 3817 -484
rect 3834 -488 3876 -456
rect 3816 -510 3876 -488
rect 3722 -526 3739 -512
rect 3771 -526 3788 -512
tri 3559 -562 3581 -540 se
rect 3581 -547 3596 -526
tri 3581 -562 3596 -547 nw
rect 3915 -547 3930 -371
tri 3930 -378 3943 -365 nw
rect 4016 -446 4031 -218
tri 3553 -568 3559 -562 se
rect 3559 -568 3568 -562
rect 3553 -584 3568 -568
tri 3568 -575 3581 -562 nw
rect 3722 -570 3739 -556
rect 3771 -570 3788 -556
tri 3915 -562 3930 -547 ne
tri 3930 -562 3952 -540 sw
rect 3553 -620 3568 -612
rect 3634 -584 3694 -570
rect 3649 -594 3694 -584
rect 3649 -612 3677 -594
tri 3553 -635 3568 -620 ne
tri 3568 -635 3590 -613 sw
rect 3634 -622 3677 -612
rect 3692 -598 3694 -594
rect 3816 -584 3876 -570
tri 3930 -575 3943 -562 ne
rect 3943 -568 3952 -562
tri 3952 -568 3958 -562 sw
rect 3816 -594 3861 -584
rect 3692 -622 3766 -598
rect 3634 -626 3766 -622
tri 3766 -626 3794 -598 sw
rect 3816 -608 3818 -594
tri 3816 -610 3818 -608 ne
rect 3830 -612 3861 -594
rect 3830 -622 3876 -612
rect 3943 -583 3958 -568
tri 3568 -647 3580 -635 ne
rect 3580 -640 3590 -635
tri 3590 -640 3595 -635 sw
rect 3479 -986 3494 -758
rect 3580 -796 3595 -640
rect 3634 -682 3662 -626
tri 3754 -644 3772 -626 ne
rect 3772 -646 3794 -626
tri 3794 -646 3814 -626 sw
tri 3830 -640 3848 -622 ne
rect 3653 -716 3662 -682
rect 3696 -655 3738 -654
rect 3696 -689 3701 -655
rect 3731 -689 3738 -655
rect 3696 -698 3738 -689
rect 3772 -655 3814 -646
rect 3772 -689 3779 -655
rect 3809 -689 3814 -655
rect 3772 -694 3814 -689
rect 3848 -682 3876 -622
tri 3921 -635 3943 -613 se
rect 3943 -620 3958 -612
tri 3943 -635 3958 -620 nw
tri 3915 -641 3921 -635 se
rect 3921 -641 3930 -635
rect 3634 -726 3662 -716
tri 3662 -726 3686 -702 sw
rect 3634 -758 3676 -726
tri 3693 -734 3694 -733 sw
rect 3693 -758 3694 -734
tri 3696 -735 3733 -698 ne
rect 3733 -726 3738 -698
tri 3738 -726 3764 -700 sw
rect 3848 -716 3857 -682
rect 3848 -726 3876 -716
rect 3733 -735 3817 -726
tri 3733 -754 3752 -735 ne
rect 3752 -754 3817 -735
rect 3634 -780 3694 -758
rect 3816 -758 3817 -754
rect 3834 -758 3876 -726
rect 3816 -780 3876 -758
rect 3722 -796 3739 -782
rect 3771 -796 3788 -782
tri 3559 -832 3581 -810 se
rect 3581 -817 3596 -796
tri 3581 -832 3596 -817 nw
rect 3915 -817 3930 -641
tri 3930 -648 3943 -635 nw
rect 4016 -716 4031 -488
tri 3553 -838 3559 -832 se
rect 3559 -838 3568 -832
rect 3553 -854 3568 -838
tri 3568 -845 3581 -832 nw
rect 3722 -840 3739 -826
rect 3771 -840 3788 -826
tri 3915 -832 3930 -817 ne
tri 3930 -832 3952 -810 sw
rect 3553 -890 3568 -882
rect 3634 -854 3694 -840
rect 3649 -864 3694 -854
rect 3649 -882 3677 -864
tri 3553 -905 3568 -890 ne
tri 3568 -905 3590 -883 sw
rect 3634 -892 3677 -882
rect 3692 -868 3694 -864
rect 3816 -854 3876 -840
tri 3930 -845 3943 -832 ne
rect 3943 -838 3952 -832
tri 3952 -838 3958 -832 sw
rect 3816 -864 3861 -854
rect 3692 -892 3766 -868
rect 3634 -896 3766 -892
tri 3766 -896 3794 -868 sw
rect 3816 -878 3818 -864
tri 3816 -880 3818 -878 ne
rect 3830 -882 3861 -864
rect 3830 -892 3876 -882
rect 3943 -853 3958 -838
tri 3568 -917 3580 -905 ne
rect 3580 -910 3590 -905
tri 3590 -910 3595 -905 sw
rect 3479 -1256 3494 -1028
rect 3580 -1066 3595 -910
rect 3634 -952 3662 -896
tri 3754 -914 3772 -896 ne
rect 3772 -916 3794 -896
tri 3794 -916 3814 -896 sw
tri 3830 -910 3848 -892 ne
rect 3653 -986 3662 -952
rect 3696 -925 3738 -924
rect 3696 -959 3701 -925
rect 3731 -959 3738 -925
rect 3696 -968 3738 -959
rect 3772 -925 3814 -916
rect 3772 -959 3779 -925
rect 3809 -959 3814 -925
rect 3772 -964 3814 -959
rect 3848 -952 3876 -892
tri 3921 -905 3943 -883 se
rect 3943 -890 3958 -882
tri 3943 -905 3958 -890 nw
tri 3915 -911 3921 -905 se
rect 3921 -911 3930 -905
rect 3634 -996 3662 -986
tri 3662 -996 3686 -972 sw
rect 3634 -1028 3676 -996
tri 3693 -1004 3694 -1003 sw
rect 3693 -1028 3694 -1004
tri 3696 -1005 3733 -968 ne
rect 3733 -996 3738 -968
tri 3738 -996 3764 -970 sw
rect 3848 -986 3857 -952
rect 3848 -996 3876 -986
rect 3733 -1005 3817 -996
tri 3733 -1024 3752 -1005 ne
rect 3752 -1024 3817 -1005
rect 3634 -1050 3694 -1028
rect 3816 -1028 3817 -1024
rect 3834 -1028 3876 -996
rect 3816 -1050 3876 -1028
rect 3722 -1066 3739 -1052
rect 3771 -1066 3788 -1052
tri 3559 -1102 3581 -1080 se
rect 3581 -1087 3596 -1066
tri 3581 -1102 3596 -1087 nw
rect 3915 -1087 3930 -911
tri 3930 -918 3943 -905 nw
rect 4016 -986 4031 -758
tri 3553 -1108 3559 -1102 se
rect 3559 -1108 3568 -1102
rect 3553 -1124 3568 -1108
tri 3568 -1115 3581 -1102 nw
rect 3722 -1110 3739 -1096
rect 3771 -1110 3788 -1096
tri 3915 -1102 3930 -1087 ne
tri 3930 -1102 3952 -1080 sw
rect 3553 -1160 3568 -1152
rect 3634 -1124 3694 -1110
rect 3649 -1134 3694 -1124
rect 3649 -1152 3677 -1134
tri 3553 -1175 3568 -1160 ne
tri 3568 -1175 3590 -1153 sw
rect 3634 -1162 3677 -1152
rect 3692 -1138 3694 -1134
rect 3816 -1124 3876 -1110
tri 3930 -1115 3943 -1102 ne
rect 3943 -1108 3952 -1102
tri 3952 -1108 3958 -1102 sw
rect 3816 -1134 3861 -1124
rect 3692 -1162 3766 -1138
rect 3634 -1166 3766 -1162
tri 3766 -1166 3794 -1138 sw
rect 3816 -1148 3818 -1134
tri 3816 -1150 3818 -1148 ne
rect 3830 -1152 3861 -1134
rect 3830 -1162 3876 -1152
rect 3943 -1123 3958 -1108
tri 3568 -1187 3580 -1175 ne
rect 3580 -1180 3590 -1175
tri 3590 -1180 3595 -1175 sw
rect 3479 -1526 3494 -1298
rect 3580 -1336 3595 -1180
rect 3634 -1222 3662 -1166
tri 3754 -1184 3772 -1166 ne
rect 3772 -1186 3794 -1166
tri 3794 -1186 3814 -1166 sw
tri 3830 -1180 3848 -1162 ne
rect 3653 -1256 3662 -1222
rect 3696 -1195 3738 -1194
rect 3696 -1229 3701 -1195
rect 3731 -1229 3738 -1195
rect 3696 -1238 3738 -1229
rect 3772 -1195 3814 -1186
rect 3772 -1229 3779 -1195
rect 3809 -1229 3814 -1195
rect 3772 -1234 3814 -1229
rect 3848 -1222 3876 -1162
tri 3921 -1175 3943 -1153 se
rect 3943 -1160 3958 -1152
tri 3943 -1175 3958 -1160 nw
tri 3915 -1181 3921 -1175 se
rect 3921 -1181 3930 -1175
rect 3634 -1266 3662 -1256
tri 3662 -1266 3686 -1242 sw
rect 3634 -1298 3676 -1266
tri 3693 -1274 3694 -1273 sw
rect 3693 -1298 3694 -1274
tri 3696 -1275 3733 -1238 ne
rect 3733 -1266 3738 -1238
tri 3738 -1266 3764 -1240 sw
rect 3848 -1256 3857 -1222
rect 3848 -1266 3876 -1256
rect 3733 -1275 3817 -1266
tri 3733 -1294 3752 -1275 ne
rect 3752 -1294 3817 -1275
rect 3634 -1320 3694 -1298
rect 3816 -1298 3817 -1294
rect 3834 -1298 3876 -1266
rect 3816 -1320 3876 -1298
rect 3722 -1336 3739 -1322
rect 3771 -1336 3788 -1322
tri 3559 -1372 3581 -1350 se
rect 3581 -1357 3596 -1336
tri 3581 -1372 3596 -1357 nw
rect 3915 -1357 3930 -1181
tri 3930 -1188 3943 -1175 nw
rect 4016 -1256 4031 -1028
tri 3553 -1378 3559 -1372 se
rect 3559 -1378 3568 -1372
rect 3553 -1394 3568 -1378
tri 3568 -1385 3581 -1372 nw
rect 3722 -1380 3739 -1366
rect 3771 -1380 3788 -1366
tri 3915 -1372 3930 -1357 ne
tri 3930 -1372 3952 -1350 sw
rect 3553 -1430 3568 -1422
rect 3634 -1394 3694 -1380
rect 3649 -1404 3694 -1394
rect 3649 -1422 3677 -1404
tri 3553 -1445 3568 -1430 ne
tri 3568 -1445 3590 -1423 sw
rect 3634 -1432 3677 -1422
rect 3692 -1408 3694 -1404
rect 3816 -1394 3876 -1380
tri 3930 -1385 3943 -1372 ne
rect 3943 -1378 3952 -1372
tri 3952 -1378 3958 -1372 sw
rect 3816 -1404 3861 -1394
rect 3692 -1432 3766 -1408
rect 3634 -1436 3766 -1432
tri 3766 -1436 3794 -1408 sw
rect 3816 -1418 3818 -1404
tri 3816 -1420 3818 -1418 ne
rect 3830 -1422 3861 -1404
rect 3830 -1432 3876 -1422
rect 3943 -1393 3958 -1378
tri 3568 -1457 3580 -1445 ne
rect 3580 -1450 3590 -1445
tri 3590 -1450 3595 -1445 sw
rect 3479 -1796 3494 -1568
rect 3580 -1606 3595 -1450
rect 3634 -1492 3662 -1436
tri 3754 -1454 3772 -1436 ne
rect 3772 -1456 3794 -1436
tri 3794 -1456 3814 -1436 sw
tri 3830 -1450 3848 -1432 ne
rect 3653 -1526 3662 -1492
rect 3696 -1465 3738 -1464
rect 3696 -1499 3701 -1465
rect 3731 -1499 3738 -1465
rect 3696 -1508 3738 -1499
rect 3772 -1465 3814 -1456
rect 3772 -1499 3779 -1465
rect 3809 -1499 3814 -1465
rect 3772 -1504 3814 -1499
rect 3848 -1492 3876 -1432
tri 3921 -1445 3943 -1423 se
rect 3943 -1430 3958 -1422
tri 3943 -1445 3958 -1430 nw
tri 3915 -1451 3921 -1445 se
rect 3921 -1451 3930 -1445
rect 3634 -1536 3662 -1526
tri 3662 -1536 3686 -1512 sw
rect 3634 -1568 3676 -1536
tri 3693 -1544 3694 -1543 sw
rect 3693 -1568 3694 -1544
tri 3696 -1545 3733 -1508 ne
rect 3733 -1536 3738 -1508
tri 3738 -1536 3764 -1510 sw
rect 3848 -1526 3857 -1492
rect 3848 -1536 3876 -1526
rect 3733 -1545 3817 -1536
tri 3733 -1564 3752 -1545 ne
rect 3752 -1564 3817 -1545
rect 3634 -1590 3694 -1568
rect 3816 -1568 3817 -1564
rect 3834 -1568 3876 -1536
rect 3816 -1590 3876 -1568
rect 3722 -1606 3739 -1592
rect 3771 -1606 3788 -1592
tri 3559 -1642 3581 -1620 se
rect 3581 -1627 3596 -1606
tri 3581 -1642 3596 -1627 nw
rect 3915 -1627 3930 -1451
tri 3930 -1458 3943 -1445 nw
rect 4016 -1526 4031 -1298
tri 3553 -1648 3559 -1642 se
rect 3559 -1648 3568 -1642
rect 3553 -1664 3568 -1648
tri 3568 -1655 3581 -1642 nw
rect 3722 -1650 3739 -1636
rect 3771 -1650 3788 -1636
tri 3915 -1642 3930 -1627 ne
tri 3930 -1642 3952 -1620 sw
rect 3553 -1700 3568 -1692
rect 3634 -1664 3694 -1650
rect 3649 -1674 3694 -1664
rect 3649 -1692 3677 -1674
tri 3553 -1715 3568 -1700 ne
tri 3568 -1715 3590 -1693 sw
rect 3634 -1702 3677 -1692
rect 3692 -1678 3694 -1674
rect 3816 -1664 3876 -1650
tri 3930 -1655 3943 -1642 ne
rect 3943 -1648 3952 -1642
tri 3952 -1648 3958 -1642 sw
rect 3816 -1674 3861 -1664
rect 3692 -1702 3766 -1678
rect 3634 -1706 3766 -1702
tri 3766 -1706 3794 -1678 sw
rect 3816 -1688 3818 -1674
tri 3816 -1690 3818 -1688 ne
rect 3830 -1692 3861 -1674
rect 3830 -1702 3876 -1692
rect 3943 -1663 3958 -1648
tri 3568 -1727 3580 -1715 ne
rect 3580 -1720 3590 -1715
tri 3590 -1720 3595 -1715 sw
rect 3479 -2066 3494 -1838
rect 3580 -1876 3595 -1720
rect 3634 -1762 3662 -1706
tri 3754 -1724 3772 -1706 ne
rect 3772 -1726 3794 -1706
tri 3794 -1726 3814 -1706 sw
tri 3830 -1720 3848 -1702 ne
rect 3653 -1796 3662 -1762
rect 3696 -1735 3738 -1734
rect 3696 -1769 3701 -1735
rect 3731 -1769 3738 -1735
rect 3696 -1778 3738 -1769
rect 3772 -1735 3814 -1726
rect 3772 -1769 3779 -1735
rect 3809 -1769 3814 -1735
rect 3772 -1774 3814 -1769
rect 3848 -1762 3876 -1702
tri 3921 -1715 3943 -1693 se
rect 3943 -1700 3958 -1692
tri 3943 -1715 3958 -1700 nw
tri 3915 -1721 3921 -1715 se
rect 3921 -1721 3930 -1715
rect 3634 -1806 3662 -1796
tri 3662 -1806 3686 -1782 sw
rect 3634 -1838 3676 -1806
tri 3693 -1814 3694 -1813 sw
rect 3693 -1838 3694 -1814
tri 3696 -1815 3733 -1778 ne
rect 3733 -1806 3738 -1778
tri 3738 -1806 3764 -1780 sw
rect 3848 -1796 3857 -1762
rect 3848 -1806 3876 -1796
rect 3733 -1815 3817 -1806
tri 3733 -1834 3752 -1815 ne
rect 3752 -1834 3817 -1815
rect 3634 -1860 3694 -1838
rect 3816 -1838 3817 -1834
rect 3834 -1838 3876 -1806
rect 3816 -1860 3876 -1838
rect 3722 -1876 3739 -1862
rect 3771 -1876 3788 -1862
tri 3559 -1912 3581 -1890 se
rect 3581 -1897 3596 -1876
tri 3581 -1912 3596 -1897 nw
rect 3915 -1897 3930 -1721
tri 3930 -1728 3943 -1715 nw
rect 4016 -1796 4031 -1568
tri 3553 -1918 3559 -1912 se
rect 3559 -1918 3568 -1912
rect 3553 -1934 3568 -1918
tri 3568 -1925 3581 -1912 nw
rect 3722 -1920 3739 -1906
rect 3771 -1920 3788 -1906
tri 3915 -1912 3930 -1897 ne
tri 3930 -1912 3952 -1890 sw
rect 3553 -1970 3568 -1962
rect 3634 -1934 3694 -1920
rect 3649 -1944 3694 -1934
rect 3649 -1962 3677 -1944
tri 3553 -1985 3568 -1970 ne
tri 3568 -1985 3590 -1963 sw
rect 3634 -1972 3677 -1962
rect 3692 -1948 3694 -1944
rect 3816 -1934 3876 -1920
tri 3930 -1925 3943 -1912 ne
rect 3943 -1918 3952 -1912
tri 3952 -1918 3958 -1912 sw
rect 3816 -1944 3861 -1934
rect 3692 -1972 3766 -1948
rect 3634 -1976 3766 -1972
tri 3766 -1976 3794 -1948 sw
rect 3816 -1958 3818 -1944
tri 3816 -1960 3818 -1958 ne
rect 3830 -1962 3861 -1944
rect 3830 -1972 3876 -1962
rect 3943 -1933 3958 -1918
tri 3568 -1997 3580 -1985 ne
rect 3580 -1990 3590 -1985
tri 3590 -1990 3595 -1985 sw
rect 3479 -2146 3494 -2108
rect 3580 -2146 3595 -1990
rect 3634 -2032 3662 -1976
tri 3754 -1994 3772 -1976 ne
rect 3772 -1996 3794 -1976
tri 3794 -1996 3814 -1976 sw
tri 3830 -1990 3848 -1972 ne
rect 3653 -2066 3662 -2032
rect 3696 -2005 3738 -2004
rect 3696 -2039 3701 -2005
rect 3731 -2039 3738 -2005
rect 3696 -2048 3738 -2039
rect 3772 -2005 3814 -1996
rect 3772 -2039 3779 -2005
rect 3809 -2039 3814 -2005
rect 3772 -2044 3814 -2039
rect 3848 -2032 3876 -1972
tri 3921 -1985 3943 -1963 se
rect 3943 -1970 3958 -1962
tri 3943 -1985 3958 -1970 nw
tri 3915 -1991 3921 -1985 se
rect 3921 -1991 3930 -1985
rect 3634 -2076 3662 -2066
tri 3662 -2076 3686 -2052 sw
rect 3634 -2108 3676 -2076
tri 3693 -2084 3694 -2083 sw
rect 3693 -2108 3694 -2084
tri 3696 -2085 3733 -2048 ne
rect 3733 -2076 3738 -2048
tri 3738 -2076 3764 -2050 sw
rect 3848 -2066 3857 -2032
rect 3848 -2076 3876 -2066
rect 3733 -2085 3817 -2076
tri 3733 -2104 3752 -2085 ne
rect 3752 -2104 3817 -2085
rect 3634 -2130 3694 -2108
rect 3816 -2108 3817 -2104
rect 3834 -2108 3876 -2076
rect 3816 -2130 3876 -2108
rect 3722 -2146 3739 -2132
rect 3771 -2146 3788 -2132
rect 3915 -2146 3930 -1991
tri 3930 -1998 3943 -1985 nw
rect 4016 -2066 4031 -1838
rect 4016 -2146 4031 -2108
rect 4059 1984 4074 2174
tri 4139 2138 4161 2160 se
rect 4161 2153 4176 2174
tri 4161 2138 4176 2153 nw
rect 4495 2153 4510 2174
tri 4133 2132 4139 2138 se
rect 4139 2132 4148 2138
rect 4133 2116 4148 2132
tri 4148 2125 4161 2138 nw
rect 4302 2130 4319 2144
rect 4351 2130 4368 2144
tri 4495 2138 4510 2153 ne
tri 4510 2138 4532 2160 sw
rect 4133 2080 4148 2088
rect 4214 2116 4274 2130
rect 4229 2106 4274 2116
rect 4229 2088 4257 2106
tri 4133 2065 4148 2080 ne
tri 4148 2065 4170 2087 sw
rect 4214 2078 4257 2088
rect 4272 2102 4274 2106
rect 4396 2116 4456 2130
tri 4510 2125 4523 2138 ne
rect 4523 2132 4532 2138
tri 4532 2132 4538 2138 sw
rect 4396 2106 4441 2116
rect 4272 2078 4346 2102
rect 4214 2074 4346 2078
tri 4346 2074 4374 2102 sw
rect 4396 2092 4398 2106
tri 4396 2090 4398 2092 ne
rect 4410 2088 4441 2106
rect 4410 2078 4456 2088
rect 4523 2117 4538 2132
tri 4148 2053 4160 2065 ne
rect 4160 2060 4170 2065
tri 4170 2060 4175 2065 sw
rect 4059 1714 4074 1942
rect 4160 1904 4175 2060
rect 4214 2018 4242 2074
tri 4334 2056 4352 2074 ne
rect 4352 2054 4374 2074
tri 4374 2054 4394 2074 sw
tri 4410 2060 4428 2078 ne
rect 4233 1984 4242 2018
rect 4276 2045 4318 2046
rect 4276 2011 4281 2045
rect 4311 2011 4318 2045
rect 4276 2002 4318 2011
rect 4352 2045 4394 2054
rect 4352 2011 4359 2045
rect 4389 2011 4394 2045
rect 4352 2006 4394 2011
rect 4428 2018 4456 2078
tri 4501 2065 4523 2087 se
rect 4523 2080 4538 2088
tri 4523 2065 4538 2080 nw
tri 4495 2059 4501 2065 se
rect 4501 2059 4510 2065
rect 4214 1974 4242 1984
tri 4242 1974 4266 1998 sw
rect 4214 1942 4256 1974
tri 4273 1966 4274 1967 sw
rect 4273 1942 4274 1966
tri 4276 1965 4313 2002 ne
rect 4313 1974 4318 2002
tri 4318 1974 4344 2000 sw
rect 4428 1984 4437 2018
rect 4428 1974 4456 1984
rect 4313 1965 4397 1974
tri 4313 1946 4332 1965 ne
rect 4332 1946 4397 1965
rect 4214 1920 4274 1942
rect 4396 1942 4397 1946
rect 4414 1942 4456 1974
rect 4396 1920 4456 1942
rect 4302 1904 4319 1918
rect 4351 1904 4368 1918
tri 4139 1868 4161 1890 se
rect 4161 1883 4176 1904
tri 4161 1868 4176 1883 nw
rect 4495 1883 4510 2059
tri 4510 2052 4523 2065 nw
rect 4596 1984 4611 2174
tri 4133 1862 4139 1868 se
rect 4139 1862 4148 1868
rect 4133 1846 4148 1862
tri 4148 1855 4161 1868 nw
rect 4302 1860 4319 1874
rect 4351 1860 4368 1874
tri 4495 1868 4510 1883 ne
tri 4510 1868 4532 1890 sw
rect 4133 1810 4148 1818
rect 4214 1846 4274 1860
rect 4229 1836 4274 1846
rect 4229 1818 4257 1836
tri 4133 1795 4148 1810 ne
tri 4148 1795 4170 1817 sw
rect 4214 1808 4257 1818
rect 4272 1832 4274 1836
rect 4396 1846 4456 1860
tri 4510 1855 4523 1868 ne
rect 4523 1862 4532 1868
tri 4532 1862 4538 1868 sw
rect 4396 1836 4441 1846
rect 4272 1808 4346 1832
rect 4214 1804 4346 1808
tri 4346 1804 4374 1832 sw
rect 4396 1822 4398 1836
tri 4396 1820 4398 1822 ne
rect 4410 1818 4441 1836
rect 4410 1808 4456 1818
rect 4523 1847 4538 1862
tri 4148 1783 4160 1795 ne
rect 4160 1790 4170 1795
tri 4170 1790 4175 1795 sw
rect 4059 1444 4074 1672
rect 4160 1634 4175 1790
rect 4214 1748 4242 1804
tri 4334 1786 4352 1804 ne
rect 4352 1784 4374 1804
tri 4374 1784 4394 1804 sw
tri 4410 1790 4428 1808 ne
rect 4233 1714 4242 1748
rect 4276 1775 4318 1776
rect 4276 1741 4281 1775
rect 4311 1741 4318 1775
rect 4276 1732 4318 1741
rect 4352 1775 4394 1784
rect 4352 1741 4359 1775
rect 4389 1741 4394 1775
rect 4352 1736 4394 1741
rect 4428 1748 4456 1808
tri 4501 1795 4523 1817 se
rect 4523 1810 4538 1818
tri 4523 1795 4538 1810 nw
tri 4495 1789 4501 1795 se
rect 4501 1789 4510 1795
rect 4214 1704 4242 1714
tri 4242 1704 4266 1728 sw
rect 4214 1672 4256 1704
tri 4273 1696 4274 1697 sw
rect 4273 1672 4274 1696
tri 4276 1695 4313 1732 ne
rect 4313 1704 4318 1732
tri 4318 1704 4344 1730 sw
rect 4428 1714 4437 1748
rect 4428 1704 4456 1714
rect 4313 1695 4397 1704
tri 4313 1676 4332 1695 ne
rect 4332 1676 4397 1695
rect 4214 1650 4274 1672
rect 4396 1672 4397 1676
rect 4414 1672 4456 1704
rect 4396 1650 4456 1672
rect 4302 1634 4319 1648
rect 4351 1634 4368 1648
tri 4139 1598 4161 1620 se
rect 4161 1613 4176 1634
tri 4161 1598 4176 1613 nw
rect 4495 1613 4510 1789
tri 4510 1782 4523 1795 nw
rect 4596 1714 4611 1942
tri 4133 1592 4139 1598 se
rect 4139 1592 4148 1598
rect 4133 1576 4148 1592
tri 4148 1585 4161 1598 nw
rect 4302 1590 4319 1604
rect 4351 1590 4368 1604
tri 4495 1598 4510 1613 ne
tri 4510 1598 4532 1620 sw
rect 4133 1540 4148 1548
rect 4214 1576 4274 1590
rect 4229 1566 4274 1576
rect 4229 1548 4257 1566
tri 4133 1525 4148 1540 ne
tri 4148 1525 4170 1547 sw
rect 4214 1538 4257 1548
rect 4272 1562 4274 1566
rect 4396 1576 4456 1590
tri 4510 1585 4523 1598 ne
rect 4523 1592 4532 1598
tri 4532 1592 4538 1598 sw
rect 4396 1566 4441 1576
rect 4272 1538 4346 1562
rect 4214 1534 4346 1538
tri 4346 1534 4374 1562 sw
rect 4396 1552 4398 1566
tri 4396 1550 4398 1552 ne
rect 4410 1548 4441 1566
rect 4410 1538 4456 1548
rect 4523 1577 4538 1592
tri 4148 1513 4160 1525 ne
rect 4160 1520 4170 1525
tri 4170 1520 4175 1525 sw
rect 4059 1174 4074 1402
rect 4160 1364 4175 1520
rect 4214 1478 4242 1534
tri 4334 1516 4352 1534 ne
rect 4352 1514 4374 1534
tri 4374 1514 4394 1534 sw
tri 4410 1520 4428 1538 ne
rect 4233 1444 4242 1478
rect 4276 1505 4318 1506
rect 4276 1471 4281 1505
rect 4311 1471 4318 1505
rect 4276 1462 4318 1471
rect 4352 1505 4394 1514
rect 4352 1471 4359 1505
rect 4389 1471 4394 1505
rect 4352 1466 4394 1471
rect 4428 1478 4456 1538
tri 4501 1525 4523 1547 se
rect 4523 1540 4538 1548
tri 4523 1525 4538 1540 nw
tri 4495 1519 4501 1525 se
rect 4501 1519 4510 1525
rect 4214 1434 4242 1444
tri 4242 1434 4266 1458 sw
rect 4214 1402 4256 1434
tri 4273 1426 4274 1427 sw
rect 4273 1402 4274 1426
tri 4276 1425 4313 1462 ne
rect 4313 1434 4318 1462
tri 4318 1434 4344 1460 sw
rect 4428 1444 4437 1478
rect 4428 1434 4456 1444
rect 4313 1425 4397 1434
tri 4313 1406 4332 1425 ne
rect 4332 1406 4397 1425
rect 4214 1380 4274 1402
rect 4396 1402 4397 1406
rect 4414 1402 4456 1434
rect 4396 1380 4456 1402
rect 4302 1364 4319 1378
rect 4351 1364 4368 1378
tri 4139 1328 4161 1350 se
rect 4161 1343 4176 1364
tri 4161 1328 4176 1343 nw
rect 4495 1343 4510 1519
tri 4510 1512 4523 1525 nw
rect 4596 1444 4611 1672
tri 4133 1322 4139 1328 se
rect 4139 1322 4148 1328
rect 4133 1306 4148 1322
tri 4148 1315 4161 1328 nw
rect 4302 1320 4319 1334
rect 4351 1320 4368 1334
tri 4495 1328 4510 1343 ne
tri 4510 1328 4532 1350 sw
rect 4133 1270 4148 1278
rect 4214 1306 4274 1320
rect 4229 1296 4274 1306
rect 4229 1278 4257 1296
tri 4133 1255 4148 1270 ne
tri 4148 1255 4170 1277 sw
rect 4214 1268 4257 1278
rect 4272 1292 4274 1296
rect 4396 1306 4456 1320
tri 4510 1315 4523 1328 ne
rect 4523 1322 4532 1328
tri 4532 1322 4538 1328 sw
rect 4396 1296 4441 1306
rect 4272 1268 4346 1292
rect 4214 1264 4346 1268
tri 4346 1264 4374 1292 sw
rect 4396 1282 4398 1296
tri 4396 1280 4398 1282 ne
rect 4410 1278 4441 1296
rect 4410 1268 4456 1278
rect 4523 1307 4538 1322
tri 4148 1243 4160 1255 ne
rect 4160 1250 4170 1255
tri 4170 1250 4175 1255 sw
rect 4059 904 4074 1132
rect 4160 1094 4175 1250
rect 4214 1208 4242 1264
tri 4334 1246 4352 1264 ne
rect 4352 1244 4374 1264
tri 4374 1244 4394 1264 sw
tri 4410 1250 4428 1268 ne
rect 4233 1174 4242 1208
rect 4276 1235 4318 1236
rect 4276 1201 4281 1235
rect 4311 1201 4318 1235
rect 4276 1192 4318 1201
rect 4352 1235 4394 1244
rect 4352 1201 4359 1235
rect 4389 1201 4394 1235
rect 4352 1196 4394 1201
rect 4428 1208 4456 1268
tri 4501 1255 4523 1277 se
rect 4523 1270 4538 1278
tri 4523 1255 4538 1270 nw
tri 4495 1249 4501 1255 se
rect 4501 1249 4510 1255
rect 4214 1164 4242 1174
tri 4242 1164 4266 1188 sw
rect 4214 1132 4256 1164
tri 4273 1156 4274 1157 sw
rect 4273 1132 4274 1156
tri 4276 1155 4313 1192 ne
rect 4313 1164 4318 1192
tri 4318 1164 4344 1190 sw
rect 4428 1174 4437 1208
rect 4428 1164 4456 1174
rect 4313 1155 4397 1164
tri 4313 1136 4332 1155 ne
rect 4332 1136 4397 1155
rect 4214 1110 4274 1132
rect 4396 1132 4397 1136
rect 4414 1132 4456 1164
rect 4396 1110 4456 1132
rect 4302 1094 4319 1108
rect 4351 1094 4368 1108
tri 4139 1058 4161 1080 se
rect 4161 1073 4176 1094
tri 4161 1058 4176 1073 nw
rect 4495 1073 4510 1249
tri 4510 1242 4523 1255 nw
rect 4596 1174 4611 1402
tri 4133 1052 4139 1058 se
rect 4139 1052 4148 1058
rect 4133 1036 4148 1052
tri 4148 1045 4161 1058 nw
rect 4302 1050 4319 1064
rect 4351 1050 4368 1064
tri 4495 1058 4510 1073 ne
tri 4510 1058 4532 1080 sw
rect 4133 1000 4148 1008
rect 4214 1036 4274 1050
rect 4229 1026 4274 1036
rect 4229 1008 4257 1026
tri 4133 985 4148 1000 ne
tri 4148 985 4170 1007 sw
rect 4214 998 4257 1008
rect 4272 1022 4274 1026
rect 4396 1036 4456 1050
tri 4510 1045 4523 1058 ne
rect 4523 1052 4532 1058
tri 4532 1052 4538 1058 sw
rect 4396 1026 4441 1036
rect 4272 998 4346 1022
rect 4214 994 4346 998
tri 4346 994 4374 1022 sw
rect 4396 1012 4398 1026
tri 4396 1010 4398 1012 ne
rect 4410 1008 4441 1026
rect 4410 998 4456 1008
rect 4523 1037 4538 1052
tri 4148 973 4160 985 ne
rect 4160 980 4170 985
tri 4170 980 4175 985 sw
rect 4059 634 4074 862
rect 4160 824 4175 980
rect 4214 938 4242 994
tri 4334 976 4352 994 ne
rect 4352 974 4374 994
tri 4374 974 4394 994 sw
tri 4410 980 4428 998 ne
rect 4233 904 4242 938
rect 4276 965 4318 966
rect 4276 931 4281 965
rect 4311 931 4318 965
rect 4276 922 4318 931
rect 4352 965 4394 974
rect 4352 931 4359 965
rect 4389 931 4394 965
rect 4352 926 4394 931
rect 4428 938 4456 998
tri 4501 985 4523 1007 se
rect 4523 1000 4538 1008
tri 4523 985 4538 1000 nw
tri 4495 979 4501 985 se
rect 4501 979 4510 985
rect 4214 894 4242 904
tri 4242 894 4266 918 sw
rect 4214 862 4256 894
tri 4273 886 4274 887 sw
rect 4273 862 4274 886
tri 4276 885 4313 922 ne
rect 4313 894 4318 922
tri 4318 894 4344 920 sw
rect 4428 904 4437 938
rect 4428 894 4456 904
rect 4313 885 4397 894
tri 4313 866 4332 885 ne
rect 4332 866 4397 885
rect 4214 840 4274 862
rect 4396 862 4397 866
rect 4414 862 4456 894
rect 4396 840 4456 862
rect 4302 824 4319 838
rect 4351 824 4368 838
tri 4139 788 4161 810 se
rect 4161 803 4176 824
tri 4161 788 4176 803 nw
rect 4495 803 4510 979
tri 4510 972 4523 985 nw
rect 4596 904 4611 1132
tri 4133 782 4139 788 se
rect 4139 782 4148 788
rect 4133 766 4148 782
tri 4148 775 4161 788 nw
rect 4302 780 4319 794
rect 4351 780 4368 794
tri 4495 788 4510 803 ne
tri 4510 788 4532 810 sw
rect 4133 730 4148 738
rect 4214 766 4274 780
rect 4229 756 4274 766
rect 4229 738 4257 756
tri 4133 715 4148 730 ne
tri 4148 715 4170 737 sw
rect 4214 728 4257 738
rect 4272 752 4274 756
rect 4396 766 4456 780
tri 4510 775 4523 788 ne
rect 4523 782 4532 788
tri 4532 782 4538 788 sw
rect 4396 756 4441 766
rect 4272 728 4346 752
rect 4214 724 4346 728
tri 4346 724 4374 752 sw
rect 4396 742 4398 756
tri 4396 740 4398 742 ne
rect 4410 738 4441 756
rect 4410 728 4456 738
rect 4523 767 4538 782
tri 4148 703 4160 715 ne
rect 4160 710 4170 715
tri 4170 710 4175 715 sw
rect 4059 364 4074 592
rect 4160 554 4175 710
rect 4214 668 4242 724
tri 4334 706 4352 724 ne
rect 4352 704 4374 724
tri 4374 704 4394 724 sw
tri 4410 710 4428 728 ne
rect 4233 634 4242 668
rect 4276 695 4318 696
rect 4276 661 4281 695
rect 4311 661 4318 695
rect 4276 652 4318 661
rect 4352 695 4394 704
rect 4352 661 4359 695
rect 4389 661 4394 695
rect 4352 656 4394 661
rect 4428 668 4456 728
tri 4501 715 4523 737 se
rect 4523 730 4538 738
tri 4523 715 4538 730 nw
tri 4495 709 4501 715 se
rect 4501 709 4510 715
rect 4214 624 4242 634
tri 4242 624 4266 648 sw
rect 4214 592 4256 624
tri 4273 616 4274 617 sw
rect 4273 592 4274 616
tri 4276 615 4313 652 ne
rect 4313 624 4318 652
tri 4318 624 4344 650 sw
rect 4428 634 4437 668
rect 4428 624 4456 634
rect 4313 615 4397 624
tri 4313 596 4332 615 ne
rect 4332 596 4397 615
rect 4214 570 4274 592
rect 4396 592 4397 596
rect 4414 592 4456 624
rect 4396 570 4456 592
rect 4302 554 4319 568
rect 4351 554 4368 568
tri 4139 518 4161 540 se
rect 4161 533 4176 554
tri 4161 518 4176 533 nw
rect 4495 533 4510 709
tri 4510 702 4523 715 nw
rect 4596 634 4611 862
tri 4133 512 4139 518 se
rect 4139 512 4148 518
rect 4133 496 4148 512
tri 4148 505 4161 518 nw
rect 4302 510 4319 524
rect 4351 510 4368 524
tri 4495 518 4510 533 ne
tri 4510 518 4532 540 sw
rect 4133 460 4148 468
rect 4214 496 4274 510
rect 4229 486 4274 496
rect 4229 468 4257 486
tri 4133 445 4148 460 ne
tri 4148 445 4170 467 sw
rect 4214 458 4257 468
rect 4272 482 4274 486
rect 4396 496 4456 510
tri 4510 505 4523 518 ne
rect 4523 512 4532 518
tri 4532 512 4538 518 sw
rect 4396 486 4441 496
rect 4272 458 4346 482
rect 4214 454 4346 458
tri 4346 454 4374 482 sw
rect 4396 472 4398 486
tri 4396 470 4398 472 ne
rect 4410 468 4441 486
rect 4410 458 4456 468
rect 4523 497 4538 512
tri 4148 433 4160 445 ne
rect 4160 440 4170 445
tri 4170 440 4175 445 sw
rect 4059 94 4074 322
rect 4160 284 4175 440
rect 4214 398 4242 454
tri 4334 436 4352 454 ne
rect 4352 434 4374 454
tri 4374 434 4394 454 sw
tri 4410 440 4428 458 ne
rect 4233 364 4242 398
rect 4276 425 4318 426
rect 4276 391 4281 425
rect 4311 391 4318 425
rect 4276 382 4318 391
rect 4352 425 4394 434
rect 4352 391 4359 425
rect 4389 391 4394 425
rect 4352 386 4394 391
rect 4428 398 4456 458
tri 4501 445 4523 467 se
rect 4523 460 4538 468
tri 4523 445 4538 460 nw
tri 4495 439 4501 445 se
rect 4501 439 4510 445
rect 4214 354 4242 364
tri 4242 354 4266 378 sw
rect 4214 322 4256 354
tri 4273 346 4274 347 sw
rect 4273 322 4274 346
tri 4276 345 4313 382 ne
rect 4313 354 4318 382
tri 4318 354 4344 380 sw
rect 4428 364 4437 398
rect 4428 354 4456 364
rect 4313 345 4397 354
tri 4313 326 4332 345 ne
rect 4332 326 4397 345
rect 4214 300 4274 322
rect 4396 322 4397 326
rect 4414 322 4456 354
rect 4396 300 4456 322
rect 4302 284 4319 298
rect 4351 284 4368 298
tri 4139 248 4161 270 se
rect 4161 263 4176 284
tri 4161 248 4176 263 nw
rect 4495 263 4510 439
tri 4510 432 4523 445 nw
rect 4596 364 4611 592
tri 4133 242 4139 248 se
rect 4139 242 4148 248
rect 4133 226 4148 242
tri 4148 235 4161 248 nw
rect 4302 240 4319 254
rect 4351 240 4368 254
tri 4495 248 4510 263 ne
tri 4510 248 4532 270 sw
rect 4133 190 4148 198
rect 4214 226 4274 240
rect 4229 216 4274 226
rect 4229 198 4257 216
tri 4133 175 4148 190 ne
tri 4148 175 4170 197 sw
rect 4214 188 4257 198
rect 4272 212 4274 216
rect 4396 226 4456 240
tri 4510 235 4523 248 ne
rect 4523 242 4532 248
tri 4532 242 4538 248 sw
rect 4396 216 4441 226
rect 4272 188 4346 212
rect 4214 184 4346 188
tri 4346 184 4374 212 sw
rect 4396 202 4398 216
tri 4396 200 4398 202 ne
rect 4410 198 4441 216
rect 4410 188 4456 198
rect 4523 227 4538 242
tri 4148 163 4160 175 ne
rect 4160 170 4170 175
tri 4170 170 4175 175 sw
rect 4059 -176 4074 52
rect 4160 14 4175 170
rect 4214 128 4242 184
tri 4334 166 4352 184 ne
rect 4352 164 4374 184
tri 4374 164 4394 184 sw
tri 4410 170 4428 188 ne
rect 4233 94 4242 128
rect 4276 155 4318 156
rect 4276 121 4281 155
rect 4311 121 4318 155
rect 4276 112 4318 121
rect 4352 155 4394 164
rect 4352 121 4359 155
rect 4389 121 4394 155
rect 4352 116 4394 121
rect 4428 128 4456 188
tri 4501 175 4523 197 se
rect 4523 190 4538 198
tri 4523 175 4538 190 nw
tri 4495 169 4501 175 se
rect 4501 169 4510 175
rect 4214 84 4242 94
tri 4242 84 4266 108 sw
rect 4214 52 4256 84
tri 4273 76 4274 77 sw
rect 4273 52 4274 76
tri 4276 75 4313 112 ne
rect 4313 84 4318 112
tri 4318 84 4344 110 sw
rect 4428 94 4437 128
rect 4428 84 4456 94
rect 4313 75 4397 84
tri 4313 56 4332 75 ne
rect 4332 56 4397 75
rect 4214 30 4274 52
rect 4396 52 4397 56
rect 4414 52 4456 84
rect 4396 30 4456 52
rect 4302 14 4319 28
rect 4351 14 4368 28
tri 4139 -22 4161 0 se
rect 4161 -7 4176 14
tri 4161 -22 4176 -7 nw
rect 4495 -7 4510 169
tri 4510 162 4523 175 nw
rect 4596 94 4611 322
tri 4133 -28 4139 -22 se
rect 4139 -28 4148 -22
rect 4133 -44 4148 -28
tri 4148 -35 4161 -22 nw
rect 4302 -30 4319 -16
rect 4351 -30 4368 -16
tri 4495 -22 4510 -7 ne
tri 4510 -22 4532 0 sw
rect 4133 -80 4148 -72
rect 4214 -44 4274 -30
rect 4229 -54 4274 -44
rect 4229 -72 4257 -54
tri 4133 -95 4148 -80 ne
tri 4148 -95 4170 -73 sw
rect 4214 -82 4257 -72
rect 4272 -58 4274 -54
rect 4396 -44 4456 -30
tri 4510 -35 4523 -22 ne
rect 4523 -28 4532 -22
tri 4532 -28 4538 -22 sw
rect 4396 -54 4441 -44
rect 4272 -82 4346 -58
rect 4214 -86 4346 -82
tri 4346 -86 4374 -58 sw
rect 4396 -68 4398 -54
tri 4396 -70 4398 -68 ne
rect 4410 -72 4441 -54
rect 4410 -82 4456 -72
rect 4523 -43 4538 -28
tri 4148 -107 4160 -95 ne
rect 4160 -100 4170 -95
tri 4170 -100 4175 -95 sw
rect 4059 -446 4074 -218
rect 4160 -256 4175 -100
rect 4214 -142 4242 -86
tri 4334 -104 4352 -86 ne
rect 4352 -106 4374 -86
tri 4374 -106 4394 -86 sw
tri 4410 -100 4428 -82 ne
rect 4233 -176 4242 -142
rect 4276 -115 4318 -114
rect 4276 -149 4281 -115
rect 4311 -149 4318 -115
rect 4276 -158 4318 -149
rect 4352 -115 4394 -106
rect 4352 -149 4359 -115
rect 4389 -149 4394 -115
rect 4352 -154 4394 -149
rect 4428 -142 4456 -82
tri 4501 -95 4523 -73 se
rect 4523 -80 4538 -72
tri 4523 -95 4538 -80 nw
tri 4495 -101 4501 -95 se
rect 4501 -101 4510 -95
rect 4214 -186 4242 -176
tri 4242 -186 4266 -162 sw
rect 4214 -218 4256 -186
tri 4273 -194 4274 -193 sw
rect 4273 -218 4274 -194
tri 4276 -195 4313 -158 ne
rect 4313 -186 4318 -158
tri 4318 -186 4344 -160 sw
rect 4428 -176 4437 -142
rect 4428 -186 4456 -176
rect 4313 -195 4397 -186
tri 4313 -214 4332 -195 ne
rect 4332 -214 4397 -195
rect 4214 -240 4274 -218
rect 4396 -218 4397 -214
rect 4414 -218 4456 -186
rect 4396 -240 4456 -218
rect 4302 -256 4319 -242
rect 4351 -256 4368 -242
tri 4139 -292 4161 -270 se
rect 4161 -277 4176 -256
tri 4161 -292 4176 -277 nw
rect 4495 -277 4510 -101
tri 4510 -108 4523 -95 nw
rect 4596 -176 4611 52
tri 4133 -298 4139 -292 se
rect 4139 -298 4148 -292
rect 4133 -314 4148 -298
tri 4148 -305 4161 -292 nw
rect 4302 -300 4319 -286
rect 4351 -300 4368 -286
tri 4495 -292 4510 -277 ne
tri 4510 -292 4532 -270 sw
rect 4133 -350 4148 -342
rect 4214 -314 4274 -300
rect 4229 -324 4274 -314
rect 4229 -342 4257 -324
tri 4133 -365 4148 -350 ne
tri 4148 -365 4170 -343 sw
rect 4214 -352 4257 -342
rect 4272 -328 4274 -324
rect 4396 -314 4456 -300
tri 4510 -305 4523 -292 ne
rect 4523 -298 4532 -292
tri 4532 -298 4538 -292 sw
rect 4396 -324 4441 -314
rect 4272 -352 4346 -328
rect 4214 -356 4346 -352
tri 4346 -356 4374 -328 sw
rect 4396 -338 4398 -324
tri 4396 -340 4398 -338 ne
rect 4410 -342 4441 -324
rect 4410 -352 4456 -342
rect 4523 -313 4538 -298
tri 4148 -377 4160 -365 ne
rect 4160 -370 4170 -365
tri 4170 -370 4175 -365 sw
rect 4059 -716 4074 -488
rect 4160 -526 4175 -370
rect 4214 -412 4242 -356
tri 4334 -374 4352 -356 ne
rect 4352 -376 4374 -356
tri 4374 -376 4394 -356 sw
tri 4410 -370 4428 -352 ne
rect 4233 -446 4242 -412
rect 4276 -385 4318 -384
rect 4276 -419 4281 -385
rect 4311 -419 4318 -385
rect 4276 -428 4318 -419
rect 4352 -385 4394 -376
rect 4352 -419 4359 -385
rect 4389 -419 4394 -385
rect 4352 -424 4394 -419
rect 4428 -412 4456 -352
tri 4501 -365 4523 -343 se
rect 4523 -350 4538 -342
tri 4523 -365 4538 -350 nw
tri 4495 -371 4501 -365 se
rect 4501 -371 4510 -365
rect 4214 -456 4242 -446
tri 4242 -456 4266 -432 sw
rect 4214 -488 4256 -456
tri 4273 -464 4274 -463 sw
rect 4273 -488 4274 -464
tri 4276 -465 4313 -428 ne
rect 4313 -456 4318 -428
tri 4318 -456 4344 -430 sw
rect 4428 -446 4437 -412
rect 4428 -456 4456 -446
rect 4313 -465 4397 -456
tri 4313 -484 4332 -465 ne
rect 4332 -484 4397 -465
rect 4214 -510 4274 -488
rect 4396 -488 4397 -484
rect 4414 -488 4456 -456
rect 4396 -510 4456 -488
rect 4302 -526 4319 -512
rect 4351 -526 4368 -512
tri 4139 -562 4161 -540 se
rect 4161 -547 4176 -526
tri 4161 -562 4176 -547 nw
rect 4495 -547 4510 -371
tri 4510 -378 4523 -365 nw
rect 4596 -446 4611 -218
tri 4133 -568 4139 -562 se
rect 4139 -568 4148 -562
rect 4133 -584 4148 -568
tri 4148 -575 4161 -562 nw
rect 4302 -570 4319 -556
rect 4351 -570 4368 -556
tri 4495 -562 4510 -547 ne
tri 4510 -562 4532 -540 sw
rect 4133 -620 4148 -612
rect 4214 -584 4274 -570
rect 4229 -594 4274 -584
rect 4229 -612 4257 -594
tri 4133 -635 4148 -620 ne
tri 4148 -635 4170 -613 sw
rect 4214 -622 4257 -612
rect 4272 -598 4274 -594
rect 4396 -584 4456 -570
tri 4510 -575 4523 -562 ne
rect 4523 -568 4532 -562
tri 4532 -568 4538 -562 sw
rect 4396 -594 4441 -584
rect 4272 -622 4346 -598
rect 4214 -626 4346 -622
tri 4346 -626 4374 -598 sw
rect 4396 -608 4398 -594
tri 4396 -610 4398 -608 ne
rect 4410 -612 4441 -594
rect 4410 -622 4456 -612
rect 4523 -583 4538 -568
tri 4148 -647 4160 -635 ne
rect 4160 -640 4170 -635
tri 4170 -640 4175 -635 sw
rect 4059 -986 4074 -758
rect 4160 -796 4175 -640
rect 4214 -682 4242 -626
tri 4334 -644 4352 -626 ne
rect 4352 -646 4374 -626
tri 4374 -646 4394 -626 sw
tri 4410 -640 4428 -622 ne
rect 4233 -716 4242 -682
rect 4276 -655 4318 -654
rect 4276 -689 4281 -655
rect 4311 -689 4318 -655
rect 4276 -698 4318 -689
rect 4352 -655 4394 -646
rect 4352 -689 4359 -655
rect 4389 -689 4394 -655
rect 4352 -694 4394 -689
rect 4428 -682 4456 -622
tri 4501 -635 4523 -613 se
rect 4523 -620 4538 -612
tri 4523 -635 4538 -620 nw
tri 4495 -641 4501 -635 se
rect 4501 -641 4510 -635
rect 4214 -726 4242 -716
tri 4242 -726 4266 -702 sw
rect 4214 -758 4256 -726
tri 4273 -734 4274 -733 sw
rect 4273 -758 4274 -734
tri 4276 -735 4313 -698 ne
rect 4313 -726 4318 -698
tri 4318 -726 4344 -700 sw
rect 4428 -716 4437 -682
rect 4428 -726 4456 -716
rect 4313 -735 4397 -726
tri 4313 -754 4332 -735 ne
rect 4332 -754 4397 -735
rect 4214 -780 4274 -758
rect 4396 -758 4397 -754
rect 4414 -758 4456 -726
rect 4396 -780 4456 -758
rect 4302 -796 4319 -782
rect 4351 -796 4368 -782
tri 4139 -832 4161 -810 se
rect 4161 -817 4176 -796
tri 4161 -832 4176 -817 nw
rect 4495 -817 4510 -641
tri 4510 -648 4523 -635 nw
rect 4596 -716 4611 -488
tri 4133 -838 4139 -832 se
rect 4139 -838 4148 -832
rect 4133 -854 4148 -838
tri 4148 -845 4161 -832 nw
rect 4302 -840 4319 -826
rect 4351 -840 4368 -826
tri 4495 -832 4510 -817 ne
tri 4510 -832 4532 -810 sw
rect 4133 -890 4148 -882
rect 4214 -854 4274 -840
rect 4229 -864 4274 -854
rect 4229 -882 4257 -864
tri 4133 -905 4148 -890 ne
tri 4148 -905 4170 -883 sw
rect 4214 -892 4257 -882
rect 4272 -868 4274 -864
rect 4396 -854 4456 -840
tri 4510 -845 4523 -832 ne
rect 4523 -838 4532 -832
tri 4532 -838 4538 -832 sw
rect 4396 -864 4441 -854
rect 4272 -892 4346 -868
rect 4214 -896 4346 -892
tri 4346 -896 4374 -868 sw
rect 4396 -878 4398 -864
tri 4396 -880 4398 -878 ne
rect 4410 -882 4441 -864
rect 4410 -892 4456 -882
rect 4523 -853 4538 -838
tri 4148 -917 4160 -905 ne
rect 4160 -910 4170 -905
tri 4170 -910 4175 -905 sw
rect 4059 -1256 4074 -1028
rect 4160 -1066 4175 -910
rect 4214 -952 4242 -896
tri 4334 -914 4352 -896 ne
rect 4352 -916 4374 -896
tri 4374 -916 4394 -896 sw
tri 4410 -910 4428 -892 ne
rect 4233 -986 4242 -952
rect 4276 -925 4318 -924
rect 4276 -959 4281 -925
rect 4311 -959 4318 -925
rect 4276 -968 4318 -959
rect 4352 -925 4394 -916
rect 4352 -959 4359 -925
rect 4389 -959 4394 -925
rect 4352 -964 4394 -959
rect 4428 -952 4456 -892
tri 4501 -905 4523 -883 se
rect 4523 -890 4538 -882
tri 4523 -905 4538 -890 nw
tri 4495 -911 4501 -905 se
rect 4501 -911 4510 -905
rect 4214 -996 4242 -986
tri 4242 -996 4266 -972 sw
rect 4214 -1028 4256 -996
tri 4273 -1004 4274 -1003 sw
rect 4273 -1028 4274 -1004
tri 4276 -1005 4313 -968 ne
rect 4313 -996 4318 -968
tri 4318 -996 4344 -970 sw
rect 4428 -986 4437 -952
rect 4428 -996 4456 -986
rect 4313 -1005 4397 -996
tri 4313 -1024 4332 -1005 ne
rect 4332 -1024 4397 -1005
rect 4214 -1050 4274 -1028
rect 4396 -1028 4397 -1024
rect 4414 -1028 4456 -996
rect 4396 -1050 4456 -1028
rect 4302 -1066 4319 -1052
rect 4351 -1066 4368 -1052
tri 4139 -1102 4161 -1080 se
rect 4161 -1087 4176 -1066
tri 4161 -1102 4176 -1087 nw
rect 4495 -1087 4510 -911
tri 4510 -918 4523 -905 nw
rect 4596 -986 4611 -758
tri 4133 -1108 4139 -1102 se
rect 4139 -1108 4148 -1102
rect 4133 -1124 4148 -1108
tri 4148 -1115 4161 -1102 nw
rect 4302 -1110 4319 -1096
rect 4351 -1110 4368 -1096
tri 4495 -1102 4510 -1087 ne
tri 4510 -1102 4532 -1080 sw
rect 4133 -1160 4148 -1152
rect 4214 -1124 4274 -1110
rect 4229 -1134 4274 -1124
rect 4229 -1152 4257 -1134
tri 4133 -1175 4148 -1160 ne
tri 4148 -1175 4170 -1153 sw
rect 4214 -1162 4257 -1152
rect 4272 -1138 4274 -1134
rect 4396 -1124 4456 -1110
tri 4510 -1115 4523 -1102 ne
rect 4523 -1108 4532 -1102
tri 4532 -1108 4538 -1102 sw
rect 4396 -1134 4441 -1124
rect 4272 -1162 4346 -1138
rect 4214 -1166 4346 -1162
tri 4346 -1166 4374 -1138 sw
rect 4396 -1148 4398 -1134
tri 4396 -1150 4398 -1148 ne
rect 4410 -1152 4441 -1134
rect 4410 -1162 4456 -1152
rect 4523 -1123 4538 -1108
tri 4148 -1187 4160 -1175 ne
rect 4160 -1180 4170 -1175
tri 4170 -1180 4175 -1175 sw
rect 4059 -1526 4074 -1298
rect 4160 -1336 4175 -1180
rect 4214 -1222 4242 -1166
tri 4334 -1184 4352 -1166 ne
rect 4352 -1186 4374 -1166
tri 4374 -1186 4394 -1166 sw
tri 4410 -1180 4428 -1162 ne
rect 4233 -1256 4242 -1222
rect 4276 -1195 4318 -1194
rect 4276 -1229 4281 -1195
rect 4311 -1229 4318 -1195
rect 4276 -1238 4318 -1229
rect 4352 -1195 4394 -1186
rect 4352 -1229 4359 -1195
rect 4389 -1229 4394 -1195
rect 4352 -1234 4394 -1229
rect 4428 -1222 4456 -1162
tri 4501 -1175 4523 -1153 se
rect 4523 -1160 4538 -1152
tri 4523 -1175 4538 -1160 nw
tri 4495 -1181 4501 -1175 se
rect 4501 -1181 4510 -1175
rect 4214 -1266 4242 -1256
tri 4242 -1266 4266 -1242 sw
rect 4214 -1298 4256 -1266
tri 4273 -1274 4274 -1273 sw
rect 4273 -1298 4274 -1274
tri 4276 -1275 4313 -1238 ne
rect 4313 -1266 4318 -1238
tri 4318 -1266 4344 -1240 sw
rect 4428 -1256 4437 -1222
rect 4428 -1266 4456 -1256
rect 4313 -1275 4397 -1266
tri 4313 -1294 4332 -1275 ne
rect 4332 -1294 4397 -1275
rect 4214 -1320 4274 -1298
rect 4396 -1298 4397 -1294
rect 4414 -1298 4456 -1266
rect 4396 -1320 4456 -1298
rect 4302 -1336 4319 -1322
rect 4351 -1336 4368 -1322
tri 4139 -1372 4161 -1350 se
rect 4161 -1357 4176 -1336
tri 4161 -1372 4176 -1357 nw
rect 4495 -1357 4510 -1181
tri 4510 -1188 4523 -1175 nw
rect 4596 -1256 4611 -1028
tri 4133 -1378 4139 -1372 se
rect 4139 -1378 4148 -1372
rect 4133 -1394 4148 -1378
tri 4148 -1385 4161 -1372 nw
rect 4302 -1380 4319 -1366
rect 4351 -1380 4368 -1366
tri 4495 -1372 4510 -1357 ne
tri 4510 -1372 4532 -1350 sw
rect 4133 -1430 4148 -1422
rect 4214 -1394 4274 -1380
rect 4229 -1404 4274 -1394
rect 4229 -1422 4257 -1404
tri 4133 -1445 4148 -1430 ne
tri 4148 -1445 4170 -1423 sw
rect 4214 -1432 4257 -1422
rect 4272 -1408 4274 -1404
rect 4396 -1394 4456 -1380
tri 4510 -1385 4523 -1372 ne
rect 4523 -1378 4532 -1372
tri 4532 -1378 4538 -1372 sw
rect 4396 -1404 4441 -1394
rect 4272 -1432 4346 -1408
rect 4214 -1436 4346 -1432
tri 4346 -1436 4374 -1408 sw
rect 4396 -1418 4398 -1404
tri 4396 -1420 4398 -1418 ne
rect 4410 -1422 4441 -1404
rect 4410 -1432 4456 -1422
rect 4523 -1393 4538 -1378
tri 4148 -1457 4160 -1445 ne
rect 4160 -1450 4170 -1445
tri 4170 -1450 4175 -1445 sw
rect 4059 -1796 4074 -1568
rect 4160 -1606 4175 -1450
rect 4214 -1492 4242 -1436
tri 4334 -1454 4352 -1436 ne
rect 4352 -1456 4374 -1436
tri 4374 -1456 4394 -1436 sw
tri 4410 -1450 4428 -1432 ne
rect 4233 -1526 4242 -1492
rect 4276 -1465 4318 -1464
rect 4276 -1499 4281 -1465
rect 4311 -1499 4318 -1465
rect 4276 -1508 4318 -1499
rect 4352 -1465 4394 -1456
rect 4352 -1499 4359 -1465
rect 4389 -1499 4394 -1465
rect 4352 -1504 4394 -1499
rect 4428 -1492 4456 -1432
tri 4501 -1445 4523 -1423 se
rect 4523 -1430 4538 -1422
tri 4523 -1445 4538 -1430 nw
tri 4495 -1451 4501 -1445 se
rect 4501 -1451 4510 -1445
rect 4214 -1536 4242 -1526
tri 4242 -1536 4266 -1512 sw
rect 4214 -1568 4256 -1536
tri 4273 -1544 4274 -1543 sw
rect 4273 -1568 4274 -1544
tri 4276 -1545 4313 -1508 ne
rect 4313 -1536 4318 -1508
tri 4318 -1536 4344 -1510 sw
rect 4428 -1526 4437 -1492
rect 4428 -1536 4456 -1526
rect 4313 -1545 4397 -1536
tri 4313 -1564 4332 -1545 ne
rect 4332 -1564 4397 -1545
rect 4214 -1590 4274 -1568
rect 4396 -1568 4397 -1564
rect 4414 -1568 4456 -1536
rect 4396 -1590 4456 -1568
rect 4302 -1606 4319 -1592
rect 4351 -1606 4368 -1592
tri 4139 -1642 4161 -1620 se
rect 4161 -1627 4176 -1606
tri 4161 -1642 4176 -1627 nw
rect 4495 -1627 4510 -1451
tri 4510 -1458 4523 -1445 nw
rect 4596 -1526 4611 -1298
tri 4133 -1648 4139 -1642 se
rect 4139 -1648 4148 -1642
rect 4133 -1664 4148 -1648
tri 4148 -1655 4161 -1642 nw
rect 4302 -1650 4319 -1636
rect 4351 -1650 4368 -1636
tri 4495 -1642 4510 -1627 ne
tri 4510 -1642 4532 -1620 sw
rect 4133 -1700 4148 -1692
rect 4214 -1664 4274 -1650
rect 4229 -1674 4274 -1664
rect 4229 -1692 4257 -1674
tri 4133 -1715 4148 -1700 ne
tri 4148 -1715 4170 -1693 sw
rect 4214 -1702 4257 -1692
rect 4272 -1678 4274 -1674
rect 4396 -1664 4456 -1650
tri 4510 -1655 4523 -1642 ne
rect 4523 -1648 4532 -1642
tri 4532 -1648 4538 -1642 sw
rect 4396 -1674 4441 -1664
rect 4272 -1702 4346 -1678
rect 4214 -1706 4346 -1702
tri 4346 -1706 4374 -1678 sw
rect 4396 -1688 4398 -1674
tri 4396 -1690 4398 -1688 ne
rect 4410 -1692 4441 -1674
rect 4410 -1702 4456 -1692
rect 4523 -1663 4538 -1648
tri 4148 -1727 4160 -1715 ne
rect 4160 -1720 4170 -1715
tri 4170 -1720 4175 -1715 sw
rect 4059 -2066 4074 -1838
rect 4160 -1876 4175 -1720
rect 4214 -1762 4242 -1706
tri 4334 -1724 4352 -1706 ne
rect 4352 -1726 4374 -1706
tri 4374 -1726 4394 -1706 sw
tri 4410 -1720 4428 -1702 ne
rect 4233 -1796 4242 -1762
rect 4276 -1735 4318 -1734
rect 4276 -1769 4281 -1735
rect 4311 -1769 4318 -1735
rect 4276 -1778 4318 -1769
rect 4352 -1735 4394 -1726
rect 4352 -1769 4359 -1735
rect 4389 -1769 4394 -1735
rect 4352 -1774 4394 -1769
rect 4428 -1762 4456 -1702
tri 4501 -1715 4523 -1693 se
rect 4523 -1700 4538 -1692
tri 4523 -1715 4538 -1700 nw
tri 4495 -1721 4501 -1715 se
rect 4501 -1721 4510 -1715
rect 4214 -1806 4242 -1796
tri 4242 -1806 4266 -1782 sw
rect 4214 -1838 4256 -1806
tri 4273 -1814 4274 -1813 sw
rect 4273 -1838 4274 -1814
tri 4276 -1815 4313 -1778 ne
rect 4313 -1806 4318 -1778
tri 4318 -1806 4344 -1780 sw
rect 4428 -1796 4437 -1762
rect 4428 -1806 4456 -1796
rect 4313 -1815 4397 -1806
tri 4313 -1834 4332 -1815 ne
rect 4332 -1834 4397 -1815
rect 4214 -1860 4274 -1838
rect 4396 -1838 4397 -1834
rect 4414 -1838 4456 -1806
rect 4396 -1860 4456 -1838
rect 4302 -1876 4319 -1862
rect 4351 -1876 4368 -1862
tri 4139 -1912 4161 -1890 se
rect 4161 -1897 4176 -1876
tri 4161 -1912 4176 -1897 nw
rect 4495 -1897 4510 -1721
tri 4510 -1728 4523 -1715 nw
rect 4596 -1796 4611 -1568
tri 4133 -1918 4139 -1912 se
rect 4139 -1918 4148 -1912
rect 4133 -1934 4148 -1918
tri 4148 -1925 4161 -1912 nw
rect 4302 -1920 4319 -1906
rect 4351 -1920 4368 -1906
tri 4495 -1912 4510 -1897 ne
tri 4510 -1912 4532 -1890 sw
rect 4133 -1970 4148 -1962
rect 4214 -1934 4274 -1920
rect 4229 -1944 4274 -1934
rect 4229 -1962 4257 -1944
tri 4133 -1985 4148 -1970 ne
tri 4148 -1985 4170 -1963 sw
rect 4214 -1972 4257 -1962
rect 4272 -1948 4274 -1944
rect 4396 -1934 4456 -1920
tri 4510 -1925 4523 -1912 ne
rect 4523 -1918 4532 -1912
tri 4532 -1918 4538 -1912 sw
rect 4396 -1944 4441 -1934
rect 4272 -1972 4346 -1948
rect 4214 -1976 4346 -1972
tri 4346 -1976 4374 -1948 sw
rect 4396 -1958 4398 -1944
tri 4396 -1960 4398 -1958 ne
rect 4410 -1962 4441 -1944
rect 4410 -1972 4456 -1962
rect 4523 -1933 4538 -1918
tri 4148 -1997 4160 -1985 ne
rect 4160 -1990 4170 -1985
tri 4170 -1990 4175 -1985 sw
rect 4059 -2146 4074 -2108
rect 4160 -2146 4175 -1990
rect 4214 -2032 4242 -1976
tri 4334 -1994 4352 -1976 ne
rect 4352 -1996 4374 -1976
tri 4374 -1996 4394 -1976 sw
tri 4410 -1990 4428 -1972 ne
rect 4233 -2066 4242 -2032
rect 4276 -2005 4318 -2004
rect 4276 -2039 4281 -2005
rect 4311 -2039 4318 -2005
rect 4276 -2048 4318 -2039
rect 4352 -2005 4394 -1996
rect 4352 -2039 4359 -2005
rect 4389 -2039 4394 -2005
rect 4352 -2044 4394 -2039
rect 4428 -2032 4456 -1972
tri 4501 -1985 4523 -1963 se
rect 4523 -1970 4538 -1962
tri 4523 -1985 4538 -1970 nw
tri 4495 -1991 4501 -1985 se
rect 4501 -1991 4510 -1985
rect 4214 -2076 4242 -2066
tri 4242 -2076 4266 -2052 sw
rect 4214 -2108 4256 -2076
tri 4273 -2084 4274 -2083 sw
rect 4273 -2108 4274 -2084
tri 4276 -2085 4313 -2048 ne
rect 4313 -2076 4318 -2048
tri 4318 -2076 4344 -2050 sw
rect 4428 -2066 4437 -2032
rect 4428 -2076 4456 -2066
rect 4313 -2085 4397 -2076
tri 4313 -2104 4332 -2085 ne
rect 4332 -2104 4397 -2085
rect 4214 -2130 4274 -2108
rect 4396 -2108 4397 -2104
rect 4414 -2108 4456 -2076
rect 4396 -2130 4456 -2108
rect 4302 -2146 4319 -2132
rect 4351 -2146 4368 -2132
rect 4495 -2146 4510 -1991
tri 4510 -1998 4523 -1985 nw
rect 4596 -2066 4611 -1838
rect 4596 -2146 4611 -2108
rect 4639 1984 4654 2174
tri 4719 2138 4741 2160 se
rect 4741 2153 4756 2174
tri 4741 2138 4756 2153 nw
rect 5075 2153 5090 2174
tri 4713 2132 4719 2138 se
rect 4719 2132 4728 2138
rect 4713 2116 4728 2132
tri 4728 2125 4741 2138 nw
rect 4882 2130 4899 2144
rect 4931 2130 4948 2144
tri 5075 2138 5090 2153 ne
tri 5090 2138 5112 2160 sw
rect 4713 2080 4728 2088
rect 4794 2116 4854 2130
rect 4809 2106 4854 2116
rect 4809 2088 4837 2106
tri 4713 2065 4728 2080 ne
tri 4728 2065 4750 2087 sw
rect 4794 2078 4837 2088
rect 4852 2102 4854 2106
rect 4976 2116 5036 2130
tri 5090 2125 5103 2138 ne
rect 5103 2132 5112 2138
tri 5112 2132 5118 2138 sw
rect 4976 2106 5021 2116
rect 4852 2078 4926 2102
rect 4794 2074 4926 2078
tri 4926 2074 4954 2102 sw
rect 4976 2092 4978 2106
tri 4976 2090 4978 2092 ne
rect 4990 2088 5021 2106
rect 4990 2078 5036 2088
rect 5103 2117 5118 2132
tri 4728 2053 4740 2065 ne
rect 4740 2060 4750 2065
tri 4750 2060 4755 2065 sw
rect 4639 1714 4654 1942
rect 4740 1904 4755 2060
rect 4794 2018 4822 2074
tri 4914 2056 4932 2074 ne
rect 4932 2054 4954 2074
tri 4954 2054 4974 2074 sw
tri 4990 2060 5008 2078 ne
rect 4813 1984 4822 2018
rect 4856 2045 4898 2046
rect 4856 2011 4861 2045
rect 4891 2011 4898 2045
rect 4856 2002 4898 2011
rect 4932 2045 4974 2054
rect 4932 2011 4939 2045
rect 4969 2011 4974 2045
rect 4932 2006 4974 2011
rect 5008 2018 5036 2078
tri 5081 2065 5103 2087 se
rect 5103 2080 5118 2088
tri 5103 2065 5118 2080 nw
tri 5075 2059 5081 2065 se
rect 5081 2059 5090 2065
rect 4794 1974 4822 1984
tri 4822 1974 4846 1998 sw
rect 4794 1942 4836 1974
tri 4853 1966 4854 1967 sw
rect 4853 1942 4854 1966
tri 4856 1965 4893 2002 ne
rect 4893 1974 4898 2002
tri 4898 1974 4924 2000 sw
rect 5008 1984 5017 2018
rect 5008 1974 5036 1984
rect 4893 1965 4977 1974
tri 4893 1946 4912 1965 ne
rect 4912 1946 4977 1965
rect 4794 1920 4854 1942
rect 4976 1942 4977 1946
rect 4994 1942 5036 1974
rect 4976 1920 5036 1942
rect 4882 1904 4899 1918
rect 4931 1904 4948 1918
tri 4719 1868 4741 1890 se
rect 4741 1883 4756 1904
tri 4741 1868 4756 1883 nw
rect 5075 1883 5090 2059
tri 5090 2052 5103 2065 nw
rect 5176 1984 5191 2174
tri 4713 1862 4719 1868 se
rect 4719 1862 4728 1868
rect 4713 1846 4728 1862
tri 4728 1855 4741 1868 nw
rect 4882 1860 4899 1874
rect 4931 1860 4948 1874
tri 5075 1868 5090 1883 ne
tri 5090 1868 5112 1890 sw
rect 4713 1810 4728 1818
rect 4794 1846 4854 1860
rect 4809 1836 4854 1846
rect 4809 1818 4837 1836
tri 4713 1795 4728 1810 ne
tri 4728 1795 4750 1817 sw
rect 4794 1808 4837 1818
rect 4852 1832 4854 1836
rect 4976 1846 5036 1860
tri 5090 1855 5103 1868 ne
rect 5103 1862 5112 1868
tri 5112 1862 5118 1868 sw
rect 4976 1836 5021 1846
rect 4852 1808 4926 1832
rect 4794 1804 4926 1808
tri 4926 1804 4954 1832 sw
rect 4976 1822 4978 1836
tri 4976 1820 4978 1822 ne
rect 4990 1818 5021 1836
rect 4990 1808 5036 1818
rect 5103 1847 5118 1862
tri 4728 1783 4740 1795 ne
rect 4740 1790 4750 1795
tri 4750 1790 4755 1795 sw
rect 4639 1444 4654 1672
rect 4740 1682 4755 1790
rect 4794 1748 4822 1804
tri 4914 1786 4932 1804 ne
rect 4932 1784 4954 1804
tri 4954 1784 4974 1804 sw
tri 4990 1790 5008 1808 ne
rect 4813 1714 4822 1748
rect 4856 1775 4898 1776
rect 4856 1741 4861 1775
rect 4891 1741 4898 1775
rect 4856 1732 4898 1741
rect 4932 1775 4974 1784
rect 4932 1741 4939 1775
rect 4969 1741 4974 1775
rect 4932 1736 4974 1741
rect 5008 1748 5036 1808
tri 5081 1795 5103 1817 se
rect 5103 1810 5118 1818
tri 5103 1795 5118 1810 nw
tri 5075 1789 5081 1795 se
rect 5081 1789 5090 1795
rect 4794 1704 4822 1714
tri 4822 1704 4846 1728 sw
rect 4740 1634 4756 1682
rect 4794 1672 4836 1704
tri 4853 1696 4854 1697 sw
rect 4853 1672 4854 1696
tri 4856 1695 4893 1732 ne
rect 4893 1704 4898 1732
tri 4898 1704 4924 1730 sw
rect 5008 1714 5017 1748
rect 5008 1704 5036 1714
rect 4893 1695 4977 1704
tri 4893 1676 4912 1695 ne
rect 4912 1676 4977 1695
rect 4794 1650 4854 1672
rect 4976 1672 4977 1676
rect 4994 1672 5036 1704
rect 4976 1650 5036 1672
rect 4882 1634 4899 1648
rect 4931 1634 4948 1648
tri 4719 1598 4741 1620 se
rect 4741 1613 4756 1634
tri 4741 1598 4756 1613 nw
rect 5075 1613 5090 1789
tri 5090 1782 5103 1795 nw
rect 5176 1714 5191 1942
tri 4713 1592 4719 1598 se
rect 4719 1592 4728 1598
rect 4713 1576 4728 1592
tri 4728 1585 4741 1598 nw
rect 4882 1590 4899 1604
rect 4931 1590 4948 1604
tri 5075 1598 5090 1613 ne
tri 5090 1598 5112 1620 sw
rect 4713 1540 4728 1548
rect 4794 1576 4854 1590
rect 4809 1566 4854 1576
rect 4809 1548 4837 1566
tri 4713 1525 4728 1540 ne
tri 4728 1525 4750 1547 sw
rect 4794 1538 4837 1548
rect 4852 1562 4854 1566
rect 4976 1576 5036 1590
tri 5090 1585 5103 1598 ne
rect 5103 1592 5112 1598
tri 5112 1592 5118 1598 sw
rect 4976 1566 5021 1576
rect 4852 1538 4926 1562
rect 4794 1534 4926 1538
tri 4926 1534 4954 1562 sw
rect 4976 1552 4978 1566
tri 4976 1550 4978 1552 ne
rect 4990 1548 5021 1566
rect 4990 1538 5036 1548
rect 5103 1577 5118 1592
tri 4728 1513 4740 1525 ne
rect 4740 1520 4750 1525
tri 4750 1520 4755 1525 sw
rect 4639 1174 4654 1402
rect 4740 1364 4755 1520
rect 4794 1478 4822 1534
tri 4914 1516 4932 1534 ne
rect 4932 1514 4954 1534
tri 4954 1514 4974 1534 sw
tri 4990 1520 5008 1538 ne
rect 4813 1444 4822 1478
rect 4856 1505 4898 1506
rect 4856 1471 4861 1505
rect 4891 1471 4898 1505
rect 4856 1462 4898 1471
rect 4932 1505 4974 1514
rect 4932 1471 4939 1505
rect 4969 1471 4974 1505
rect 4932 1466 4974 1471
rect 5008 1478 5036 1538
tri 5081 1525 5103 1547 se
rect 5103 1540 5118 1548
tri 5103 1525 5118 1540 nw
tri 5075 1519 5081 1525 se
rect 5081 1519 5090 1525
rect 4794 1434 4822 1444
tri 4822 1434 4846 1458 sw
rect 4794 1402 4836 1434
tri 4853 1426 4854 1427 sw
rect 4853 1402 4854 1426
tri 4856 1425 4893 1462 ne
rect 4893 1434 4898 1462
tri 4898 1434 4924 1460 sw
rect 5008 1444 5017 1478
rect 5008 1434 5036 1444
rect 4893 1425 4977 1434
tri 4893 1406 4912 1425 ne
rect 4912 1406 4977 1425
rect 4794 1380 4854 1402
rect 4976 1402 4977 1406
rect 4994 1402 5036 1434
rect 4976 1380 5036 1402
rect 4882 1364 4899 1378
rect 4931 1364 4948 1378
tri 4719 1328 4741 1350 se
rect 4741 1343 4756 1364
tri 4741 1328 4756 1343 nw
rect 5075 1343 5090 1519
tri 5090 1512 5103 1525 nw
rect 5176 1444 5191 1672
tri 4713 1322 4719 1328 se
rect 4719 1322 4728 1328
rect 4713 1306 4728 1322
tri 4728 1315 4741 1328 nw
rect 4882 1320 4899 1334
rect 4931 1320 4948 1334
tri 5075 1328 5090 1343 ne
tri 5090 1328 5112 1350 sw
rect 4713 1270 4728 1278
rect 4794 1306 4854 1320
rect 4809 1296 4854 1306
rect 4809 1278 4837 1296
tri 4713 1255 4728 1270 ne
tri 4728 1255 4750 1277 sw
rect 4794 1268 4837 1278
rect 4852 1292 4854 1296
rect 4976 1306 5036 1320
tri 5090 1315 5103 1328 ne
rect 5103 1322 5112 1328
tri 5112 1322 5118 1328 sw
rect 4976 1296 5021 1306
rect 4852 1268 4926 1292
rect 4794 1264 4926 1268
tri 4926 1264 4954 1292 sw
rect 4976 1282 4978 1296
tri 4976 1280 4978 1282 ne
rect 4990 1278 5021 1296
rect 4990 1268 5036 1278
rect 5103 1307 5118 1322
tri 4728 1243 4740 1255 ne
rect 4740 1250 4750 1255
tri 4750 1250 4755 1255 sw
rect 4639 903 4654 1132
rect 4740 1141 4755 1250
rect 4794 1208 4822 1264
tri 4914 1246 4932 1264 ne
rect 4932 1244 4954 1264
tri 4954 1244 4974 1264 sw
tri 4990 1250 5008 1268 ne
rect 4813 1174 4822 1208
rect 4856 1235 4898 1236
rect 4856 1201 4861 1235
rect 4891 1201 4898 1235
rect 4856 1192 4898 1201
rect 4932 1235 4974 1244
rect 4932 1201 4939 1235
rect 4969 1201 4974 1235
rect 4932 1196 4974 1201
rect 5008 1208 5036 1268
tri 5081 1255 5103 1277 se
rect 5103 1270 5118 1278
tri 5103 1255 5118 1270 nw
tri 5075 1249 5081 1255 se
rect 5081 1249 5090 1255
rect 4794 1164 4822 1174
tri 4822 1164 4846 1188 sw
rect 4740 1094 4756 1141
rect 4794 1132 4836 1164
tri 4853 1156 4854 1157 sw
rect 4853 1132 4854 1156
tri 4856 1155 4893 1192 ne
rect 4893 1164 4898 1192
tri 4898 1164 4924 1190 sw
rect 5008 1174 5017 1208
rect 5008 1164 5036 1174
rect 4893 1155 4977 1164
tri 4893 1136 4912 1155 ne
rect 4912 1136 4977 1155
rect 4794 1110 4854 1132
rect 4976 1132 4977 1136
rect 4994 1132 5036 1164
rect 4976 1110 5036 1132
rect 4882 1094 4899 1108
rect 4931 1094 4948 1108
tri 4719 1057 4741 1079 se
rect 4741 1072 4756 1094
tri 4741 1057 4756 1072 nw
rect 5075 1072 5090 1249
tri 5090 1242 5103 1255 nw
rect 5176 1174 5191 1402
tri 4713 1051 4719 1057 se
rect 4719 1051 4728 1057
rect 4713 1035 4728 1051
tri 4728 1044 4741 1057 nw
rect 4882 1049 4899 1063
rect 4931 1049 4948 1063
tri 5075 1057 5090 1072 ne
tri 5090 1057 5112 1079 sw
rect 4713 999 4728 1007
rect 4794 1035 4854 1049
rect 4809 1025 4854 1035
rect 4809 1007 4837 1025
tri 4713 984 4728 999 ne
tri 4728 984 4750 1006 sw
rect 4794 997 4837 1007
rect 4852 1021 4854 1025
rect 4976 1035 5036 1049
tri 5090 1044 5103 1057 ne
rect 5103 1051 5112 1057
tri 5112 1051 5118 1057 sw
rect 4976 1025 5021 1035
rect 4852 997 4926 1021
rect 4794 993 4926 997
tri 4926 993 4954 1021 sw
rect 4976 1011 4978 1025
tri 4976 1009 4978 1011 ne
rect 4990 1007 5021 1025
rect 4990 997 5036 1007
rect 5103 1036 5118 1051
tri 4728 972 4740 984 ne
rect 4740 979 4750 984
tri 4750 979 4755 984 sw
rect 4639 633 4654 861
rect 4740 823 4755 979
rect 4794 937 4822 993
tri 4914 975 4932 993 ne
rect 4932 973 4954 993
tri 4954 973 4974 993 sw
tri 4990 979 5008 997 ne
rect 4813 903 4822 937
rect 4856 964 4898 965
rect 4856 930 4861 964
rect 4891 930 4898 964
rect 4856 921 4898 930
rect 4932 964 4974 973
rect 4932 930 4939 964
rect 4969 930 4974 964
rect 4932 925 4974 930
rect 5008 937 5036 997
tri 5081 984 5103 1006 se
rect 5103 999 5118 1007
tri 5103 984 5118 999 nw
tri 5075 978 5081 984 se
rect 5081 978 5090 984
rect 4794 893 4822 903
tri 4822 893 4846 917 sw
rect 4794 861 4836 893
tri 4853 885 4854 886 sw
rect 4853 861 4854 885
tri 4856 884 4893 921 ne
rect 4893 893 4898 921
tri 4898 893 4924 919 sw
rect 5008 903 5017 937
rect 5008 893 5036 903
rect 4893 884 4977 893
tri 4893 865 4912 884 ne
rect 4912 865 4977 884
rect 4794 839 4854 861
rect 4976 861 4977 865
rect 4994 861 5036 893
rect 4976 839 5036 861
rect 4882 823 4899 837
rect 4931 823 4948 837
tri 4719 787 4741 809 se
rect 4741 802 4756 823
tri 4741 787 4756 802 nw
rect 5075 802 5090 978
tri 5090 971 5103 984 nw
rect 5176 903 5191 1132
tri 4713 781 4719 787 se
rect 4719 781 4728 787
rect 4713 765 4728 781
tri 4728 774 4741 787 nw
rect 4882 779 4899 793
rect 4931 779 4948 793
tri 5075 787 5090 802 ne
tri 5090 787 5112 809 sw
rect 4713 729 4728 737
rect 4794 765 4854 779
rect 4809 755 4854 765
rect 4809 737 4837 755
tri 4713 714 4728 729 ne
tri 4728 714 4750 736 sw
rect 4794 727 4837 737
rect 4852 751 4854 755
rect 4976 765 5036 779
tri 5090 774 5103 787 ne
rect 5103 781 5112 787
tri 5112 781 5118 787 sw
rect 4976 755 5021 765
rect 4852 727 4926 751
rect 4794 723 4926 727
tri 4926 723 4954 751 sw
rect 4976 741 4978 755
tri 4976 739 4978 741 ne
rect 4990 737 5021 755
rect 4990 727 5036 737
rect 5103 766 5118 781
tri 4728 702 4740 714 ne
rect 4740 709 4750 714
tri 4750 709 4755 714 sw
rect 4639 363 4654 591
rect 4740 601 4755 709
rect 4794 667 4822 723
tri 4914 705 4932 723 ne
rect 4932 703 4954 723
tri 4954 703 4974 723 sw
tri 4990 709 5008 727 ne
rect 4813 633 4822 667
rect 4856 694 4898 695
rect 4856 660 4861 694
rect 4891 660 4898 694
rect 4856 651 4898 660
rect 4932 694 4974 703
rect 4932 660 4939 694
rect 4969 660 4974 694
rect 4932 655 4974 660
rect 5008 667 5036 727
tri 5081 714 5103 736 se
rect 5103 729 5118 737
tri 5103 714 5118 729 nw
tri 5075 708 5081 714 se
rect 5081 708 5090 714
rect 4794 623 4822 633
tri 4822 623 4846 647 sw
rect 4740 553 4756 601
rect 4794 591 4836 623
tri 4853 615 4854 616 sw
rect 4853 591 4854 615
tri 4856 614 4893 651 ne
rect 4893 623 4898 651
tri 4898 623 4924 649 sw
rect 5008 633 5017 667
rect 5008 623 5036 633
rect 4893 614 4977 623
tri 4893 595 4912 614 ne
rect 4912 595 4977 614
rect 4794 569 4854 591
rect 4976 591 4977 595
rect 4994 591 5036 623
rect 4976 569 5036 591
rect 4882 553 4899 567
rect 4931 553 4948 567
tri 4719 517 4741 539 se
rect 4741 532 4756 553
tri 4741 517 4756 532 nw
rect 5075 532 5090 708
tri 5090 701 5103 714 nw
rect 5176 633 5191 861
tri 4713 511 4719 517 se
rect 4719 511 4728 517
rect 4713 495 4728 511
tri 4728 504 4741 517 nw
rect 4882 509 4899 523
rect 4931 509 4948 523
tri 5075 517 5090 532 ne
tri 5090 517 5112 539 sw
rect 4713 459 4728 467
rect 4794 495 4854 509
rect 4809 485 4854 495
rect 4809 467 4837 485
tri 4713 444 4728 459 ne
tri 4728 444 4750 466 sw
rect 4794 457 4837 467
rect 4852 481 4854 485
rect 4976 495 5036 509
tri 5090 504 5103 517 ne
rect 5103 511 5112 517
tri 5112 511 5118 517 sw
rect 4976 485 5021 495
rect 4852 457 4926 481
rect 4794 453 4926 457
tri 4926 453 4954 481 sw
rect 4976 471 4978 485
tri 4976 469 4978 471 ne
rect 4990 467 5021 485
rect 4990 457 5036 467
rect 5103 496 5118 511
tri 4728 432 4740 444 ne
rect 4740 439 4750 444
tri 4750 439 4755 444 sw
rect 4639 93 4654 321
rect 4740 283 4755 439
rect 4794 397 4822 453
tri 4914 435 4932 453 ne
rect 4932 433 4954 453
tri 4954 433 4974 453 sw
tri 4990 439 5008 457 ne
rect 4813 363 4822 397
rect 4856 424 4898 425
rect 4856 390 4861 424
rect 4891 390 4898 424
rect 4856 381 4898 390
rect 4932 424 4974 433
rect 4932 390 4939 424
rect 4969 390 4974 424
rect 4932 385 4974 390
rect 5008 397 5036 457
tri 5081 444 5103 466 se
rect 5103 459 5118 467
tri 5103 444 5118 459 nw
tri 5075 438 5081 444 se
rect 5081 438 5090 444
rect 4794 353 4822 363
tri 4822 353 4846 377 sw
rect 4794 321 4836 353
tri 4853 345 4854 346 sw
rect 4853 321 4854 345
tri 4856 344 4893 381 ne
rect 4893 353 4898 381
tri 4898 353 4924 379 sw
rect 5008 363 5017 397
rect 5008 353 5036 363
rect 4893 344 4977 353
tri 4893 325 4912 344 ne
rect 4912 325 4977 344
rect 4794 299 4854 321
rect 4976 321 4977 325
rect 4994 321 5036 353
rect 4976 299 5036 321
rect 4882 283 4899 297
rect 4931 283 4948 297
tri 4719 247 4741 269 se
rect 4741 262 4756 283
tri 4741 247 4756 262 nw
rect 5075 262 5090 438
tri 5090 431 5103 444 nw
rect 5176 363 5191 591
tri 4713 241 4719 247 se
rect 4719 241 4728 247
rect 4713 225 4728 241
tri 4728 234 4741 247 nw
rect 4882 239 4899 253
rect 4931 239 4948 253
tri 5075 247 5090 262 ne
tri 5090 247 5112 269 sw
rect 4713 189 4728 197
rect 4794 225 4854 239
rect 4809 215 4854 225
rect 4809 197 4837 215
tri 4713 174 4728 189 ne
tri 4728 174 4750 196 sw
rect 4794 187 4837 197
rect 4852 211 4854 215
rect 4976 225 5036 239
tri 5090 234 5103 247 ne
rect 5103 241 5112 247
tri 5112 241 5118 247 sw
rect 4976 215 5021 225
rect 4852 187 4926 211
rect 4794 183 4926 187
tri 4926 183 4954 211 sw
rect 4976 201 4978 215
tri 4976 199 4978 201 ne
rect 4990 197 5021 215
rect 4990 187 5036 197
rect 5103 226 5118 241
tri 4728 162 4740 174 ne
rect 4740 169 4750 174
tri 4750 169 4755 174 sw
rect 4639 -177 4654 51
rect 4740 61 4755 169
rect 4794 127 4822 183
tri 4914 165 4932 183 ne
rect 4932 163 4954 183
tri 4954 163 4974 183 sw
tri 4990 169 5008 187 ne
rect 4813 93 4822 127
rect 4856 154 4898 155
rect 4856 120 4861 154
rect 4891 120 4898 154
rect 4856 111 4898 120
rect 4932 154 4974 163
rect 4932 120 4939 154
rect 4969 120 4974 154
rect 4932 115 4974 120
rect 5008 127 5036 187
tri 5081 174 5103 196 se
rect 5103 189 5118 197
tri 5103 174 5118 189 nw
tri 5075 168 5081 174 se
rect 5081 168 5090 174
rect 4794 83 4822 93
tri 4822 83 4846 107 sw
rect 4740 13 4756 61
rect 4794 51 4836 83
tri 4853 75 4854 76 sw
rect 4853 51 4854 75
tri 4856 74 4893 111 ne
rect 4893 83 4898 111
tri 4898 83 4924 109 sw
rect 5008 93 5017 127
rect 5008 83 5036 93
rect 4893 74 4977 83
tri 4893 55 4912 74 ne
rect 4912 55 4977 74
rect 4794 29 4854 51
rect 4976 51 4977 55
rect 4994 51 5036 83
rect 4976 29 5036 51
rect 4882 13 4899 27
rect 4931 13 4948 27
tri 4719 -23 4741 -1 se
rect 4741 -8 4756 13
tri 4741 -23 4756 -8 nw
rect 5075 -8 5090 168
tri 5090 161 5103 174 nw
rect 5176 93 5191 321
tri 4713 -29 4719 -23 se
rect 4719 -29 4728 -23
rect 4713 -45 4728 -29
tri 4728 -36 4741 -23 nw
rect 4882 -31 4899 -17
rect 4931 -31 4948 -17
tri 5075 -23 5090 -8 ne
tri 5090 -23 5112 -1 sw
rect 4713 -81 4728 -73
rect 4794 -45 4854 -31
rect 4809 -55 4854 -45
rect 4809 -73 4837 -55
tri 4713 -96 4728 -81 ne
tri 4728 -96 4750 -74 sw
rect 4794 -83 4837 -73
rect 4852 -59 4854 -55
rect 4976 -45 5036 -31
tri 5090 -36 5103 -23 ne
rect 5103 -29 5112 -23
tri 5112 -29 5118 -23 sw
rect 4976 -55 5021 -45
rect 4852 -83 4926 -59
rect 4794 -87 4926 -83
tri 4926 -87 4954 -59 sw
rect 4976 -69 4978 -55
tri 4976 -71 4978 -69 ne
rect 4990 -73 5021 -55
rect 4990 -83 5036 -73
rect 5103 -44 5118 -29
tri 4728 -108 4740 -96 ne
rect 4740 -101 4750 -96
tri 4750 -101 4755 -96 sw
rect 4639 -447 4654 -219
rect 4740 -257 4755 -101
rect 4794 -143 4822 -87
tri 4914 -105 4932 -87 ne
rect 4932 -107 4954 -87
tri 4954 -107 4974 -87 sw
tri 4990 -101 5008 -83 ne
rect 4813 -177 4822 -143
rect 4856 -116 4898 -115
rect 4856 -150 4861 -116
rect 4891 -150 4898 -116
rect 4856 -159 4898 -150
rect 4932 -116 4974 -107
rect 4932 -150 4939 -116
rect 4969 -150 4974 -116
rect 4932 -155 4974 -150
rect 5008 -143 5036 -83
tri 5081 -96 5103 -74 se
rect 5103 -81 5118 -73
tri 5103 -96 5118 -81 nw
tri 5075 -102 5081 -96 se
rect 5081 -102 5090 -96
rect 4794 -187 4822 -177
tri 4822 -187 4846 -163 sw
rect 4794 -219 4836 -187
tri 4853 -195 4854 -194 sw
rect 4853 -219 4854 -195
tri 4856 -196 4893 -159 ne
rect 4893 -187 4898 -159
tri 4898 -187 4924 -161 sw
rect 5008 -177 5017 -143
rect 5008 -187 5036 -177
rect 4893 -196 4977 -187
tri 4893 -215 4912 -196 ne
rect 4912 -215 4977 -196
rect 4794 -241 4854 -219
rect 4976 -219 4977 -215
rect 4994 -219 5036 -187
rect 4976 -241 5036 -219
rect 4882 -257 4899 -243
rect 4931 -257 4948 -243
tri 4719 -293 4741 -271 se
rect 4741 -278 4756 -257
tri 4741 -293 4756 -278 nw
rect 5075 -278 5090 -102
tri 5090 -109 5103 -96 nw
rect 5176 -177 5191 51
tri 4713 -299 4719 -293 se
rect 4719 -299 4728 -293
rect 4713 -315 4728 -299
tri 4728 -306 4741 -293 nw
rect 4882 -301 4899 -287
rect 4931 -301 4948 -287
tri 5075 -293 5090 -278 ne
tri 5090 -293 5112 -271 sw
rect 4713 -351 4728 -343
rect 4794 -315 4854 -301
rect 4809 -325 4854 -315
rect 4809 -343 4837 -325
tri 4713 -366 4728 -351 ne
tri 4728 -366 4750 -344 sw
rect 4794 -353 4837 -343
rect 4852 -329 4854 -325
rect 4976 -315 5036 -301
tri 5090 -306 5103 -293 ne
rect 5103 -299 5112 -293
tri 5112 -299 5118 -293 sw
rect 4976 -325 5021 -315
rect 4852 -353 4926 -329
rect 4794 -357 4926 -353
tri 4926 -357 4954 -329 sw
rect 4976 -339 4978 -325
tri 4976 -341 4978 -339 ne
rect 4990 -343 5021 -325
rect 4990 -353 5036 -343
rect 5103 -314 5118 -299
tri 4728 -378 4740 -366 ne
rect 4740 -371 4750 -366
tri 4750 -371 4755 -366 sw
rect 4639 -717 4654 -489
rect 4740 -479 4755 -371
rect 4794 -413 4822 -357
tri 4914 -375 4932 -357 ne
rect 4932 -377 4954 -357
tri 4954 -377 4974 -357 sw
tri 4990 -371 5008 -353 ne
rect 4813 -447 4822 -413
rect 4856 -386 4898 -385
rect 4856 -420 4861 -386
rect 4891 -420 4898 -386
rect 4856 -429 4898 -420
rect 4932 -386 4974 -377
rect 4932 -420 4939 -386
rect 4969 -420 4974 -386
rect 4932 -425 4974 -420
rect 5008 -413 5036 -353
tri 5081 -366 5103 -344 se
rect 5103 -351 5118 -343
tri 5103 -366 5118 -351 nw
tri 5075 -372 5081 -366 se
rect 5081 -372 5090 -366
rect 4794 -457 4822 -447
tri 4822 -457 4846 -433 sw
rect 4740 -527 4756 -479
rect 4794 -489 4836 -457
tri 4853 -465 4854 -464 sw
rect 4853 -489 4854 -465
tri 4856 -466 4893 -429 ne
rect 4893 -457 4898 -429
tri 4898 -457 4924 -431 sw
rect 5008 -447 5017 -413
rect 5008 -457 5036 -447
rect 4893 -466 4977 -457
tri 4893 -485 4912 -466 ne
rect 4912 -485 4977 -466
rect 4794 -511 4854 -489
rect 4976 -489 4977 -485
rect 4994 -489 5036 -457
rect 4976 -511 5036 -489
rect 4882 -527 4899 -513
rect 4931 -527 4948 -513
tri 4719 -563 4741 -541 se
rect 4741 -548 4756 -527
tri 4741 -563 4756 -548 nw
rect 5075 -548 5090 -372
tri 5090 -379 5103 -366 nw
rect 5176 -447 5191 -219
tri 4713 -569 4719 -563 se
rect 4719 -569 4728 -563
rect 4713 -585 4728 -569
tri 4728 -576 4741 -563 nw
rect 4882 -571 4899 -557
rect 4931 -571 4948 -557
tri 5075 -563 5090 -548 ne
tri 5090 -563 5112 -541 sw
rect 4713 -621 4728 -613
rect 4794 -585 4854 -571
rect 4809 -595 4854 -585
rect 4809 -613 4837 -595
tri 4713 -636 4728 -621 ne
tri 4728 -636 4750 -614 sw
rect 4794 -623 4837 -613
rect 4852 -599 4854 -595
rect 4976 -585 5036 -571
tri 5090 -576 5103 -563 ne
rect 5103 -569 5112 -563
tri 5112 -569 5118 -563 sw
rect 4976 -595 5021 -585
rect 4852 -623 4926 -599
rect 4794 -627 4926 -623
tri 4926 -627 4954 -599 sw
rect 4976 -609 4978 -595
tri 4976 -611 4978 -609 ne
rect 4990 -613 5021 -595
rect 4990 -623 5036 -613
rect 5103 -584 5118 -569
tri 4728 -648 4740 -636 ne
rect 4740 -641 4750 -636
tri 4750 -641 4755 -636 sw
rect 4639 -987 4654 -759
rect 4740 -797 4755 -641
rect 4794 -683 4822 -627
tri 4914 -645 4932 -627 ne
rect 4932 -647 4954 -627
tri 4954 -647 4974 -627 sw
tri 4990 -641 5008 -623 ne
rect 4813 -717 4822 -683
rect 4856 -656 4898 -655
rect 4856 -690 4861 -656
rect 4891 -690 4898 -656
rect 4856 -699 4898 -690
rect 4932 -656 4974 -647
rect 4932 -690 4939 -656
rect 4969 -690 4974 -656
rect 4932 -695 4974 -690
rect 5008 -683 5036 -623
tri 5081 -636 5103 -614 se
rect 5103 -621 5118 -613
tri 5103 -636 5118 -621 nw
tri 5075 -642 5081 -636 se
rect 5081 -642 5090 -636
rect 4794 -727 4822 -717
tri 4822 -727 4846 -703 sw
rect 4794 -759 4836 -727
tri 4853 -735 4854 -734 sw
rect 4853 -759 4854 -735
tri 4856 -736 4893 -699 ne
rect 4893 -727 4898 -699
tri 4898 -727 4924 -701 sw
rect 5008 -717 5017 -683
rect 5008 -727 5036 -717
rect 4893 -736 4977 -727
tri 4893 -755 4912 -736 ne
rect 4912 -755 4977 -736
rect 4794 -781 4854 -759
rect 4976 -759 4977 -755
rect 4994 -759 5036 -727
rect 4976 -781 5036 -759
rect 4882 -797 4899 -783
rect 4931 -797 4948 -783
tri 4719 -833 4741 -811 se
rect 4741 -818 4756 -797
tri 4741 -833 4756 -818 nw
rect 5075 -818 5090 -642
tri 5090 -649 5103 -636 nw
rect 5176 -717 5191 -489
tri 4713 -839 4719 -833 se
rect 4719 -839 4728 -833
rect 4713 -855 4728 -839
tri 4728 -846 4741 -833 nw
rect 4882 -841 4899 -827
rect 4931 -841 4948 -827
tri 5075 -833 5090 -818 ne
tri 5090 -833 5112 -811 sw
rect 4713 -891 4728 -883
rect 4794 -855 4854 -841
rect 4809 -865 4854 -855
rect 4809 -883 4837 -865
tri 4713 -906 4728 -891 ne
tri 4728 -906 4750 -884 sw
rect 4794 -893 4837 -883
rect 4852 -869 4854 -865
rect 4976 -855 5036 -841
tri 5090 -846 5103 -833 ne
rect 5103 -839 5112 -833
tri 5112 -839 5118 -833 sw
rect 4976 -865 5021 -855
rect 4852 -893 4926 -869
rect 4794 -897 4926 -893
tri 4926 -897 4954 -869 sw
rect 4976 -879 4978 -865
tri 4976 -881 4978 -879 ne
rect 4990 -883 5021 -865
rect 4990 -893 5036 -883
rect 5103 -854 5118 -839
tri 4728 -918 4740 -906 ne
rect 4740 -911 4750 -906
tri 4750 -911 4755 -906 sw
rect 4639 -1257 4654 -1029
rect 4740 -1019 4755 -911
rect 4794 -953 4822 -897
tri 4914 -915 4932 -897 ne
rect 4932 -917 4954 -897
tri 4954 -917 4974 -897 sw
tri 4990 -911 5008 -893 ne
rect 4813 -987 4822 -953
rect 4856 -926 4898 -925
rect 4856 -960 4861 -926
rect 4891 -960 4898 -926
rect 4856 -969 4898 -960
rect 4932 -926 4974 -917
rect 4932 -960 4939 -926
rect 4969 -960 4974 -926
rect 4932 -965 4974 -960
rect 5008 -953 5036 -893
tri 5081 -906 5103 -884 se
rect 5103 -891 5118 -883
tri 5103 -906 5118 -891 nw
tri 5075 -912 5081 -906 se
rect 5081 -912 5090 -906
rect 4794 -997 4822 -987
tri 4822 -997 4846 -973 sw
rect 4740 -1067 4756 -1019
rect 4794 -1029 4836 -997
tri 4853 -1005 4854 -1004 sw
rect 4853 -1029 4854 -1005
tri 4856 -1006 4893 -969 ne
rect 4893 -997 4898 -969
tri 4898 -997 4924 -971 sw
rect 5008 -987 5017 -953
rect 5008 -997 5036 -987
rect 4893 -1006 4977 -997
tri 4893 -1025 4912 -1006 ne
rect 4912 -1025 4977 -1006
rect 4794 -1051 4854 -1029
rect 4976 -1029 4977 -1025
rect 4994 -1029 5036 -997
rect 4976 -1051 5036 -1029
rect 4882 -1067 4899 -1053
rect 4931 -1067 4948 -1053
tri 4719 -1103 4741 -1081 se
rect 4741 -1088 4756 -1067
tri 4741 -1103 4756 -1088 nw
rect 5075 -1088 5090 -912
tri 5090 -919 5103 -906 nw
rect 5176 -987 5191 -759
tri 4713 -1109 4719 -1103 se
rect 4719 -1109 4728 -1103
rect 4713 -1125 4728 -1109
tri 4728 -1116 4741 -1103 nw
rect 4882 -1111 4899 -1097
rect 4931 -1111 4948 -1097
tri 5075 -1103 5090 -1088 ne
tri 5090 -1103 5112 -1081 sw
rect 4713 -1161 4728 -1153
rect 4794 -1125 4854 -1111
rect 4809 -1135 4854 -1125
rect 4809 -1153 4837 -1135
tri 4713 -1176 4728 -1161 ne
tri 4728 -1176 4750 -1154 sw
rect 4794 -1163 4837 -1153
rect 4852 -1139 4854 -1135
rect 4976 -1125 5036 -1111
tri 5090 -1116 5103 -1103 ne
rect 5103 -1109 5112 -1103
tri 5112 -1109 5118 -1103 sw
rect 4976 -1135 5021 -1125
rect 4852 -1163 4926 -1139
rect 4794 -1167 4926 -1163
tri 4926 -1167 4954 -1139 sw
rect 4976 -1149 4978 -1135
tri 4976 -1151 4978 -1149 ne
rect 4990 -1153 5021 -1135
rect 4990 -1163 5036 -1153
rect 5103 -1124 5118 -1109
tri 4728 -1188 4740 -1176 ne
rect 4740 -1181 4750 -1176
tri 4750 -1181 4755 -1176 sw
rect 4639 -1527 4654 -1299
rect 4740 -1337 4755 -1181
rect 4794 -1223 4822 -1167
tri 4914 -1185 4932 -1167 ne
rect 4932 -1187 4954 -1167
tri 4954 -1187 4974 -1167 sw
tri 4990 -1181 5008 -1163 ne
rect 4813 -1257 4822 -1223
rect 4856 -1196 4898 -1195
rect 4856 -1230 4861 -1196
rect 4891 -1230 4898 -1196
rect 4856 -1239 4898 -1230
rect 4932 -1196 4974 -1187
rect 4932 -1230 4939 -1196
rect 4969 -1230 4974 -1196
rect 4932 -1235 4974 -1230
rect 5008 -1223 5036 -1163
tri 5081 -1176 5103 -1154 se
rect 5103 -1161 5118 -1153
tri 5103 -1176 5118 -1161 nw
tri 5075 -1182 5081 -1176 se
rect 5081 -1182 5090 -1176
rect 4794 -1267 4822 -1257
tri 4822 -1267 4846 -1243 sw
rect 4794 -1299 4836 -1267
tri 4853 -1275 4854 -1274 sw
rect 4853 -1299 4854 -1275
tri 4856 -1276 4893 -1239 ne
rect 4893 -1267 4898 -1239
tri 4898 -1267 4924 -1241 sw
rect 5008 -1257 5017 -1223
rect 5008 -1267 5036 -1257
rect 4893 -1276 4977 -1267
tri 4893 -1295 4912 -1276 ne
rect 4912 -1295 4977 -1276
rect 4794 -1321 4854 -1299
rect 4976 -1299 4977 -1295
rect 4994 -1299 5036 -1267
rect 4976 -1321 5036 -1299
rect 4882 -1337 4899 -1323
rect 4931 -1337 4948 -1323
tri 4719 -1373 4741 -1351 se
rect 4741 -1358 4756 -1337
tri 4741 -1373 4756 -1358 nw
rect 5075 -1358 5090 -1182
tri 5090 -1189 5103 -1176 nw
rect 5176 -1257 5191 -1029
tri 4713 -1379 4719 -1373 se
rect 4719 -1379 4728 -1373
rect 4713 -1395 4728 -1379
tri 4728 -1386 4741 -1373 nw
rect 4882 -1381 4899 -1367
rect 4931 -1381 4948 -1367
tri 5075 -1373 5090 -1358 ne
tri 5090 -1373 5112 -1351 sw
rect 4713 -1431 4728 -1423
rect 4794 -1395 4854 -1381
rect 4809 -1405 4854 -1395
rect 4809 -1423 4837 -1405
tri 4713 -1446 4728 -1431 ne
tri 4728 -1446 4750 -1424 sw
rect 4794 -1433 4837 -1423
rect 4852 -1409 4854 -1405
rect 4976 -1395 5036 -1381
tri 5090 -1386 5103 -1373 ne
rect 5103 -1379 5112 -1373
tri 5112 -1379 5118 -1373 sw
rect 4976 -1405 5021 -1395
rect 4852 -1433 4926 -1409
rect 4794 -1437 4926 -1433
tri 4926 -1437 4954 -1409 sw
rect 4976 -1419 4978 -1405
tri 4976 -1421 4978 -1419 ne
rect 4990 -1423 5021 -1405
rect 4990 -1433 5036 -1423
rect 5103 -1394 5118 -1379
tri 4728 -1458 4740 -1446 ne
rect 4740 -1451 4750 -1446
tri 4750 -1451 4755 -1446 sw
rect 4639 -1797 4654 -1569
rect 4740 -1559 4755 -1451
rect 4794 -1493 4822 -1437
tri 4914 -1455 4932 -1437 ne
rect 4932 -1457 4954 -1437
tri 4954 -1457 4974 -1437 sw
tri 4990 -1451 5008 -1433 ne
rect 4813 -1527 4822 -1493
rect 4856 -1466 4898 -1465
rect 4856 -1500 4861 -1466
rect 4891 -1500 4898 -1466
rect 4856 -1509 4898 -1500
rect 4932 -1466 4974 -1457
rect 4932 -1500 4939 -1466
rect 4969 -1500 4974 -1466
rect 4932 -1505 4974 -1500
rect 5008 -1493 5036 -1433
tri 5081 -1446 5103 -1424 se
rect 5103 -1431 5118 -1423
tri 5103 -1446 5118 -1431 nw
tri 5075 -1452 5081 -1446 se
rect 5081 -1452 5090 -1446
rect 4794 -1537 4822 -1527
tri 4822 -1537 4846 -1513 sw
rect 4740 -1607 4756 -1559
rect 4794 -1569 4836 -1537
tri 4853 -1545 4854 -1544 sw
rect 4853 -1569 4854 -1545
tri 4856 -1546 4893 -1509 ne
rect 4893 -1537 4898 -1509
tri 4898 -1537 4924 -1511 sw
rect 5008 -1527 5017 -1493
rect 5008 -1537 5036 -1527
rect 4893 -1546 4977 -1537
tri 4893 -1565 4912 -1546 ne
rect 4912 -1565 4977 -1546
rect 4794 -1591 4854 -1569
rect 4976 -1569 4977 -1565
rect 4994 -1569 5036 -1537
rect 4976 -1591 5036 -1569
rect 4882 -1607 4899 -1593
rect 4931 -1607 4948 -1593
tri 4719 -1643 4741 -1621 se
rect 4741 -1628 4756 -1607
tri 4741 -1643 4756 -1628 nw
rect 5075 -1628 5090 -1452
tri 5090 -1459 5103 -1446 nw
rect 5176 -1527 5191 -1299
tri 4713 -1649 4719 -1643 se
rect 4719 -1649 4728 -1643
rect 4713 -1665 4728 -1649
tri 4728 -1656 4741 -1643 nw
rect 4882 -1651 4899 -1637
rect 4931 -1651 4948 -1637
tri 5075 -1643 5090 -1628 ne
tri 5090 -1643 5112 -1621 sw
rect 4713 -1701 4728 -1693
rect 4794 -1665 4854 -1651
rect 4809 -1675 4854 -1665
rect 4809 -1693 4837 -1675
tri 4713 -1716 4728 -1701 ne
tri 4728 -1716 4750 -1694 sw
rect 4794 -1703 4837 -1693
rect 4852 -1679 4854 -1675
rect 4976 -1665 5036 -1651
tri 5090 -1656 5103 -1643 ne
rect 5103 -1649 5112 -1643
tri 5112 -1649 5118 -1643 sw
rect 4976 -1675 5021 -1665
rect 4852 -1703 4926 -1679
rect 4794 -1707 4926 -1703
tri 4926 -1707 4954 -1679 sw
rect 4976 -1689 4978 -1675
tri 4976 -1691 4978 -1689 ne
rect 4990 -1693 5021 -1675
rect 4990 -1703 5036 -1693
rect 5103 -1664 5118 -1649
tri 4728 -1728 4740 -1716 ne
rect 4740 -1721 4750 -1716
tri 4750 -1721 4755 -1716 sw
rect 4639 -2067 4654 -1839
rect 4740 -1877 4755 -1721
rect 4794 -1763 4822 -1707
tri 4914 -1725 4932 -1707 ne
rect 4932 -1727 4954 -1707
tri 4954 -1727 4974 -1707 sw
tri 4990 -1721 5008 -1703 ne
rect 4813 -1797 4822 -1763
rect 4856 -1736 4898 -1735
rect 4856 -1770 4861 -1736
rect 4891 -1770 4898 -1736
rect 4856 -1779 4898 -1770
rect 4932 -1736 4974 -1727
rect 4932 -1770 4939 -1736
rect 4969 -1770 4974 -1736
rect 4932 -1775 4974 -1770
rect 5008 -1763 5036 -1703
tri 5081 -1716 5103 -1694 se
rect 5103 -1701 5118 -1693
tri 5103 -1716 5118 -1701 nw
tri 5075 -1722 5081 -1716 se
rect 5081 -1722 5090 -1716
rect 4794 -1807 4822 -1797
tri 4822 -1807 4846 -1783 sw
rect 4794 -1839 4836 -1807
tri 4853 -1815 4854 -1814 sw
rect 4853 -1839 4854 -1815
tri 4856 -1816 4893 -1779 ne
rect 4893 -1807 4898 -1779
tri 4898 -1807 4924 -1781 sw
rect 5008 -1797 5017 -1763
rect 5008 -1807 5036 -1797
rect 4893 -1816 4977 -1807
tri 4893 -1835 4912 -1816 ne
rect 4912 -1835 4977 -1816
rect 4794 -1861 4854 -1839
rect 4976 -1839 4977 -1835
rect 4994 -1839 5036 -1807
rect 4976 -1861 5036 -1839
rect 4882 -1877 4899 -1863
rect 4931 -1877 4948 -1863
tri 4719 -1913 4741 -1891 se
rect 4741 -1898 4756 -1877
tri 4741 -1913 4756 -1898 nw
rect 5075 -1898 5090 -1722
tri 5090 -1729 5103 -1716 nw
rect 5176 -1797 5191 -1569
tri 4713 -1919 4719 -1913 se
rect 4719 -1919 4728 -1913
rect 4713 -1935 4728 -1919
tri 4728 -1926 4741 -1913 nw
rect 4882 -1921 4899 -1907
rect 4931 -1921 4948 -1907
tri 5075 -1913 5090 -1898 ne
tri 5090 -1913 5112 -1891 sw
rect 4713 -1971 4728 -1963
rect 4794 -1935 4854 -1921
rect 4809 -1945 4854 -1935
rect 4809 -1963 4837 -1945
tri 4713 -1986 4728 -1971 ne
tri 4728 -1986 4750 -1964 sw
rect 4794 -1973 4837 -1963
rect 4852 -1949 4854 -1945
rect 4976 -1935 5036 -1921
tri 5090 -1926 5103 -1913 ne
rect 5103 -1919 5112 -1913
tri 5112 -1919 5118 -1913 sw
rect 4976 -1945 5021 -1935
rect 4852 -1973 4926 -1949
rect 4794 -1977 4926 -1973
tri 4926 -1977 4954 -1949 sw
rect 4976 -1959 4978 -1945
tri 4976 -1961 4978 -1959 ne
rect 4990 -1963 5021 -1945
rect 4990 -1973 5036 -1963
rect 5103 -1934 5118 -1919
tri 4728 -1998 4740 -1986 ne
rect 4740 -1991 4750 -1986
tri 4750 -1991 4755 -1986 sw
rect 4639 -2147 4654 -2109
rect 4740 -2147 4755 -1991
rect 4794 -2033 4822 -1977
tri 4914 -1995 4932 -1977 ne
rect 4932 -1997 4954 -1977
tri 4954 -1997 4974 -1977 sw
tri 4990 -1991 5008 -1973 ne
rect 4813 -2067 4822 -2033
rect 4856 -2006 4898 -2005
rect 4856 -2040 4861 -2006
rect 4891 -2040 4898 -2006
rect 4856 -2049 4898 -2040
rect 4932 -2006 4974 -1997
rect 4932 -2040 4939 -2006
rect 4969 -2040 4974 -2006
rect 4932 -2045 4974 -2040
rect 5008 -2033 5036 -1973
tri 5081 -1986 5103 -1964 se
rect 5103 -1971 5118 -1963
tri 5103 -1986 5118 -1971 nw
tri 5075 -1992 5081 -1986 se
rect 5081 -1992 5090 -1986
rect 4794 -2077 4822 -2067
tri 4822 -2077 4846 -2053 sw
rect 4794 -2109 4836 -2077
tri 4853 -2085 4854 -2084 sw
rect 4853 -2109 4854 -2085
tri 4856 -2086 4893 -2049 ne
rect 4893 -2077 4898 -2049
tri 4898 -2077 4924 -2051 sw
rect 5008 -2067 5017 -2033
rect 5008 -2077 5036 -2067
rect 4893 -2086 4977 -2077
tri 4893 -2105 4912 -2086 ne
rect 4912 -2105 4977 -2086
rect 4794 -2131 4854 -2109
rect 4976 -2109 4977 -2105
rect 4994 -2109 5036 -2077
rect 4976 -2131 5036 -2109
rect 4882 -2147 4899 -2133
rect 4931 -2147 4948 -2133
rect 5075 -2147 5090 -1992
tri 5090 -1999 5103 -1986 nw
rect 5176 -2067 5191 -1839
rect 5176 -2147 5191 -2109
rect 5219 1984 5234 2174
tri 5299 2138 5321 2160 se
rect 5321 2153 5336 2174
tri 5321 2138 5336 2153 nw
rect 5655 2153 5670 2174
tri 5293 2132 5299 2138 se
rect 5299 2132 5308 2138
rect 5293 2116 5308 2132
tri 5308 2125 5321 2138 nw
rect 5462 2130 5479 2144
rect 5511 2130 5528 2144
tri 5655 2138 5670 2153 ne
tri 5670 2138 5692 2160 sw
rect 5293 2080 5308 2088
rect 5374 2116 5434 2130
rect 5389 2106 5434 2116
rect 5389 2088 5417 2106
tri 5293 2065 5308 2080 ne
tri 5308 2065 5330 2087 sw
rect 5374 2078 5417 2088
rect 5432 2102 5434 2106
rect 5556 2116 5616 2130
tri 5670 2125 5683 2138 ne
rect 5683 2132 5692 2138
tri 5692 2132 5698 2138 sw
rect 5556 2106 5601 2116
rect 5432 2078 5506 2102
rect 5374 2074 5506 2078
tri 5506 2074 5534 2102 sw
rect 5556 2092 5558 2106
tri 5556 2090 5558 2092 ne
rect 5570 2088 5601 2106
rect 5570 2078 5616 2088
rect 5683 2117 5698 2132
tri 5308 2053 5320 2065 ne
rect 5320 2060 5330 2065
tri 5330 2060 5335 2065 sw
rect 5219 1714 5234 1942
rect 5320 1904 5335 2060
rect 5374 2018 5402 2074
tri 5494 2056 5512 2074 ne
rect 5512 2054 5534 2074
tri 5534 2054 5554 2074 sw
tri 5570 2060 5588 2078 ne
rect 5393 1984 5402 2018
rect 5436 2045 5478 2046
rect 5436 2011 5441 2045
rect 5471 2011 5478 2045
rect 5436 2002 5478 2011
rect 5512 2045 5554 2054
rect 5512 2011 5519 2045
rect 5549 2011 5554 2045
rect 5512 2006 5554 2011
rect 5588 2018 5616 2078
tri 5661 2065 5683 2087 se
rect 5683 2080 5698 2088
tri 5683 2065 5698 2080 nw
tri 5655 2059 5661 2065 se
rect 5661 2059 5670 2065
rect 5374 1974 5402 1984
tri 5402 1974 5426 1998 sw
rect 5374 1942 5416 1974
tri 5433 1966 5434 1967 sw
rect 5433 1942 5434 1966
tri 5436 1965 5473 2002 ne
rect 5473 1974 5478 2002
tri 5478 1974 5504 2000 sw
rect 5588 1984 5597 2018
rect 5588 1974 5616 1984
rect 5473 1965 5557 1974
tri 5473 1946 5492 1965 ne
rect 5492 1946 5557 1965
rect 5374 1920 5434 1942
rect 5556 1942 5557 1946
rect 5574 1942 5616 1974
rect 5556 1920 5616 1942
rect 5462 1904 5479 1918
rect 5511 1904 5528 1918
tri 5299 1868 5321 1890 se
rect 5321 1883 5336 1904
tri 5321 1868 5336 1883 nw
rect 5655 1883 5670 2059
tri 5670 2052 5683 2065 nw
rect 5756 1984 5771 2174
tri 5293 1862 5299 1868 se
rect 5299 1862 5308 1868
rect 5293 1846 5308 1862
tri 5308 1855 5321 1868 nw
rect 5462 1860 5479 1874
rect 5511 1860 5528 1874
tri 5655 1868 5670 1883 ne
tri 5670 1868 5692 1890 sw
rect 5293 1810 5308 1818
rect 5374 1846 5434 1860
rect 5389 1836 5434 1846
rect 5389 1818 5417 1836
tri 5293 1795 5308 1810 ne
tri 5308 1795 5330 1817 sw
rect 5374 1808 5417 1818
rect 5432 1832 5434 1836
rect 5556 1846 5616 1860
tri 5670 1855 5683 1868 ne
rect 5683 1862 5692 1868
tri 5692 1862 5698 1868 sw
rect 5556 1836 5601 1846
rect 5432 1808 5506 1832
rect 5374 1804 5506 1808
tri 5506 1804 5534 1832 sw
rect 5556 1822 5558 1836
tri 5556 1820 5558 1822 ne
rect 5570 1818 5601 1836
rect 5570 1808 5616 1818
rect 5683 1847 5698 1862
tri 5308 1783 5320 1795 ne
rect 5320 1790 5330 1795
tri 5330 1790 5335 1795 sw
rect 5219 1444 5234 1672
rect 5320 1682 5335 1790
rect 5374 1748 5402 1804
tri 5494 1786 5512 1804 ne
rect 5512 1784 5534 1804
tri 5534 1784 5554 1804 sw
tri 5570 1790 5588 1808 ne
rect 5393 1714 5402 1748
rect 5436 1775 5478 1776
rect 5436 1741 5441 1775
rect 5471 1741 5478 1775
rect 5436 1732 5478 1741
rect 5512 1775 5554 1784
rect 5512 1741 5519 1775
rect 5549 1741 5554 1775
rect 5512 1736 5554 1741
rect 5588 1748 5616 1808
tri 5661 1795 5683 1817 se
rect 5683 1810 5698 1818
tri 5683 1795 5698 1810 nw
tri 5655 1789 5661 1795 se
rect 5661 1789 5670 1795
rect 5374 1704 5402 1714
tri 5402 1704 5426 1728 sw
rect 5320 1634 5336 1682
rect 5374 1672 5416 1704
tri 5433 1696 5434 1697 sw
rect 5433 1672 5434 1696
tri 5436 1695 5473 1732 ne
rect 5473 1704 5478 1732
tri 5478 1704 5504 1730 sw
rect 5588 1714 5597 1748
rect 5588 1704 5616 1714
rect 5473 1695 5557 1704
tri 5473 1676 5492 1695 ne
rect 5492 1676 5557 1695
rect 5374 1650 5434 1672
rect 5556 1672 5557 1676
rect 5574 1672 5616 1704
rect 5556 1650 5616 1672
rect 5462 1634 5479 1648
rect 5511 1634 5528 1648
tri 5299 1598 5321 1620 se
rect 5321 1613 5336 1634
tri 5321 1598 5336 1613 nw
rect 5655 1613 5670 1789
tri 5670 1782 5683 1795 nw
rect 5756 1714 5771 1942
tri 5293 1592 5299 1598 se
rect 5299 1592 5308 1598
rect 5293 1576 5308 1592
tri 5308 1585 5321 1598 nw
rect 5462 1590 5479 1604
rect 5511 1590 5528 1604
tri 5655 1598 5670 1613 ne
tri 5670 1598 5692 1620 sw
rect 5293 1540 5308 1548
rect 5374 1576 5434 1590
rect 5389 1566 5434 1576
rect 5389 1548 5417 1566
tri 5293 1525 5308 1540 ne
tri 5308 1525 5330 1547 sw
rect 5374 1538 5417 1548
rect 5432 1562 5434 1566
rect 5556 1576 5616 1590
tri 5670 1585 5683 1598 ne
rect 5683 1592 5692 1598
tri 5692 1592 5698 1598 sw
rect 5556 1566 5601 1576
rect 5432 1538 5506 1562
rect 5374 1534 5506 1538
tri 5506 1534 5534 1562 sw
rect 5556 1552 5558 1566
tri 5556 1550 5558 1552 ne
rect 5570 1548 5601 1566
rect 5570 1538 5616 1548
rect 5683 1577 5698 1592
tri 5308 1513 5320 1525 ne
rect 5320 1520 5330 1525
tri 5330 1520 5335 1525 sw
rect 5219 1174 5234 1402
rect 5320 1364 5335 1520
rect 5374 1478 5402 1534
tri 5494 1516 5512 1534 ne
rect 5512 1514 5534 1534
tri 5534 1514 5554 1534 sw
tri 5570 1520 5588 1538 ne
rect 5393 1444 5402 1478
rect 5436 1505 5478 1506
rect 5436 1471 5441 1505
rect 5471 1471 5478 1505
rect 5436 1462 5478 1471
rect 5512 1505 5554 1514
rect 5512 1471 5519 1505
rect 5549 1471 5554 1505
rect 5512 1466 5554 1471
rect 5588 1478 5616 1538
tri 5661 1525 5683 1547 se
rect 5683 1540 5698 1548
tri 5683 1525 5698 1540 nw
tri 5655 1519 5661 1525 se
rect 5661 1519 5670 1525
rect 5374 1434 5402 1444
tri 5402 1434 5426 1458 sw
rect 5374 1402 5416 1434
tri 5433 1426 5434 1427 sw
rect 5433 1402 5434 1426
tri 5436 1425 5473 1462 ne
rect 5473 1434 5478 1462
tri 5478 1434 5504 1460 sw
rect 5588 1444 5597 1478
rect 5588 1434 5616 1444
rect 5473 1425 5557 1434
tri 5473 1406 5492 1425 ne
rect 5492 1406 5557 1425
rect 5374 1380 5434 1402
rect 5556 1402 5557 1406
rect 5574 1402 5616 1434
rect 5556 1380 5616 1402
rect 5462 1364 5479 1378
rect 5511 1364 5528 1378
tri 5299 1328 5321 1350 se
rect 5321 1343 5336 1364
tri 5321 1328 5336 1343 nw
rect 5655 1343 5670 1519
tri 5670 1512 5683 1525 nw
rect 5756 1444 5771 1672
tri 5293 1322 5299 1328 se
rect 5299 1322 5308 1328
rect 5293 1306 5308 1322
tri 5308 1315 5321 1328 nw
rect 5462 1320 5479 1334
rect 5511 1320 5528 1334
tri 5655 1328 5670 1343 ne
tri 5670 1328 5692 1350 sw
rect 5293 1270 5308 1278
rect 5374 1306 5434 1320
rect 5389 1296 5434 1306
rect 5389 1278 5417 1296
tri 5293 1255 5308 1270 ne
tri 5308 1255 5330 1277 sw
rect 5374 1268 5417 1278
rect 5432 1292 5434 1296
rect 5556 1306 5616 1320
tri 5670 1315 5683 1328 ne
rect 5683 1322 5692 1328
tri 5692 1322 5698 1328 sw
rect 5556 1296 5601 1306
rect 5432 1268 5506 1292
rect 5374 1264 5506 1268
tri 5506 1264 5534 1292 sw
rect 5556 1282 5558 1296
tri 5556 1280 5558 1282 ne
rect 5570 1278 5601 1296
rect 5570 1268 5616 1278
rect 5683 1307 5698 1322
tri 5308 1243 5320 1255 ne
rect 5320 1250 5330 1255
tri 5330 1250 5335 1255 sw
rect 5219 903 5234 1132
rect 5320 1141 5335 1250
rect 5374 1208 5402 1264
tri 5494 1246 5512 1264 ne
rect 5512 1244 5534 1264
tri 5534 1244 5554 1264 sw
tri 5570 1250 5588 1268 ne
rect 5393 1174 5402 1208
rect 5436 1235 5478 1236
rect 5436 1201 5441 1235
rect 5471 1201 5478 1235
rect 5436 1192 5478 1201
rect 5512 1235 5554 1244
rect 5512 1201 5519 1235
rect 5549 1201 5554 1235
rect 5512 1196 5554 1201
rect 5588 1208 5616 1268
tri 5661 1255 5683 1277 se
rect 5683 1270 5698 1278
tri 5683 1255 5698 1270 nw
tri 5655 1249 5661 1255 se
rect 5661 1249 5670 1255
rect 5374 1164 5402 1174
tri 5402 1164 5426 1188 sw
rect 5320 1094 5336 1141
rect 5374 1132 5416 1164
tri 5433 1156 5434 1157 sw
rect 5433 1132 5434 1156
tri 5436 1155 5473 1192 ne
rect 5473 1164 5478 1192
tri 5478 1164 5504 1190 sw
rect 5588 1174 5597 1208
rect 5588 1164 5616 1174
rect 5473 1155 5557 1164
tri 5473 1136 5492 1155 ne
rect 5492 1136 5557 1155
rect 5374 1110 5434 1132
rect 5556 1132 5557 1136
rect 5574 1132 5616 1164
rect 5556 1110 5616 1132
rect 5462 1094 5479 1108
rect 5511 1094 5528 1108
tri 5299 1057 5321 1079 se
rect 5321 1072 5336 1094
tri 5321 1057 5336 1072 nw
rect 5655 1072 5670 1249
tri 5670 1242 5683 1255 nw
rect 5756 1174 5771 1402
tri 5293 1051 5299 1057 se
rect 5299 1051 5308 1057
rect 5293 1035 5308 1051
tri 5308 1044 5321 1057 nw
rect 5462 1049 5479 1063
rect 5511 1049 5528 1063
tri 5655 1057 5670 1072 ne
tri 5670 1057 5692 1079 sw
rect 5293 999 5308 1007
rect 5374 1035 5434 1049
rect 5389 1025 5434 1035
rect 5389 1007 5417 1025
tri 5293 984 5308 999 ne
tri 5308 984 5330 1006 sw
rect 5374 997 5417 1007
rect 5432 1021 5434 1025
rect 5556 1035 5616 1049
tri 5670 1044 5683 1057 ne
rect 5683 1051 5692 1057
tri 5692 1051 5698 1057 sw
rect 5556 1025 5601 1035
rect 5432 997 5506 1021
rect 5374 993 5506 997
tri 5506 993 5534 1021 sw
rect 5556 1011 5558 1025
tri 5556 1009 5558 1011 ne
rect 5570 1007 5601 1025
rect 5570 997 5616 1007
rect 5683 1036 5698 1051
tri 5308 972 5320 984 ne
rect 5320 979 5330 984
tri 5330 979 5335 984 sw
rect 5219 633 5234 861
rect 5320 823 5335 979
rect 5374 937 5402 993
tri 5494 975 5512 993 ne
rect 5512 973 5534 993
tri 5534 973 5554 993 sw
tri 5570 979 5588 997 ne
rect 5393 903 5402 937
rect 5436 964 5478 965
rect 5436 930 5441 964
rect 5471 930 5478 964
rect 5436 921 5478 930
rect 5512 964 5554 973
rect 5512 930 5519 964
rect 5549 930 5554 964
rect 5512 925 5554 930
rect 5588 937 5616 997
tri 5661 984 5683 1006 se
rect 5683 999 5698 1007
tri 5683 984 5698 999 nw
tri 5655 978 5661 984 se
rect 5661 978 5670 984
rect 5374 893 5402 903
tri 5402 893 5426 917 sw
rect 5374 861 5416 893
tri 5433 885 5434 886 sw
rect 5433 861 5434 885
tri 5436 884 5473 921 ne
rect 5473 893 5478 921
tri 5478 893 5504 919 sw
rect 5588 903 5597 937
rect 5588 893 5616 903
rect 5473 884 5557 893
tri 5473 865 5492 884 ne
rect 5492 865 5557 884
rect 5374 839 5434 861
rect 5556 861 5557 865
rect 5574 861 5616 893
rect 5556 839 5616 861
rect 5462 823 5479 837
rect 5511 823 5528 837
tri 5299 787 5321 809 se
rect 5321 802 5336 823
tri 5321 787 5336 802 nw
rect 5655 802 5670 978
tri 5670 971 5683 984 nw
rect 5756 903 5771 1132
tri 5293 781 5299 787 se
rect 5299 781 5308 787
rect 5293 765 5308 781
tri 5308 774 5321 787 nw
rect 5462 779 5479 793
rect 5511 779 5528 793
tri 5655 787 5670 802 ne
tri 5670 787 5692 809 sw
rect 5293 729 5308 737
rect 5374 765 5434 779
rect 5389 755 5434 765
rect 5389 737 5417 755
tri 5293 714 5308 729 ne
tri 5308 714 5330 736 sw
rect 5374 727 5417 737
rect 5432 751 5434 755
rect 5556 765 5616 779
tri 5670 774 5683 787 ne
rect 5683 781 5692 787
tri 5692 781 5698 787 sw
rect 5556 755 5601 765
rect 5432 727 5506 751
rect 5374 723 5506 727
tri 5506 723 5534 751 sw
rect 5556 741 5558 755
tri 5556 739 5558 741 ne
rect 5570 737 5601 755
rect 5570 727 5616 737
rect 5683 766 5698 781
tri 5308 702 5320 714 ne
rect 5320 709 5330 714
tri 5330 709 5335 714 sw
rect 5219 363 5234 591
rect 5320 601 5335 709
rect 5374 667 5402 723
tri 5494 705 5512 723 ne
rect 5512 703 5534 723
tri 5534 703 5554 723 sw
tri 5570 709 5588 727 ne
rect 5393 633 5402 667
rect 5436 694 5478 695
rect 5436 660 5441 694
rect 5471 660 5478 694
rect 5436 651 5478 660
rect 5512 694 5554 703
rect 5512 660 5519 694
rect 5549 660 5554 694
rect 5512 655 5554 660
rect 5588 667 5616 727
tri 5661 714 5683 736 se
rect 5683 729 5698 737
tri 5683 714 5698 729 nw
tri 5655 708 5661 714 se
rect 5661 708 5670 714
rect 5374 623 5402 633
tri 5402 623 5426 647 sw
rect 5320 553 5336 601
rect 5374 591 5416 623
tri 5433 615 5434 616 sw
rect 5433 591 5434 615
tri 5436 614 5473 651 ne
rect 5473 623 5478 651
tri 5478 623 5504 649 sw
rect 5588 633 5597 667
rect 5588 623 5616 633
rect 5473 614 5557 623
tri 5473 595 5492 614 ne
rect 5492 595 5557 614
rect 5374 569 5434 591
rect 5556 591 5557 595
rect 5574 591 5616 623
rect 5556 569 5616 591
rect 5462 553 5479 567
rect 5511 553 5528 567
tri 5299 517 5321 539 se
rect 5321 532 5336 553
tri 5321 517 5336 532 nw
rect 5655 532 5670 708
tri 5670 701 5683 714 nw
rect 5756 633 5771 861
tri 5293 511 5299 517 se
rect 5299 511 5308 517
rect 5293 495 5308 511
tri 5308 504 5321 517 nw
rect 5462 509 5479 523
rect 5511 509 5528 523
tri 5655 517 5670 532 ne
tri 5670 517 5692 539 sw
rect 5293 459 5308 467
rect 5374 495 5434 509
rect 5389 485 5434 495
rect 5389 467 5417 485
tri 5293 444 5308 459 ne
tri 5308 444 5330 466 sw
rect 5374 457 5417 467
rect 5432 481 5434 485
rect 5556 495 5616 509
tri 5670 504 5683 517 ne
rect 5683 511 5692 517
tri 5692 511 5698 517 sw
rect 5556 485 5601 495
rect 5432 457 5506 481
rect 5374 453 5506 457
tri 5506 453 5534 481 sw
rect 5556 471 5558 485
tri 5556 469 5558 471 ne
rect 5570 467 5601 485
rect 5570 457 5616 467
rect 5683 496 5698 511
tri 5308 432 5320 444 ne
rect 5320 439 5330 444
tri 5330 439 5335 444 sw
rect 5219 93 5234 321
rect 5320 283 5335 439
rect 5374 397 5402 453
tri 5494 435 5512 453 ne
rect 5512 433 5534 453
tri 5534 433 5554 453 sw
tri 5570 439 5588 457 ne
rect 5393 363 5402 397
rect 5436 424 5478 425
rect 5436 390 5441 424
rect 5471 390 5478 424
rect 5436 381 5478 390
rect 5512 424 5554 433
rect 5512 390 5519 424
rect 5549 390 5554 424
rect 5512 385 5554 390
rect 5588 397 5616 457
tri 5661 444 5683 466 se
rect 5683 459 5698 467
tri 5683 444 5698 459 nw
tri 5655 438 5661 444 se
rect 5661 438 5670 444
rect 5374 353 5402 363
tri 5402 353 5426 377 sw
rect 5374 321 5416 353
tri 5433 345 5434 346 sw
rect 5433 321 5434 345
tri 5436 344 5473 381 ne
rect 5473 353 5478 381
tri 5478 353 5504 379 sw
rect 5588 363 5597 397
rect 5588 353 5616 363
rect 5473 344 5557 353
tri 5473 325 5492 344 ne
rect 5492 325 5557 344
rect 5374 299 5434 321
rect 5556 321 5557 325
rect 5574 321 5616 353
rect 5556 299 5616 321
rect 5462 283 5479 297
rect 5511 283 5528 297
tri 5299 247 5321 269 se
rect 5321 262 5336 283
tri 5321 247 5336 262 nw
rect 5655 262 5670 438
tri 5670 431 5683 444 nw
rect 5756 363 5771 591
tri 5293 241 5299 247 se
rect 5299 241 5308 247
rect 5293 225 5308 241
tri 5308 234 5321 247 nw
rect 5462 239 5479 253
rect 5511 239 5528 253
tri 5655 247 5670 262 ne
tri 5670 247 5692 269 sw
rect 5293 189 5308 197
rect 5374 225 5434 239
rect 5389 215 5434 225
rect 5389 197 5417 215
tri 5293 174 5308 189 ne
tri 5308 174 5330 196 sw
rect 5374 187 5417 197
rect 5432 211 5434 215
rect 5556 225 5616 239
tri 5670 234 5683 247 ne
rect 5683 241 5692 247
tri 5692 241 5698 247 sw
rect 5556 215 5601 225
rect 5432 187 5506 211
rect 5374 183 5506 187
tri 5506 183 5534 211 sw
rect 5556 201 5558 215
tri 5556 199 5558 201 ne
rect 5570 197 5601 215
rect 5570 187 5616 197
rect 5683 226 5698 241
tri 5308 162 5320 174 ne
rect 5320 169 5330 174
tri 5330 169 5335 174 sw
rect 5219 -177 5234 51
rect 5320 61 5335 169
rect 5374 127 5402 183
tri 5494 165 5512 183 ne
rect 5512 163 5534 183
tri 5534 163 5554 183 sw
tri 5570 169 5588 187 ne
rect 5393 93 5402 127
rect 5436 154 5478 155
rect 5436 120 5441 154
rect 5471 120 5478 154
rect 5436 111 5478 120
rect 5512 154 5554 163
rect 5512 120 5519 154
rect 5549 120 5554 154
rect 5512 115 5554 120
rect 5588 127 5616 187
tri 5661 174 5683 196 se
rect 5683 189 5698 197
tri 5683 174 5698 189 nw
tri 5655 168 5661 174 se
rect 5661 168 5670 174
rect 5374 83 5402 93
tri 5402 83 5426 107 sw
rect 5320 13 5336 61
rect 5374 51 5416 83
tri 5433 75 5434 76 sw
rect 5433 51 5434 75
tri 5436 74 5473 111 ne
rect 5473 83 5478 111
tri 5478 83 5504 109 sw
rect 5588 93 5597 127
rect 5588 83 5616 93
rect 5473 74 5557 83
tri 5473 55 5492 74 ne
rect 5492 55 5557 74
rect 5374 29 5434 51
rect 5556 51 5557 55
rect 5574 51 5616 83
rect 5556 29 5616 51
rect 5462 13 5479 27
rect 5511 13 5528 27
tri 5299 -23 5321 -1 se
rect 5321 -8 5336 13
tri 5321 -23 5336 -8 nw
rect 5655 -8 5670 168
tri 5670 161 5683 174 nw
rect 5756 93 5771 321
tri 5293 -29 5299 -23 se
rect 5299 -29 5308 -23
rect 5293 -45 5308 -29
tri 5308 -36 5321 -23 nw
rect 5462 -31 5479 -17
rect 5511 -31 5528 -17
tri 5655 -23 5670 -8 ne
tri 5670 -23 5692 -1 sw
rect 5293 -81 5308 -73
rect 5374 -45 5434 -31
rect 5389 -55 5434 -45
rect 5389 -73 5417 -55
tri 5293 -96 5308 -81 ne
tri 5308 -96 5330 -74 sw
rect 5374 -83 5417 -73
rect 5432 -59 5434 -55
rect 5556 -45 5616 -31
tri 5670 -36 5683 -23 ne
rect 5683 -29 5692 -23
tri 5692 -29 5698 -23 sw
rect 5556 -55 5601 -45
rect 5432 -83 5506 -59
rect 5374 -87 5506 -83
tri 5506 -87 5534 -59 sw
rect 5556 -69 5558 -55
tri 5556 -71 5558 -69 ne
rect 5570 -73 5601 -55
rect 5570 -83 5616 -73
rect 5683 -44 5698 -29
tri 5308 -108 5320 -96 ne
rect 5320 -101 5330 -96
tri 5330 -101 5335 -96 sw
rect 5219 -447 5234 -219
rect 5320 -257 5335 -101
rect 5374 -143 5402 -87
tri 5494 -105 5512 -87 ne
rect 5512 -107 5534 -87
tri 5534 -107 5554 -87 sw
tri 5570 -101 5588 -83 ne
rect 5393 -177 5402 -143
rect 5436 -116 5478 -115
rect 5436 -150 5441 -116
rect 5471 -150 5478 -116
rect 5436 -159 5478 -150
rect 5512 -116 5554 -107
rect 5512 -150 5519 -116
rect 5549 -150 5554 -116
rect 5512 -155 5554 -150
rect 5588 -143 5616 -83
tri 5661 -96 5683 -74 se
rect 5683 -81 5698 -73
tri 5683 -96 5698 -81 nw
tri 5655 -102 5661 -96 se
rect 5661 -102 5670 -96
rect 5374 -187 5402 -177
tri 5402 -187 5426 -163 sw
rect 5374 -219 5416 -187
tri 5433 -195 5434 -194 sw
rect 5433 -219 5434 -195
tri 5436 -196 5473 -159 ne
rect 5473 -187 5478 -159
tri 5478 -187 5504 -161 sw
rect 5588 -177 5597 -143
rect 5588 -187 5616 -177
rect 5473 -196 5557 -187
tri 5473 -215 5492 -196 ne
rect 5492 -215 5557 -196
rect 5374 -241 5434 -219
rect 5556 -219 5557 -215
rect 5574 -219 5616 -187
rect 5556 -241 5616 -219
rect 5462 -257 5479 -243
rect 5511 -257 5528 -243
tri 5299 -293 5321 -271 se
rect 5321 -278 5336 -257
tri 5321 -293 5336 -278 nw
rect 5655 -278 5670 -102
tri 5670 -109 5683 -96 nw
rect 5756 -177 5771 51
tri 5293 -299 5299 -293 se
rect 5299 -299 5308 -293
rect 5293 -315 5308 -299
tri 5308 -306 5321 -293 nw
rect 5462 -301 5479 -287
rect 5511 -301 5528 -287
tri 5655 -293 5670 -278 ne
tri 5670 -293 5692 -271 sw
rect 5293 -351 5308 -343
rect 5374 -315 5434 -301
rect 5389 -325 5434 -315
rect 5389 -343 5417 -325
tri 5293 -366 5308 -351 ne
tri 5308 -366 5330 -344 sw
rect 5374 -353 5417 -343
rect 5432 -329 5434 -325
rect 5556 -315 5616 -301
tri 5670 -306 5683 -293 ne
rect 5683 -299 5692 -293
tri 5692 -299 5698 -293 sw
rect 5556 -325 5601 -315
rect 5432 -353 5506 -329
rect 5374 -357 5506 -353
tri 5506 -357 5534 -329 sw
rect 5556 -339 5558 -325
tri 5556 -341 5558 -339 ne
rect 5570 -343 5601 -325
rect 5570 -353 5616 -343
rect 5683 -314 5698 -299
tri 5308 -378 5320 -366 ne
rect 5320 -371 5330 -366
tri 5330 -371 5335 -366 sw
rect 5219 -717 5234 -489
rect 5320 -479 5335 -371
rect 5374 -413 5402 -357
tri 5494 -375 5512 -357 ne
rect 5512 -377 5534 -357
tri 5534 -377 5554 -357 sw
tri 5570 -371 5588 -353 ne
rect 5393 -447 5402 -413
rect 5436 -386 5478 -385
rect 5436 -420 5441 -386
rect 5471 -420 5478 -386
rect 5436 -429 5478 -420
rect 5512 -386 5554 -377
rect 5512 -420 5519 -386
rect 5549 -420 5554 -386
rect 5512 -425 5554 -420
rect 5588 -413 5616 -353
tri 5661 -366 5683 -344 se
rect 5683 -351 5698 -343
tri 5683 -366 5698 -351 nw
tri 5655 -372 5661 -366 se
rect 5661 -372 5670 -366
rect 5374 -457 5402 -447
tri 5402 -457 5426 -433 sw
rect 5320 -527 5336 -479
rect 5374 -489 5416 -457
tri 5433 -465 5434 -464 sw
rect 5433 -489 5434 -465
tri 5436 -466 5473 -429 ne
rect 5473 -457 5478 -429
tri 5478 -457 5504 -431 sw
rect 5588 -447 5597 -413
rect 5588 -457 5616 -447
rect 5473 -466 5557 -457
tri 5473 -485 5492 -466 ne
rect 5492 -485 5557 -466
rect 5374 -511 5434 -489
rect 5556 -489 5557 -485
rect 5574 -489 5616 -457
rect 5556 -511 5616 -489
rect 5462 -527 5479 -513
rect 5511 -527 5528 -513
tri 5299 -563 5321 -541 se
rect 5321 -548 5336 -527
tri 5321 -563 5336 -548 nw
rect 5655 -548 5670 -372
tri 5670 -379 5683 -366 nw
rect 5756 -447 5771 -219
tri 5293 -569 5299 -563 se
rect 5299 -569 5308 -563
rect 5293 -585 5308 -569
tri 5308 -576 5321 -563 nw
rect 5462 -571 5479 -557
rect 5511 -571 5528 -557
tri 5655 -563 5670 -548 ne
tri 5670 -563 5692 -541 sw
rect 5293 -621 5308 -613
rect 5374 -585 5434 -571
rect 5389 -595 5434 -585
rect 5389 -613 5417 -595
tri 5293 -636 5308 -621 ne
tri 5308 -636 5330 -614 sw
rect 5374 -623 5417 -613
rect 5432 -599 5434 -595
rect 5556 -585 5616 -571
tri 5670 -576 5683 -563 ne
rect 5683 -569 5692 -563
tri 5692 -569 5698 -563 sw
rect 5556 -595 5601 -585
rect 5432 -623 5506 -599
rect 5374 -627 5506 -623
tri 5506 -627 5534 -599 sw
rect 5556 -609 5558 -595
tri 5556 -611 5558 -609 ne
rect 5570 -613 5601 -595
rect 5570 -623 5616 -613
rect 5683 -584 5698 -569
tri 5308 -648 5320 -636 ne
rect 5320 -641 5330 -636
tri 5330 -641 5335 -636 sw
rect 5219 -987 5234 -759
rect 5320 -797 5335 -641
rect 5374 -683 5402 -627
tri 5494 -645 5512 -627 ne
rect 5512 -647 5534 -627
tri 5534 -647 5554 -627 sw
tri 5570 -641 5588 -623 ne
rect 5393 -717 5402 -683
rect 5436 -656 5478 -655
rect 5436 -690 5441 -656
rect 5471 -690 5478 -656
rect 5436 -699 5478 -690
rect 5512 -656 5554 -647
rect 5512 -690 5519 -656
rect 5549 -690 5554 -656
rect 5512 -695 5554 -690
rect 5588 -683 5616 -623
tri 5661 -636 5683 -614 se
rect 5683 -621 5698 -613
tri 5683 -636 5698 -621 nw
tri 5655 -642 5661 -636 se
rect 5661 -642 5670 -636
rect 5374 -727 5402 -717
tri 5402 -727 5426 -703 sw
rect 5374 -759 5416 -727
tri 5433 -735 5434 -734 sw
rect 5433 -759 5434 -735
tri 5436 -736 5473 -699 ne
rect 5473 -727 5478 -699
tri 5478 -727 5504 -701 sw
rect 5588 -717 5597 -683
rect 5588 -727 5616 -717
rect 5473 -736 5557 -727
tri 5473 -755 5492 -736 ne
rect 5492 -755 5557 -736
rect 5374 -781 5434 -759
rect 5556 -759 5557 -755
rect 5574 -759 5616 -727
rect 5556 -781 5616 -759
rect 5462 -797 5479 -783
rect 5511 -797 5528 -783
tri 5299 -833 5321 -811 se
rect 5321 -818 5336 -797
tri 5321 -833 5336 -818 nw
rect 5655 -818 5670 -642
tri 5670 -649 5683 -636 nw
rect 5756 -717 5771 -489
tri 5293 -839 5299 -833 se
rect 5299 -839 5308 -833
rect 5293 -855 5308 -839
tri 5308 -846 5321 -833 nw
rect 5462 -841 5479 -827
rect 5511 -841 5528 -827
tri 5655 -833 5670 -818 ne
tri 5670 -833 5692 -811 sw
rect 5293 -891 5308 -883
rect 5374 -855 5434 -841
rect 5389 -865 5434 -855
rect 5389 -883 5417 -865
tri 5293 -906 5308 -891 ne
tri 5308 -906 5330 -884 sw
rect 5374 -893 5417 -883
rect 5432 -869 5434 -865
rect 5556 -855 5616 -841
tri 5670 -846 5683 -833 ne
rect 5683 -839 5692 -833
tri 5692 -839 5698 -833 sw
rect 5556 -865 5601 -855
rect 5432 -893 5506 -869
rect 5374 -897 5506 -893
tri 5506 -897 5534 -869 sw
rect 5556 -879 5558 -865
tri 5556 -881 5558 -879 ne
rect 5570 -883 5601 -865
rect 5570 -893 5616 -883
rect 5683 -854 5698 -839
tri 5308 -918 5320 -906 ne
rect 5320 -911 5330 -906
tri 5330 -911 5335 -906 sw
rect 5219 -1257 5234 -1029
rect 5320 -1019 5335 -911
rect 5374 -953 5402 -897
tri 5494 -915 5512 -897 ne
rect 5512 -917 5534 -897
tri 5534 -917 5554 -897 sw
tri 5570 -911 5588 -893 ne
rect 5393 -987 5402 -953
rect 5436 -926 5478 -925
rect 5436 -960 5441 -926
rect 5471 -960 5478 -926
rect 5436 -969 5478 -960
rect 5512 -926 5554 -917
rect 5512 -960 5519 -926
rect 5549 -960 5554 -926
rect 5512 -965 5554 -960
rect 5588 -953 5616 -893
tri 5661 -906 5683 -884 se
rect 5683 -891 5698 -883
tri 5683 -906 5698 -891 nw
tri 5655 -912 5661 -906 se
rect 5661 -912 5670 -906
rect 5374 -997 5402 -987
tri 5402 -997 5426 -973 sw
rect 5320 -1067 5336 -1019
rect 5374 -1029 5416 -997
tri 5433 -1005 5434 -1004 sw
rect 5433 -1029 5434 -1005
tri 5436 -1006 5473 -969 ne
rect 5473 -997 5478 -969
tri 5478 -997 5504 -971 sw
rect 5588 -987 5597 -953
rect 5588 -997 5616 -987
rect 5473 -1006 5557 -997
tri 5473 -1025 5492 -1006 ne
rect 5492 -1025 5557 -1006
rect 5374 -1051 5434 -1029
rect 5556 -1029 5557 -1025
rect 5574 -1029 5616 -997
rect 5556 -1051 5616 -1029
rect 5462 -1067 5479 -1053
rect 5511 -1067 5528 -1053
tri 5299 -1103 5321 -1081 se
rect 5321 -1088 5336 -1067
tri 5321 -1103 5336 -1088 nw
rect 5655 -1088 5670 -912
tri 5670 -919 5683 -906 nw
rect 5756 -987 5771 -759
tri 5293 -1109 5299 -1103 se
rect 5299 -1109 5308 -1103
rect 5293 -1125 5308 -1109
tri 5308 -1116 5321 -1103 nw
rect 5462 -1111 5479 -1097
rect 5511 -1111 5528 -1097
tri 5655 -1103 5670 -1088 ne
tri 5670 -1103 5692 -1081 sw
rect 5293 -1161 5308 -1153
rect 5374 -1125 5434 -1111
rect 5389 -1135 5434 -1125
rect 5389 -1153 5417 -1135
tri 5293 -1176 5308 -1161 ne
tri 5308 -1176 5330 -1154 sw
rect 5374 -1163 5417 -1153
rect 5432 -1139 5434 -1135
rect 5556 -1125 5616 -1111
tri 5670 -1116 5683 -1103 ne
rect 5683 -1109 5692 -1103
tri 5692 -1109 5698 -1103 sw
rect 5556 -1135 5601 -1125
rect 5432 -1163 5506 -1139
rect 5374 -1167 5506 -1163
tri 5506 -1167 5534 -1139 sw
rect 5556 -1149 5558 -1135
tri 5556 -1151 5558 -1149 ne
rect 5570 -1153 5601 -1135
rect 5570 -1163 5616 -1153
rect 5683 -1124 5698 -1109
tri 5308 -1188 5320 -1176 ne
rect 5320 -1181 5330 -1176
tri 5330 -1181 5335 -1176 sw
rect 5219 -1527 5234 -1299
rect 5320 -1337 5335 -1181
rect 5374 -1223 5402 -1167
tri 5494 -1185 5512 -1167 ne
rect 5512 -1187 5534 -1167
tri 5534 -1187 5554 -1167 sw
tri 5570 -1181 5588 -1163 ne
rect 5393 -1257 5402 -1223
rect 5436 -1196 5478 -1195
rect 5436 -1230 5441 -1196
rect 5471 -1230 5478 -1196
rect 5436 -1239 5478 -1230
rect 5512 -1196 5554 -1187
rect 5512 -1230 5519 -1196
rect 5549 -1230 5554 -1196
rect 5512 -1235 5554 -1230
rect 5588 -1223 5616 -1163
tri 5661 -1176 5683 -1154 se
rect 5683 -1161 5698 -1153
tri 5683 -1176 5698 -1161 nw
tri 5655 -1182 5661 -1176 se
rect 5661 -1182 5670 -1176
rect 5374 -1267 5402 -1257
tri 5402 -1267 5426 -1243 sw
rect 5374 -1299 5416 -1267
tri 5433 -1275 5434 -1274 sw
rect 5433 -1299 5434 -1275
tri 5436 -1276 5473 -1239 ne
rect 5473 -1267 5478 -1239
tri 5478 -1267 5504 -1241 sw
rect 5588 -1257 5597 -1223
rect 5588 -1267 5616 -1257
rect 5473 -1276 5557 -1267
tri 5473 -1295 5492 -1276 ne
rect 5492 -1295 5557 -1276
rect 5374 -1321 5434 -1299
rect 5556 -1299 5557 -1295
rect 5574 -1299 5616 -1267
rect 5556 -1321 5616 -1299
rect 5462 -1337 5479 -1323
rect 5511 -1337 5528 -1323
tri 5299 -1373 5321 -1351 se
rect 5321 -1358 5336 -1337
tri 5321 -1373 5336 -1358 nw
rect 5655 -1358 5670 -1182
tri 5670 -1189 5683 -1176 nw
rect 5756 -1257 5771 -1029
tri 5293 -1379 5299 -1373 se
rect 5299 -1379 5308 -1373
rect 5293 -1395 5308 -1379
tri 5308 -1386 5321 -1373 nw
rect 5462 -1381 5479 -1367
rect 5511 -1381 5528 -1367
tri 5655 -1373 5670 -1358 ne
tri 5670 -1373 5692 -1351 sw
rect 5293 -1431 5308 -1423
rect 5374 -1395 5434 -1381
rect 5389 -1405 5434 -1395
rect 5389 -1423 5417 -1405
tri 5293 -1446 5308 -1431 ne
tri 5308 -1446 5330 -1424 sw
rect 5374 -1433 5417 -1423
rect 5432 -1409 5434 -1405
rect 5556 -1395 5616 -1381
tri 5670 -1386 5683 -1373 ne
rect 5683 -1379 5692 -1373
tri 5692 -1379 5698 -1373 sw
rect 5556 -1405 5601 -1395
rect 5432 -1433 5506 -1409
rect 5374 -1437 5506 -1433
tri 5506 -1437 5534 -1409 sw
rect 5556 -1419 5558 -1405
tri 5556 -1421 5558 -1419 ne
rect 5570 -1423 5601 -1405
rect 5570 -1433 5616 -1423
rect 5683 -1394 5698 -1379
tri 5308 -1458 5320 -1446 ne
rect 5320 -1451 5330 -1446
tri 5330 -1451 5335 -1446 sw
rect 5219 -1797 5234 -1569
rect 5320 -1559 5335 -1451
rect 5374 -1493 5402 -1437
tri 5494 -1455 5512 -1437 ne
rect 5512 -1457 5534 -1437
tri 5534 -1457 5554 -1437 sw
tri 5570 -1451 5588 -1433 ne
rect 5393 -1527 5402 -1493
rect 5436 -1466 5478 -1465
rect 5436 -1500 5441 -1466
rect 5471 -1500 5478 -1466
rect 5436 -1509 5478 -1500
rect 5512 -1466 5554 -1457
rect 5512 -1500 5519 -1466
rect 5549 -1500 5554 -1466
rect 5512 -1505 5554 -1500
rect 5588 -1493 5616 -1433
tri 5661 -1446 5683 -1424 se
rect 5683 -1431 5698 -1423
tri 5683 -1446 5698 -1431 nw
tri 5655 -1452 5661 -1446 se
rect 5661 -1452 5670 -1446
rect 5374 -1537 5402 -1527
tri 5402 -1537 5426 -1513 sw
rect 5320 -1607 5336 -1559
rect 5374 -1569 5416 -1537
tri 5433 -1545 5434 -1544 sw
rect 5433 -1569 5434 -1545
tri 5436 -1546 5473 -1509 ne
rect 5473 -1537 5478 -1509
tri 5478 -1537 5504 -1511 sw
rect 5588 -1527 5597 -1493
rect 5588 -1537 5616 -1527
rect 5473 -1546 5557 -1537
tri 5473 -1565 5492 -1546 ne
rect 5492 -1565 5557 -1546
rect 5374 -1591 5434 -1569
rect 5556 -1569 5557 -1565
rect 5574 -1569 5616 -1537
rect 5556 -1591 5616 -1569
rect 5462 -1607 5479 -1593
rect 5511 -1607 5528 -1593
tri 5299 -1643 5321 -1621 se
rect 5321 -1628 5336 -1607
tri 5321 -1643 5336 -1628 nw
rect 5655 -1628 5670 -1452
tri 5670 -1459 5683 -1446 nw
rect 5756 -1527 5771 -1299
tri 5293 -1649 5299 -1643 se
rect 5299 -1649 5308 -1643
rect 5293 -1665 5308 -1649
tri 5308 -1656 5321 -1643 nw
rect 5462 -1651 5479 -1637
rect 5511 -1651 5528 -1637
tri 5655 -1643 5670 -1628 ne
tri 5670 -1643 5692 -1621 sw
rect 5293 -1701 5308 -1693
rect 5374 -1665 5434 -1651
rect 5389 -1675 5434 -1665
rect 5389 -1693 5417 -1675
tri 5293 -1716 5308 -1701 ne
tri 5308 -1716 5330 -1694 sw
rect 5374 -1703 5417 -1693
rect 5432 -1679 5434 -1675
rect 5556 -1665 5616 -1651
tri 5670 -1656 5683 -1643 ne
rect 5683 -1649 5692 -1643
tri 5692 -1649 5698 -1643 sw
rect 5556 -1675 5601 -1665
rect 5432 -1703 5506 -1679
rect 5374 -1707 5506 -1703
tri 5506 -1707 5534 -1679 sw
rect 5556 -1689 5558 -1675
tri 5556 -1691 5558 -1689 ne
rect 5570 -1693 5601 -1675
rect 5570 -1703 5616 -1693
rect 5683 -1664 5698 -1649
tri 5308 -1728 5320 -1716 ne
rect 5320 -1721 5330 -1716
tri 5330 -1721 5335 -1716 sw
rect 5219 -2067 5234 -1839
rect 5320 -1877 5335 -1721
rect 5374 -1763 5402 -1707
tri 5494 -1725 5512 -1707 ne
rect 5512 -1727 5534 -1707
tri 5534 -1727 5554 -1707 sw
tri 5570 -1721 5588 -1703 ne
rect 5393 -1797 5402 -1763
rect 5436 -1736 5478 -1735
rect 5436 -1770 5441 -1736
rect 5471 -1770 5478 -1736
rect 5436 -1779 5478 -1770
rect 5512 -1736 5554 -1727
rect 5512 -1770 5519 -1736
rect 5549 -1770 5554 -1736
rect 5512 -1775 5554 -1770
rect 5588 -1763 5616 -1703
tri 5661 -1716 5683 -1694 se
rect 5683 -1701 5698 -1693
tri 5683 -1716 5698 -1701 nw
tri 5655 -1722 5661 -1716 se
rect 5661 -1722 5670 -1716
rect 5374 -1807 5402 -1797
tri 5402 -1807 5426 -1783 sw
rect 5374 -1839 5416 -1807
tri 5433 -1815 5434 -1814 sw
rect 5433 -1839 5434 -1815
tri 5436 -1816 5473 -1779 ne
rect 5473 -1807 5478 -1779
tri 5478 -1807 5504 -1781 sw
rect 5588 -1797 5597 -1763
rect 5588 -1807 5616 -1797
rect 5473 -1816 5557 -1807
tri 5473 -1835 5492 -1816 ne
rect 5492 -1835 5557 -1816
rect 5374 -1861 5434 -1839
rect 5556 -1839 5557 -1835
rect 5574 -1839 5616 -1807
rect 5556 -1861 5616 -1839
rect 5462 -1877 5479 -1863
rect 5511 -1877 5528 -1863
tri 5299 -1913 5321 -1891 se
rect 5321 -1898 5336 -1877
tri 5321 -1913 5336 -1898 nw
rect 5655 -1898 5670 -1722
tri 5670 -1729 5683 -1716 nw
rect 5756 -1797 5771 -1569
tri 5293 -1919 5299 -1913 se
rect 5299 -1919 5308 -1913
rect 5293 -1935 5308 -1919
tri 5308 -1926 5321 -1913 nw
rect 5462 -1921 5479 -1907
rect 5511 -1921 5528 -1907
tri 5655 -1913 5670 -1898 ne
tri 5670 -1913 5692 -1891 sw
rect 5293 -1971 5308 -1963
rect 5374 -1935 5434 -1921
rect 5389 -1945 5434 -1935
rect 5389 -1963 5417 -1945
tri 5293 -1986 5308 -1971 ne
tri 5308 -1986 5330 -1964 sw
rect 5374 -1973 5417 -1963
rect 5432 -1949 5434 -1945
rect 5556 -1935 5616 -1921
tri 5670 -1926 5683 -1913 ne
rect 5683 -1919 5692 -1913
tri 5692 -1919 5698 -1913 sw
rect 5556 -1945 5601 -1935
rect 5432 -1973 5506 -1949
rect 5374 -1977 5506 -1973
tri 5506 -1977 5534 -1949 sw
rect 5556 -1959 5558 -1945
tri 5556 -1961 5558 -1959 ne
rect 5570 -1963 5601 -1945
rect 5570 -1973 5616 -1963
rect 5683 -1934 5698 -1919
tri 5308 -1998 5320 -1986 ne
rect 5320 -1991 5330 -1986
tri 5330 -1991 5335 -1986 sw
rect 5219 -2147 5234 -2109
rect 5320 -2147 5335 -1991
rect 5374 -2033 5402 -1977
tri 5494 -1995 5512 -1977 ne
rect 5512 -1997 5534 -1977
tri 5534 -1997 5554 -1977 sw
tri 5570 -1991 5588 -1973 ne
rect 5393 -2067 5402 -2033
rect 5436 -2006 5478 -2005
rect 5436 -2040 5441 -2006
rect 5471 -2040 5478 -2006
rect 5436 -2049 5478 -2040
rect 5512 -2006 5554 -1997
rect 5512 -2040 5519 -2006
rect 5549 -2040 5554 -2006
rect 5512 -2045 5554 -2040
rect 5588 -2033 5616 -1973
tri 5661 -1986 5683 -1964 se
rect 5683 -1971 5698 -1963
tri 5683 -1986 5698 -1971 nw
tri 5655 -1992 5661 -1986 se
rect 5661 -1992 5670 -1986
rect 5374 -2077 5402 -2067
tri 5402 -2077 5426 -2053 sw
rect 5374 -2109 5416 -2077
tri 5433 -2085 5434 -2084 sw
rect 5433 -2109 5434 -2085
tri 5436 -2086 5473 -2049 ne
rect 5473 -2077 5478 -2049
tri 5478 -2077 5504 -2051 sw
rect 5588 -2067 5597 -2033
rect 5588 -2077 5616 -2067
rect 5473 -2086 5557 -2077
tri 5473 -2105 5492 -2086 ne
rect 5492 -2105 5557 -2086
rect 5374 -2131 5434 -2109
rect 5556 -2109 5557 -2105
rect 5574 -2109 5616 -2077
rect 5556 -2131 5616 -2109
rect 5462 -2147 5479 -2133
rect 5511 -2147 5528 -2133
rect 5655 -2147 5670 -1992
tri 5670 -1999 5683 -1986 nw
rect 5756 -2067 5771 -1839
rect 5756 -2147 5771 -2109
rect 5799 1984 5814 2174
tri 5879 2138 5901 2160 se
rect 5901 2153 5916 2174
tri 5901 2138 5916 2153 nw
rect 6235 2153 6250 2174
tri 5873 2132 5879 2138 se
rect 5879 2132 5888 2138
rect 5873 2116 5888 2132
tri 5888 2125 5901 2138 nw
rect 6042 2130 6059 2144
rect 6091 2130 6108 2144
tri 6235 2138 6250 2153 ne
tri 6250 2138 6272 2160 sw
rect 5873 2080 5888 2088
rect 5954 2116 6014 2130
rect 5969 2106 6014 2116
rect 5969 2088 5997 2106
tri 5873 2065 5888 2080 ne
tri 5888 2065 5910 2087 sw
rect 5954 2078 5997 2088
rect 6012 2102 6014 2106
rect 6136 2116 6196 2130
tri 6250 2125 6263 2138 ne
rect 6263 2132 6272 2138
tri 6272 2132 6278 2138 sw
rect 6136 2106 6181 2116
rect 6012 2078 6086 2102
rect 5954 2074 6086 2078
tri 6086 2074 6114 2102 sw
rect 6136 2092 6138 2106
tri 6136 2090 6138 2092 ne
rect 6150 2088 6181 2106
rect 6150 2078 6196 2088
rect 6263 2117 6278 2132
tri 5888 2053 5900 2065 ne
rect 5900 2060 5910 2065
tri 5910 2060 5915 2065 sw
rect 5799 1714 5814 1942
rect 5900 1904 5915 2060
rect 5954 2018 5982 2074
tri 6074 2056 6092 2074 ne
rect 6092 2054 6114 2074
tri 6114 2054 6134 2074 sw
tri 6150 2060 6168 2078 ne
rect 5973 1984 5982 2018
rect 6016 2045 6058 2046
rect 6016 2011 6021 2045
rect 6051 2011 6058 2045
rect 6016 2002 6058 2011
rect 6092 2045 6134 2054
rect 6092 2011 6099 2045
rect 6129 2011 6134 2045
rect 6092 2006 6134 2011
rect 6168 2018 6196 2078
tri 6241 2065 6263 2087 se
rect 6263 2080 6278 2088
tri 6263 2065 6278 2080 nw
tri 6235 2059 6241 2065 se
rect 6241 2059 6250 2065
rect 5954 1974 5982 1984
tri 5982 1974 6006 1998 sw
rect 5954 1942 5996 1974
tri 6013 1966 6014 1967 sw
rect 6013 1942 6014 1966
tri 6016 1965 6053 2002 ne
rect 6053 1974 6058 2002
tri 6058 1974 6084 2000 sw
rect 6168 1984 6177 2018
rect 6168 1974 6196 1984
rect 6053 1965 6137 1974
tri 6053 1946 6072 1965 ne
rect 6072 1946 6137 1965
rect 5954 1920 6014 1942
rect 6136 1942 6137 1946
rect 6154 1942 6196 1974
rect 6136 1920 6196 1942
rect 6042 1904 6059 1918
rect 6091 1904 6108 1918
tri 5879 1868 5901 1890 se
rect 5901 1883 5916 1904
tri 5901 1868 5916 1883 nw
rect 6235 1883 6250 2059
tri 6250 2052 6263 2065 nw
rect 6336 1984 6351 2174
tri 5873 1862 5879 1868 se
rect 5879 1862 5888 1868
rect 5873 1846 5888 1862
tri 5888 1855 5901 1868 nw
rect 6042 1860 6059 1874
rect 6091 1860 6108 1874
tri 6235 1868 6250 1883 ne
tri 6250 1868 6272 1890 sw
rect 5873 1810 5888 1818
rect 5954 1846 6014 1860
rect 5969 1836 6014 1846
rect 5969 1818 5997 1836
tri 5873 1795 5888 1810 ne
tri 5888 1795 5910 1817 sw
rect 5954 1808 5997 1818
rect 6012 1832 6014 1836
rect 6136 1846 6196 1860
tri 6250 1855 6263 1868 ne
rect 6263 1862 6272 1868
tri 6272 1862 6278 1868 sw
rect 6136 1836 6181 1846
rect 6012 1808 6086 1832
rect 5954 1804 6086 1808
tri 6086 1804 6114 1832 sw
rect 6136 1822 6138 1836
tri 6136 1820 6138 1822 ne
rect 6150 1818 6181 1836
rect 6150 1808 6196 1818
rect 6263 1847 6278 1862
tri 5888 1783 5900 1795 ne
rect 5900 1790 5910 1795
tri 5910 1790 5915 1795 sw
rect 5799 1444 5814 1672
rect 5900 1682 5915 1790
rect 5954 1748 5982 1804
tri 6074 1786 6092 1804 ne
rect 6092 1784 6114 1804
tri 6114 1784 6134 1804 sw
tri 6150 1790 6168 1808 ne
rect 5973 1714 5982 1748
rect 6016 1775 6058 1776
rect 6016 1741 6021 1775
rect 6051 1741 6058 1775
rect 6016 1732 6058 1741
rect 6092 1775 6134 1784
rect 6092 1741 6099 1775
rect 6129 1741 6134 1775
rect 6092 1736 6134 1741
rect 6168 1748 6196 1808
tri 6241 1795 6263 1817 se
rect 6263 1810 6278 1818
tri 6263 1795 6278 1810 nw
tri 6235 1789 6241 1795 se
rect 6241 1789 6250 1795
rect 5954 1704 5982 1714
tri 5982 1704 6006 1728 sw
rect 5900 1634 5916 1682
rect 5954 1672 5996 1704
tri 6013 1696 6014 1697 sw
rect 6013 1672 6014 1696
tri 6016 1695 6053 1732 ne
rect 6053 1704 6058 1732
tri 6058 1704 6084 1730 sw
rect 6168 1714 6177 1748
rect 6168 1704 6196 1714
rect 6053 1695 6137 1704
tri 6053 1676 6072 1695 ne
rect 6072 1676 6137 1695
rect 5954 1650 6014 1672
rect 6136 1672 6137 1676
rect 6154 1672 6196 1704
rect 6136 1650 6196 1672
rect 6042 1634 6059 1648
rect 6091 1634 6108 1648
tri 5879 1598 5901 1620 se
rect 5901 1613 5916 1634
tri 5901 1598 5916 1613 nw
rect 6235 1613 6250 1789
tri 6250 1782 6263 1795 nw
rect 6336 1714 6351 1942
tri 5873 1592 5879 1598 se
rect 5879 1592 5888 1598
rect 5873 1576 5888 1592
tri 5888 1585 5901 1598 nw
rect 6042 1590 6059 1604
rect 6091 1590 6108 1604
tri 6235 1598 6250 1613 ne
tri 6250 1598 6272 1620 sw
rect 5873 1540 5888 1548
rect 5954 1576 6014 1590
rect 5969 1566 6014 1576
rect 5969 1548 5997 1566
tri 5873 1525 5888 1540 ne
tri 5888 1525 5910 1547 sw
rect 5954 1538 5997 1548
rect 6012 1562 6014 1566
rect 6136 1576 6196 1590
tri 6250 1585 6263 1598 ne
rect 6263 1592 6272 1598
tri 6272 1592 6278 1598 sw
rect 6136 1566 6181 1576
rect 6012 1538 6086 1562
rect 5954 1534 6086 1538
tri 6086 1534 6114 1562 sw
rect 6136 1552 6138 1566
tri 6136 1550 6138 1552 ne
rect 6150 1548 6181 1566
rect 6150 1538 6196 1548
rect 6263 1577 6278 1592
tri 5888 1513 5900 1525 ne
rect 5900 1520 5910 1525
tri 5910 1520 5915 1525 sw
rect 5799 1174 5814 1402
rect 5900 1364 5915 1520
rect 5954 1478 5982 1534
tri 6074 1516 6092 1534 ne
rect 6092 1514 6114 1534
tri 6114 1514 6134 1534 sw
tri 6150 1520 6168 1538 ne
rect 5973 1444 5982 1478
rect 6016 1505 6058 1506
rect 6016 1471 6021 1505
rect 6051 1471 6058 1505
rect 6016 1462 6058 1471
rect 6092 1505 6134 1514
rect 6092 1471 6099 1505
rect 6129 1471 6134 1505
rect 6092 1466 6134 1471
rect 6168 1478 6196 1538
tri 6241 1525 6263 1547 se
rect 6263 1540 6278 1548
tri 6263 1525 6278 1540 nw
tri 6235 1519 6241 1525 se
rect 6241 1519 6250 1525
rect 5954 1434 5982 1444
tri 5982 1434 6006 1458 sw
rect 5954 1402 5996 1434
tri 6013 1426 6014 1427 sw
rect 6013 1402 6014 1426
tri 6016 1425 6053 1462 ne
rect 6053 1434 6058 1462
tri 6058 1434 6084 1460 sw
rect 6168 1444 6177 1478
rect 6168 1434 6196 1444
rect 6053 1425 6137 1434
tri 6053 1406 6072 1425 ne
rect 6072 1406 6137 1425
rect 5954 1380 6014 1402
rect 6136 1402 6137 1406
rect 6154 1402 6196 1434
rect 6136 1380 6196 1402
rect 6042 1364 6059 1378
rect 6091 1364 6108 1378
tri 5879 1328 5901 1350 se
rect 5901 1343 5916 1364
tri 5901 1328 5916 1343 nw
rect 6235 1343 6250 1519
tri 6250 1512 6263 1525 nw
rect 6336 1444 6351 1672
tri 5873 1322 5879 1328 se
rect 5879 1322 5888 1328
rect 5873 1306 5888 1322
tri 5888 1315 5901 1328 nw
rect 6042 1320 6059 1334
rect 6091 1320 6108 1334
tri 6235 1328 6250 1343 ne
tri 6250 1328 6272 1350 sw
rect 5873 1270 5888 1278
rect 5954 1306 6014 1320
rect 5969 1296 6014 1306
rect 5969 1278 5997 1296
tri 5873 1255 5888 1270 ne
tri 5888 1255 5910 1277 sw
rect 5954 1268 5997 1278
rect 6012 1292 6014 1296
rect 6136 1306 6196 1320
tri 6250 1315 6263 1328 ne
rect 6263 1322 6272 1328
tri 6272 1322 6278 1328 sw
rect 6136 1296 6181 1306
rect 6012 1268 6086 1292
rect 5954 1264 6086 1268
tri 6086 1264 6114 1292 sw
rect 6136 1282 6138 1296
tri 6136 1280 6138 1282 ne
rect 6150 1278 6181 1296
rect 6150 1268 6196 1278
rect 6263 1307 6278 1322
tri 5888 1243 5900 1255 ne
rect 5900 1250 5910 1255
tri 5910 1250 5915 1255 sw
rect 5799 903 5814 1132
rect 5900 1141 5915 1250
rect 5954 1208 5982 1264
tri 6074 1246 6092 1264 ne
rect 6092 1244 6114 1264
tri 6114 1244 6134 1264 sw
tri 6150 1250 6168 1268 ne
rect 5973 1174 5982 1208
rect 6016 1235 6058 1236
rect 6016 1201 6021 1235
rect 6051 1201 6058 1235
rect 6016 1192 6058 1201
rect 6092 1235 6134 1244
rect 6092 1201 6099 1235
rect 6129 1201 6134 1235
rect 6092 1196 6134 1201
rect 6168 1208 6196 1268
tri 6241 1255 6263 1277 se
rect 6263 1270 6278 1278
tri 6263 1255 6278 1270 nw
tri 6235 1249 6241 1255 se
rect 6241 1249 6250 1255
rect 5954 1164 5982 1174
tri 5982 1164 6006 1188 sw
rect 5900 1094 5916 1141
rect 5954 1132 5996 1164
tri 6013 1156 6014 1157 sw
rect 6013 1132 6014 1156
tri 6016 1155 6053 1192 ne
rect 6053 1164 6058 1192
tri 6058 1164 6084 1190 sw
rect 6168 1174 6177 1208
rect 6168 1164 6196 1174
rect 6053 1155 6137 1164
tri 6053 1136 6072 1155 ne
rect 6072 1136 6137 1155
rect 5954 1110 6014 1132
rect 6136 1132 6137 1136
rect 6154 1132 6196 1164
rect 6136 1110 6196 1132
rect 6042 1094 6059 1108
rect 6091 1094 6108 1108
tri 5879 1057 5901 1079 se
rect 5901 1072 5916 1094
tri 5901 1057 5916 1072 nw
rect 6235 1072 6250 1249
tri 6250 1242 6263 1255 nw
rect 6336 1174 6351 1402
tri 5873 1051 5879 1057 se
rect 5879 1051 5888 1057
rect 5873 1035 5888 1051
tri 5888 1044 5901 1057 nw
rect 6042 1049 6059 1063
rect 6091 1049 6108 1063
tri 6235 1057 6250 1072 ne
tri 6250 1057 6272 1079 sw
rect 5873 999 5888 1007
rect 5954 1035 6014 1049
rect 5969 1025 6014 1035
rect 5969 1007 5997 1025
tri 5873 984 5888 999 ne
tri 5888 984 5910 1006 sw
rect 5954 997 5997 1007
rect 6012 1021 6014 1025
rect 6136 1035 6196 1049
tri 6250 1044 6263 1057 ne
rect 6263 1051 6272 1057
tri 6272 1051 6278 1057 sw
rect 6136 1025 6181 1035
rect 6012 997 6086 1021
rect 5954 993 6086 997
tri 6086 993 6114 1021 sw
rect 6136 1011 6138 1025
tri 6136 1009 6138 1011 ne
rect 6150 1007 6181 1025
rect 6150 997 6196 1007
rect 6263 1036 6278 1051
tri 5888 972 5900 984 ne
rect 5900 979 5910 984
tri 5910 979 5915 984 sw
rect 5799 633 5814 861
rect 5900 823 5915 979
rect 5954 937 5982 993
tri 6074 975 6092 993 ne
rect 6092 973 6114 993
tri 6114 973 6134 993 sw
tri 6150 979 6168 997 ne
rect 5973 903 5982 937
rect 6016 964 6058 965
rect 6016 930 6021 964
rect 6051 930 6058 964
rect 6016 921 6058 930
rect 6092 964 6134 973
rect 6092 930 6099 964
rect 6129 930 6134 964
rect 6092 925 6134 930
rect 6168 937 6196 997
tri 6241 984 6263 1006 se
rect 6263 999 6278 1007
tri 6263 984 6278 999 nw
tri 6235 978 6241 984 se
rect 6241 978 6250 984
rect 5954 893 5982 903
tri 5982 893 6006 917 sw
rect 5954 861 5996 893
tri 6013 885 6014 886 sw
rect 6013 861 6014 885
tri 6016 884 6053 921 ne
rect 6053 893 6058 921
tri 6058 893 6084 919 sw
rect 6168 903 6177 937
rect 6168 893 6196 903
rect 6053 884 6137 893
tri 6053 865 6072 884 ne
rect 6072 865 6137 884
rect 5954 839 6014 861
rect 6136 861 6137 865
rect 6154 861 6196 893
rect 6136 839 6196 861
rect 6042 823 6059 837
rect 6091 823 6108 837
tri 5879 787 5901 809 se
rect 5901 802 5916 823
tri 5901 787 5916 802 nw
rect 6235 802 6250 978
tri 6250 971 6263 984 nw
rect 6336 903 6351 1132
tri 5873 781 5879 787 se
rect 5879 781 5888 787
rect 5873 765 5888 781
tri 5888 774 5901 787 nw
rect 6042 779 6059 793
rect 6091 779 6108 793
tri 6235 787 6250 802 ne
tri 6250 787 6272 809 sw
rect 5873 729 5888 737
rect 5954 765 6014 779
rect 5969 755 6014 765
rect 5969 737 5997 755
tri 5873 714 5888 729 ne
tri 5888 714 5910 736 sw
rect 5954 727 5997 737
rect 6012 751 6014 755
rect 6136 765 6196 779
tri 6250 774 6263 787 ne
rect 6263 781 6272 787
tri 6272 781 6278 787 sw
rect 6136 755 6181 765
rect 6012 727 6086 751
rect 5954 723 6086 727
tri 6086 723 6114 751 sw
rect 6136 741 6138 755
tri 6136 739 6138 741 ne
rect 6150 737 6181 755
rect 6150 727 6196 737
rect 6263 766 6278 781
tri 5888 702 5900 714 ne
rect 5900 709 5910 714
tri 5910 709 5915 714 sw
rect 5799 363 5814 591
rect 5900 601 5915 709
rect 5954 667 5982 723
tri 6074 705 6092 723 ne
rect 6092 703 6114 723
tri 6114 703 6134 723 sw
tri 6150 709 6168 727 ne
rect 5973 633 5982 667
rect 6016 694 6058 695
rect 6016 660 6021 694
rect 6051 660 6058 694
rect 6016 651 6058 660
rect 6092 694 6134 703
rect 6092 660 6099 694
rect 6129 660 6134 694
rect 6092 655 6134 660
rect 6168 667 6196 727
tri 6241 714 6263 736 se
rect 6263 729 6278 737
tri 6263 714 6278 729 nw
tri 6235 708 6241 714 se
rect 6241 708 6250 714
rect 5954 623 5982 633
tri 5982 623 6006 647 sw
rect 5900 553 5916 601
rect 5954 591 5996 623
tri 6013 615 6014 616 sw
rect 6013 591 6014 615
tri 6016 614 6053 651 ne
rect 6053 623 6058 651
tri 6058 623 6084 649 sw
rect 6168 633 6177 667
rect 6168 623 6196 633
rect 6053 614 6137 623
tri 6053 595 6072 614 ne
rect 6072 595 6137 614
rect 5954 569 6014 591
rect 6136 591 6137 595
rect 6154 591 6196 623
rect 6136 569 6196 591
rect 6042 553 6059 567
rect 6091 553 6108 567
tri 5879 517 5901 539 se
rect 5901 532 5916 553
tri 5901 517 5916 532 nw
rect 6235 532 6250 708
tri 6250 701 6263 714 nw
rect 6336 633 6351 861
tri 5873 511 5879 517 se
rect 5879 511 5888 517
rect 5873 495 5888 511
tri 5888 504 5901 517 nw
rect 6042 509 6059 523
rect 6091 509 6108 523
tri 6235 517 6250 532 ne
tri 6250 517 6272 539 sw
rect 5873 459 5888 467
rect 5954 495 6014 509
rect 5969 485 6014 495
rect 5969 467 5997 485
tri 5873 444 5888 459 ne
tri 5888 444 5910 466 sw
rect 5954 457 5997 467
rect 6012 481 6014 485
rect 6136 495 6196 509
tri 6250 504 6263 517 ne
rect 6263 511 6272 517
tri 6272 511 6278 517 sw
rect 6136 485 6181 495
rect 6012 457 6086 481
rect 5954 453 6086 457
tri 6086 453 6114 481 sw
rect 6136 471 6138 485
tri 6136 469 6138 471 ne
rect 6150 467 6181 485
rect 6150 457 6196 467
rect 6263 496 6278 511
tri 5888 432 5900 444 ne
rect 5900 439 5910 444
tri 5910 439 5915 444 sw
rect 5799 93 5814 321
rect 5900 283 5915 439
rect 5954 397 5982 453
tri 6074 435 6092 453 ne
rect 6092 433 6114 453
tri 6114 433 6134 453 sw
tri 6150 439 6168 457 ne
rect 5973 363 5982 397
rect 6016 424 6058 425
rect 6016 390 6021 424
rect 6051 390 6058 424
rect 6016 381 6058 390
rect 6092 424 6134 433
rect 6092 390 6099 424
rect 6129 390 6134 424
rect 6092 385 6134 390
rect 6168 397 6196 457
tri 6241 444 6263 466 se
rect 6263 459 6278 467
tri 6263 444 6278 459 nw
tri 6235 438 6241 444 se
rect 6241 438 6250 444
rect 5954 353 5982 363
tri 5982 353 6006 377 sw
rect 5954 321 5996 353
tri 6013 345 6014 346 sw
rect 6013 321 6014 345
tri 6016 344 6053 381 ne
rect 6053 353 6058 381
tri 6058 353 6084 379 sw
rect 6168 363 6177 397
rect 6168 353 6196 363
rect 6053 344 6137 353
tri 6053 325 6072 344 ne
rect 6072 325 6137 344
rect 5954 299 6014 321
rect 6136 321 6137 325
rect 6154 321 6196 353
rect 6136 299 6196 321
rect 6042 283 6059 297
rect 6091 283 6108 297
tri 5879 247 5901 269 se
rect 5901 262 5916 283
tri 5901 247 5916 262 nw
rect 6235 262 6250 438
tri 6250 431 6263 444 nw
rect 6336 363 6351 591
tri 5873 241 5879 247 se
rect 5879 241 5888 247
rect 5873 225 5888 241
tri 5888 234 5901 247 nw
rect 6042 239 6059 253
rect 6091 239 6108 253
tri 6235 247 6250 262 ne
tri 6250 247 6272 269 sw
rect 5873 189 5888 197
rect 5954 225 6014 239
rect 5969 215 6014 225
rect 5969 197 5997 215
tri 5873 174 5888 189 ne
tri 5888 174 5910 196 sw
rect 5954 187 5997 197
rect 6012 211 6014 215
rect 6136 225 6196 239
tri 6250 234 6263 247 ne
rect 6263 241 6272 247
tri 6272 241 6278 247 sw
rect 6136 215 6181 225
rect 6012 187 6086 211
rect 5954 183 6086 187
tri 6086 183 6114 211 sw
rect 6136 201 6138 215
tri 6136 199 6138 201 ne
rect 6150 197 6181 215
rect 6150 187 6196 197
rect 6263 226 6278 241
tri 5888 162 5900 174 ne
rect 5900 169 5910 174
tri 5910 169 5915 174 sw
rect 5799 -177 5814 51
rect 5900 61 5915 169
rect 5954 127 5982 183
tri 6074 165 6092 183 ne
rect 6092 163 6114 183
tri 6114 163 6134 183 sw
tri 6150 169 6168 187 ne
rect 5973 93 5982 127
rect 6016 154 6058 155
rect 6016 120 6021 154
rect 6051 120 6058 154
rect 6016 111 6058 120
rect 6092 154 6134 163
rect 6092 120 6099 154
rect 6129 120 6134 154
rect 6092 115 6134 120
rect 6168 127 6196 187
tri 6241 174 6263 196 se
rect 6263 189 6278 197
tri 6263 174 6278 189 nw
tri 6235 168 6241 174 se
rect 6241 168 6250 174
rect 5954 83 5982 93
tri 5982 83 6006 107 sw
rect 5900 13 5916 61
rect 5954 51 5996 83
tri 6013 75 6014 76 sw
rect 6013 51 6014 75
tri 6016 74 6053 111 ne
rect 6053 83 6058 111
tri 6058 83 6084 109 sw
rect 6168 93 6177 127
rect 6168 83 6196 93
rect 6053 74 6137 83
tri 6053 55 6072 74 ne
rect 6072 55 6137 74
rect 5954 29 6014 51
rect 6136 51 6137 55
rect 6154 51 6196 83
rect 6136 29 6196 51
rect 6042 13 6059 27
rect 6091 13 6108 27
tri 5879 -23 5901 -1 se
rect 5901 -8 5916 13
tri 5901 -23 5916 -8 nw
rect 6235 -8 6250 168
tri 6250 161 6263 174 nw
rect 6336 93 6351 321
tri 5873 -29 5879 -23 se
rect 5879 -29 5888 -23
rect 5873 -45 5888 -29
tri 5888 -36 5901 -23 nw
rect 6042 -31 6059 -17
rect 6091 -31 6108 -17
tri 6235 -23 6250 -8 ne
tri 6250 -23 6272 -1 sw
rect 5873 -81 5888 -73
rect 5954 -45 6014 -31
rect 5969 -55 6014 -45
rect 5969 -73 5997 -55
tri 5873 -96 5888 -81 ne
tri 5888 -96 5910 -74 sw
rect 5954 -83 5997 -73
rect 6012 -59 6014 -55
rect 6136 -45 6196 -31
tri 6250 -36 6263 -23 ne
rect 6263 -29 6272 -23
tri 6272 -29 6278 -23 sw
rect 6136 -55 6181 -45
rect 6012 -83 6086 -59
rect 5954 -87 6086 -83
tri 6086 -87 6114 -59 sw
rect 6136 -69 6138 -55
tri 6136 -71 6138 -69 ne
rect 6150 -73 6181 -55
rect 6150 -83 6196 -73
rect 6263 -44 6278 -29
tri 5888 -108 5900 -96 ne
rect 5900 -101 5910 -96
tri 5910 -101 5915 -96 sw
rect 5799 -447 5814 -219
rect 5900 -257 5915 -101
rect 5954 -143 5982 -87
tri 6074 -105 6092 -87 ne
rect 6092 -107 6114 -87
tri 6114 -107 6134 -87 sw
tri 6150 -101 6168 -83 ne
rect 5973 -177 5982 -143
rect 6016 -116 6058 -115
rect 6016 -150 6021 -116
rect 6051 -150 6058 -116
rect 6016 -159 6058 -150
rect 6092 -116 6134 -107
rect 6092 -150 6099 -116
rect 6129 -150 6134 -116
rect 6092 -155 6134 -150
rect 6168 -143 6196 -83
tri 6241 -96 6263 -74 se
rect 6263 -81 6278 -73
tri 6263 -96 6278 -81 nw
tri 6235 -102 6241 -96 se
rect 6241 -102 6250 -96
rect 5954 -187 5982 -177
tri 5982 -187 6006 -163 sw
rect 5954 -219 5996 -187
tri 6013 -195 6014 -194 sw
rect 6013 -219 6014 -195
tri 6016 -196 6053 -159 ne
rect 6053 -187 6058 -159
tri 6058 -187 6084 -161 sw
rect 6168 -177 6177 -143
rect 6168 -187 6196 -177
rect 6053 -196 6137 -187
tri 6053 -215 6072 -196 ne
rect 6072 -215 6137 -196
rect 5954 -241 6014 -219
rect 6136 -219 6137 -215
rect 6154 -219 6196 -187
rect 6136 -241 6196 -219
rect 6042 -257 6059 -243
rect 6091 -257 6108 -243
tri 5879 -293 5901 -271 se
rect 5901 -278 5916 -257
tri 5901 -293 5916 -278 nw
rect 6235 -278 6250 -102
tri 6250 -109 6263 -96 nw
rect 6336 -177 6351 51
tri 5873 -299 5879 -293 se
rect 5879 -299 5888 -293
rect 5873 -315 5888 -299
tri 5888 -306 5901 -293 nw
rect 6042 -301 6059 -287
rect 6091 -301 6108 -287
tri 6235 -293 6250 -278 ne
tri 6250 -293 6272 -271 sw
rect 5873 -351 5888 -343
rect 5954 -315 6014 -301
rect 5969 -325 6014 -315
rect 5969 -343 5997 -325
tri 5873 -366 5888 -351 ne
tri 5888 -366 5910 -344 sw
rect 5954 -353 5997 -343
rect 6012 -329 6014 -325
rect 6136 -315 6196 -301
tri 6250 -306 6263 -293 ne
rect 6263 -299 6272 -293
tri 6272 -299 6278 -293 sw
rect 6136 -325 6181 -315
rect 6012 -353 6086 -329
rect 5954 -357 6086 -353
tri 6086 -357 6114 -329 sw
rect 6136 -339 6138 -325
tri 6136 -341 6138 -339 ne
rect 6150 -343 6181 -325
rect 6150 -353 6196 -343
rect 6263 -314 6278 -299
tri 5888 -378 5900 -366 ne
rect 5900 -371 5910 -366
tri 5910 -371 5915 -366 sw
rect 5799 -717 5814 -489
rect 5900 -479 5915 -371
rect 5954 -413 5982 -357
tri 6074 -375 6092 -357 ne
rect 6092 -377 6114 -357
tri 6114 -377 6134 -357 sw
tri 6150 -371 6168 -353 ne
rect 5973 -447 5982 -413
rect 6016 -386 6058 -385
rect 6016 -420 6021 -386
rect 6051 -420 6058 -386
rect 6016 -429 6058 -420
rect 6092 -386 6134 -377
rect 6092 -420 6099 -386
rect 6129 -420 6134 -386
rect 6092 -425 6134 -420
rect 6168 -413 6196 -353
tri 6241 -366 6263 -344 se
rect 6263 -351 6278 -343
tri 6263 -366 6278 -351 nw
tri 6235 -372 6241 -366 se
rect 6241 -372 6250 -366
rect 5954 -457 5982 -447
tri 5982 -457 6006 -433 sw
rect 5900 -527 5916 -479
rect 5954 -489 5996 -457
tri 6013 -465 6014 -464 sw
rect 6013 -489 6014 -465
tri 6016 -466 6053 -429 ne
rect 6053 -457 6058 -429
tri 6058 -457 6084 -431 sw
rect 6168 -447 6177 -413
rect 6168 -457 6196 -447
rect 6053 -466 6137 -457
tri 6053 -485 6072 -466 ne
rect 6072 -485 6137 -466
rect 5954 -511 6014 -489
rect 6136 -489 6137 -485
rect 6154 -489 6196 -457
rect 6136 -511 6196 -489
rect 6042 -527 6059 -513
rect 6091 -527 6108 -513
tri 5879 -563 5901 -541 se
rect 5901 -548 5916 -527
tri 5901 -563 5916 -548 nw
rect 6235 -548 6250 -372
tri 6250 -379 6263 -366 nw
rect 6336 -447 6351 -219
tri 5873 -569 5879 -563 se
rect 5879 -569 5888 -563
rect 5873 -585 5888 -569
tri 5888 -576 5901 -563 nw
rect 6042 -571 6059 -557
rect 6091 -571 6108 -557
tri 6235 -563 6250 -548 ne
tri 6250 -563 6272 -541 sw
rect 5873 -621 5888 -613
rect 5954 -585 6014 -571
rect 5969 -595 6014 -585
rect 5969 -613 5997 -595
tri 5873 -636 5888 -621 ne
tri 5888 -636 5910 -614 sw
rect 5954 -623 5997 -613
rect 6012 -599 6014 -595
rect 6136 -585 6196 -571
tri 6250 -576 6263 -563 ne
rect 6263 -569 6272 -563
tri 6272 -569 6278 -563 sw
rect 6136 -595 6181 -585
rect 6012 -623 6086 -599
rect 5954 -627 6086 -623
tri 6086 -627 6114 -599 sw
rect 6136 -609 6138 -595
tri 6136 -611 6138 -609 ne
rect 6150 -613 6181 -595
rect 6150 -623 6196 -613
rect 6263 -584 6278 -569
tri 5888 -648 5900 -636 ne
rect 5900 -641 5910 -636
tri 5910 -641 5915 -636 sw
rect 5799 -987 5814 -759
rect 5900 -797 5915 -641
rect 5954 -683 5982 -627
tri 6074 -645 6092 -627 ne
rect 6092 -647 6114 -627
tri 6114 -647 6134 -627 sw
tri 6150 -641 6168 -623 ne
rect 5973 -717 5982 -683
rect 6016 -656 6058 -655
rect 6016 -690 6021 -656
rect 6051 -690 6058 -656
rect 6016 -699 6058 -690
rect 6092 -656 6134 -647
rect 6092 -690 6099 -656
rect 6129 -690 6134 -656
rect 6092 -695 6134 -690
rect 6168 -683 6196 -623
tri 6241 -636 6263 -614 se
rect 6263 -621 6278 -613
tri 6263 -636 6278 -621 nw
tri 6235 -642 6241 -636 se
rect 6241 -642 6250 -636
rect 5954 -727 5982 -717
tri 5982 -727 6006 -703 sw
rect 5954 -759 5996 -727
tri 6013 -735 6014 -734 sw
rect 6013 -759 6014 -735
tri 6016 -736 6053 -699 ne
rect 6053 -727 6058 -699
tri 6058 -727 6084 -701 sw
rect 6168 -717 6177 -683
rect 6168 -727 6196 -717
rect 6053 -736 6137 -727
tri 6053 -755 6072 -736 ne
rect 6072 -755 6137 -736
rect 5954 -781 6014 -759
rect 6136 -759 6137 -755
rect 6154 -759 6196 -727
rect 6136 -781 6196 -759
rect 6042 -797 6059 -783
rect 6091 -797 6108 -783
tri 5879 -833 5901 -811 se
rect 5901 -818 5916 -797
tri 5901 -833 5916 -818 nw
rect 6235 -818 6250 -642
tri 6250 -649 6263 -636 nw
rect 6336 -717 6351 -489
tri 5873 -839 5879 -833 se
rect 5879 -839 5888 -833
rect 5873 -855 5888 -839
tri 5888 -846 5901 -833 nw
rect 6042 -841 6059 -827
rect 6091 -841 6108 -827
tri 6235 -833 6250 -818 ne
tri 6250 -833 6272 -811 sw
rect 5873 -891 5888 -883
rect 5954 -855 6014 -841
rect 5969 -865 6014 -855
rect 5969 -883 5997 -865
tri 5873 -906 5888 -891 ne
tri 5888 -906 5910 -884 sw
rect 5954 -893 5997 -883
rect 6012 -869 6014 -865
rect 6136 -855 6196 -841
tri 6250 -846 6263 -833 ne
rect 6263 -839 6272 -833
tri 6272 -839 6278 -833 sw
rect 6136 -865 6181 -855
rect 6012 -893 6086 -869
rect 5954 -897 6086 -893
tri 6086 -897 6114 -869 sw
rect 6136 -879 6138 -865
tri 6136 -881 6138 -879 ne
rect 6150 -883 6181 -865
rect 6150 -893 6196 -883
rect 6263 -854 6278 -839
tri 5888 -918 5900 -906 ne
rect 5900 -911 5910 -906
tri 5910 -911 5915 -906 sw
rect 5799 -1257 5814 -1029
rect 5900 -1019 5915 -911
rect 5954 -953 5982 -897
tri 6074 -915 6092 -897 ne
rect 6092 -917 6114 -897
tri 6114 -917 6134 -897 sw
tri 6150 -911 6168 -893 ne
rect 5973 -987 5982 -953
rect 6016 -926 6058 -925
rect 6016 -960 6021 -926
rect 6051 -960 6058 -926
rect 6016 -969 6058 -960
rect 6092 -926 6134 -917
rect 6092 -960 6099 -926
rect 6129 -960 6134 -926
rect 6092 -965 6134 -960
rect 6168 -953 6196 -893
tri 6241 -906 6263 -884 se
rect 6263 -891 6278 -883
tri 6263 -906 6278 -891 nw
tri 6235 -912 6241 -906 se
rect 6241 -912 6250 -906
rect 5954 -997 5982 -987
tri 5982 -997 6006 -973 sw
rect 5900 -1067 5916 -1019
rect 5954 -1029 5996 -997
tri 6013 -1005 6014 -1004 sw
rect 6013 -1029 6014 -1005
tri 6016 -1006 6053 -969 ne
rect 6053 -997 6058 -969
tri 6058 -997 6084 -971 sw
rect 6168 -987 6177 -953
rect 6168 -997 6196 -987
rect 6053 -1006 6137 -997
tri 6053 -1025 6072 -1006 ne
rect 6072 -1025 6137 -1006
rect 5954 -1051 6014 -1029
rect 6136 -1029 6137 -1025
rect 6154 -1029 6196 -997
rect 6136 -1051 6196 -1029
rect 6042 -1067 6059 -1053
rect 6091 -1067 6108 -1053
tri 5879 -1103 5901 -1081 se
rect 5901 -1088 5916 -1067
tri 5901 -1103 5916 -1088 nw
rect 6235 -1088 6250 -912
tri 6250 -919 6263 -906 nw
rect 6336 -987 6351 -759
tri 5873 -1109 5879 -1103 se
rect 5879 -1109 5888 -1103
rect 5873 -1125 5888 -1109
tri 5888 -1116 5901 -1103 nw
rect 6042 -1111 6059 -1097
rect 6091 -1111 6108 -1097
tri 6235 -1103 6250 -1088 ne
tri 6250 -1103 6272 -1081 sw
rect 5873 -1161 5888 -1153
rect 5954 -1125 6014 -1111
rect 5969 -1135 6014 -1125
rect 5969 -1153 5997 -1135
tri 5873 -1176 5888 -1161 ne
tri 5888 -1176 5910 -1154 sw
rect 5954 -1163 5997 -1153
rect 6012 -1139 6014 -1135
rect 6136 -1125 6196 -1111
tri 6250 -1116 6263 -1103 ne
rect 6263 -1109 6272 -1103
tri 6272 -1109 6278 -1103 sw
rect 6136 -1135 6181 -1125
rect 6012 -1163 6086 -1139
rect 5954 -1167 6086 -1163
tri 6086 -1167 6114 -1139 sw
rect 6136 -1149 6138 -1135
tri 6136 -1151 6138 -1149 ne
rect 6150 -1153 6181 -1135
rect 6150 -1163 6196 -1153
rect 6263 -1124 6278 -1109
tri 5888 -1188 5900 -1176 ne
rect 5900 -1181 5910 -1176
tri 5910 -1181 5915 -1176 sw
rect 5799 -1527 5814 -1299
rect 5900 -1337 5915 -1181
rect 5954 -1223 5982 -1167
tri 6074 -1185 6092 -1167 ne
rect 6092 -1187 6114 -1167
tri 6114 -1187 6134 -1167 sw
tri 6150 -1181 6168 -1163 ne
rect 5973 -1257 5982 -1223
rect 6016 -1196 6058 -1195
rect 6016 -1230 6021 -1196
rect 6051 -1230 6058 -1196
rect 6016 -1239 6058 -1230
rect 6092 -1196 6134 -1187
rect 6092 -1230 6099 -1196
rect 6129 -1230 6134 -1196
rect 6092 -1235 6134 -1230
rect 6168 -1223 6196 -1163
tri 6241 -1176 6263 -1154 se
rect 6263 -1161 6278 -1153
tri 6263 -1176 6278 -1161 nw
tri 6235 -1182 6241 -1176 se
rect 6241 -1182 6250 -1176
rect 5954 -1267 5982 -1257
tri 5982 -1267 6006 -1243 sw
rect 5954 -1299 5996 -1267
tri 6013 -1275 6014 -1274 sw
rect 6013 -1299 6014 -1275
tri 6016 -1276 6053 -1239 ne
rect 6053 -1267 6058 -1239
tri 6058 -1267 6084 -1241 sw
rect 6168 -1257 6177 -1223
rect 6168 -1267 6196 -1257
rect 6053 -1276 6137 -1267
tri 6053 -1295 6072 -1276 ne
rect 6072 -1295 6137 -1276
rect 5954 -1321 6014 -1299
rect 6136 -1299 6137 -1295
rect 6154 -1299 6196 -1267
rect 6136 -1321 6196 -1299
rect 6042 -1337 6059 -1323
rect 6091 -1337 6108 -1323
tri 5879 -1373 5901 -1351 se
rect 5901 -1358 5916 -1337
tri 5901 -1373 5916 -1358 nw
rect 6235 -1358 6250 -1182
tri 6250 -1189 6263 -1176 nw
rect 6336 -1257 6351 -1029
tri 5873 -1379 5879 -1373 se
rect 5879 -1379 5888 -1373
rect 5873 -1395 5888 -1379
tri 5888 -1386 5901 -1373 nw
rect 6042 -1381 6059 -1367
rect 6091 -1381 6108 -1367
tri 6235 -1373 6250 -1358 ne
tri 6250 -1373 6272 -1351 sw
rect 5873 -1431 5888 -1423
rect 5954 -1395 6014 -1381
rect 5969 -1405 6014 -1395
rect 5969 -1423 5997 -1405
tri 5873 -1446 5888 -1431 ne
tri 5888 -1446 5910 -1424 sw
rect 5954 -1433 5997 -1423
rect 6012 -1409 6014 -1405
rect 6136 -1395 6196 -1381
tri 6250 -1386 6263 -1373 ne
rect 6263 -1379 6272 -1373
tri 6272 -1379 6278 -1373 sw
rect 6136 -1405 6181 -1395
rect 6012 -1433 6086 -1409
rect 5954 -1437 6086 -1433
tri 6086 -1437 6114 -1409 sw
rect 6136 -1419 6138 -1405
tri 6136 -1421 6138 -1419 ne
rect 6150 -1423 6181 -1405
rect 6150 -1433 6196 -1423
rect 6263 -1394 6278 -1379
tri 5888 -1458 5900 -1446 ne
rect 5900 -1451 5910 -1446
tri 5910 -1451 5915 -1446 sw
rect 5799 -1797 5814 -1569
rect 5900 -1559 5915 -1451
rect 5954 -1493 5982 -1437
tri 6074 -1455 6092 -1437 ne
rect 6092 -1457 6114 -1437
tri 6114 -1457 6134 -1437 sw
tri 6150 -1451 6168 -1433 ne
rect 5973 -1527 5982 -1493
rect 6016 -1466 6058 -1465
rect 6016 -1500 6021 -1466
rect 6051 -1500 6058 -1466
rect 6016 -1509 6058 -1500
rect 6092 -1466 6134 -1457
rect 6092 -1500 6099 -1466
rect 6129 -1500 6134 -1466
rect 6092 -1505 6134 -1500
rect 6168 -1493 6196 -1433
tri 6241 -1446 6263 -1424 se
rect 6263 -1431 6278 -1423
tri 6263 -1446 6278 -1431 nw
tri 6235 -1452 6241 -1446 se
rect 6241 -1452 6250 -1446
rect 5954 -1537 5982 -1527
tri 5982 -1537 6006 -1513 sw
rect 5900 -1607 5916 -1559
rect 5954 -1569 5996 -1537
tri 6013 -1545 6014 -1544 sw
rect 6013 -1569 6014 -1545
tri 6016 -1546 6053 -1509 ne
rect 6053 -1537 6058 -1509
tri 6058 -1537 6084 -1511 sw
rect 6168 -1527 6177 -1493
rect 6168 -1537 6196 -1527
rect 6053 -1546 6137 -1537
tri 6053 -1565 6072 -1546 ne
rect 6072 -1565 6137 -1546
rect 5954 -1591 6014 -1569
rect 6136 -1569 6137 -1565
rect 6154 -1569 6196 -1537
rect 6136 -1591 6196 -1569
rect 6042 -1607 6059 -1593
rect 6091 -1607 6108 -1593
tri 5879 -1643 5901 -1621 se
rect 5901 -1628 5916 -1607
tri 5901 -1643 5916 -1628 nw
rect 6235 -1628 6250 -1452
tri 6250 -1459 6263 -1446 nw
rect 6336 -1527 6351 -1299
tri 5873 -1649 5879 -1643 se
rect 5879 -1649 5888 -1643
rect 5873 -1665 5888 -1649
tri 5888 -1656 5901 -1643 nw
rect 6042 -1651 6059 -1637
rect 6091 -1651 6108 -1637
tri 6235 -1643 6250 -1628 ne
tri 6250 -1643 6272 -1621 sw
rect 5873 -1701 5888 -1693
rect 5954 -1665 6014 -1651
rect 5969 -1675 6014 -1665
rect 5969 -1693 5997 -1675
tri 5873 -1716 5888 -1701 ne
tri 5888 -1716 5910 -1694 sw
rect 5954 -1703 5997 -1693
rect 6012 -1679 6014 -1675
rect 6136 -1665 6196 -1651
tri 6250 -1656 6263 -1643 ne
rect 6263 -1649 6272 -1643
tri 6272 -1649 6278 -1643 sw
rect 6136 -1675 6181 -1665
rect 6012 -1703 6086 -1679
rect 5954 -1707 6086 -1703
tri 6086 -1707 6114 -1679 sw
rect 6136 -1689 6138 -1675
tri 6136 -1691 6138 -1689 ne
rect 6150 -1693 6181 -1675
rect 6150 -1703 6196 -1693
rect 6263 -1664 6278 -1649
tri 5888 -1728 5900 -1716 ne
rect 5900 -1721 5910 -1716
tri 5910 -1721 5915 -1716 sw
rect 5799 -2067 5814 -1839
rect 5900 -1877 5915 -1721
rect 5954 -1763 5982 -1707
tri 6074 -1725 6092 -1707 ne
rect 6092 -1727 6114 -1707
tri 6114 -1727 6134 -1707 sw
tri 6150 -1721 6168 -1703 ne
rect 5973 -1797 5982 -1763
rect 6016 -1736 6058 -1735
rect 6016 -1770 6021 -1736
rect 6051 -1770 6058 -1736
rect 6016 -1779 6058 -1770
rect 6092 -1736 6134 -1727
rect 6092 -1770 6099 -1736
rect 6129 -1770 6134 -1736
rect 6092 -1775 6134 -1770
rect 6168 -1763 6196 -1703
tri 6241 -1716 6263 -1694 se
rect 6263 -1701 6278 -1693
tri 6263 -1716 6278 -1701 nw
tri 6235 -1722 6241 -1716 se
rect 6241 -1722 6250 -1716
rect 5954 -1807 5982 -1797
tri 5982 -1807 6006 -1783 sw
rect 5954 -1839 5996 -1807
tri 6013 -1815 6014 -1814 sw
rect 6013 -1839 6014 -1815
tri 6016 -1816 6053 -1779 ne
rect 6053 -1807 6058 -1779
tri 6058 -1807 6084 -1781 sw
rect 6168 -1797 6177 -1763
rect 6168 -1807 6196 -1797
rect 6053 -1816 6137 -1807
tri 6053 -1835 6072 -1816 ne
rect 6072 -1835 6137 -1816
rect 5954 -1861 6014 -1839
rect 6136 -1839 6137 -1835
rect 6154 -1839 6196 -1807
rect 6136 -1861 6196 -1839
rect 6042 -1877 6059 -1863
rect 6091 -1877 6108 -1863
tri 5879 -1913 5901 -1891 se
rect 5901 -1898 5916 -1877
tri 5901 -1913 5916 -1898 nw
rect 6235 -1898 6250 -1722
tri 6250 -1729 6263 -1716 nw
rect 6336 -1797 6351 -1569
tri 5873 -1919 5879 -1913 se
rect 5879 -1919 5888 -1913
rect 5873 -1935 5888 -1919
tri 5888 -1926 5901 -1913 nw
rect 6042 -1921 6059 -1907
rect 6091 -1921 6108 -1907
tri 6235 -1913 6250 -1898 ne
tri 6250 -1913 6272 -1891 sw
rect 5873 -1971 5888 -1963
rect 5954 -1935 6014 -1921
rect 5969 -1945 6014 -1935
rect 5969 -1963 5997 -1945
tri 5873 -1986 5888 -1971 ne
tri 5888 -1986 5910 -1964 sw
rect 5954 -1973 5997 -1963
rect 6012 -1949 6014 -1945
rect 6136 -1935 6196 -1921
tri 6250 -1926 6263 -1913 ne
rect 6263 -1919 6272 -1913
tri 6272 -1919 6278 -1913 sw
rect 6136 -1945 6181 -1935
rect 6012 -1973 6086 -1949
rect 5954 -1977 6086 -1973
tri 6086 -1977 6114 -1949 sw
rect 6136 -1959 6138 -1945
tri 6136 -1961 6138 -1959 ne
rect 6150 -1963 6181 -1945
rect 6150 -1973 6196 -1963
rect 6263 -1934 6278 -1919
tri 5888 -1998 5900 -1986 ne
rect 5900 -1991 5910 -1986
tri 5910 -1991 5915 -1986 sw
rect 5799 -2147 5814 -2109
rect 5900 -2147 5915 -1991
rect 5954 -2033 5982 -1977
tri 6074 -1995 6092 -1977 ne
rect 6092 -1997 6114 -1977
tri 6114 -1997 6134 -1977 sw
tri 6150 -1991 6168 -1973 ne
rect 5973 -2067 5982 -2033
rect 6016 -2006 6058 -2005
rect 6016 -2040 6021 -2006
rect 6051 -2040 6058 -2006
rect 6016 -2049 6058 -2040
rect 6092 -2006 6134 -1997
rect 6092 -2040 6099 -2006
rect 6129 -2040 6134 -2006
rect 6092 -2045 6134 -2040
rect 6168 -2033 6196 -1973
tri 6241 -1986 6263 -1964 se
rect 6263 -1971 6278 -1963
tri 6263 -1986 6278 -1971 nw
tri 6235 -1992 6241 -1986 se
rect 6241 -1992 6250 -1986
rect 5954 -2077 5982 -2067
tri 5982 -2077 6006 -2053 sw
rect 5954 -2109 5996 -2077
tri 6013 -2085 6014 -2084 sw
rect 6013 -2109 6014 -2085
tri 6016 -2086 6053 -2049 ne
rect 6053 -2077 6058 -2049
tri 6058 -2077 6084 -2051 sw
rect 6168 -2067 6177 -2033
rect 6168 -2077 6196 -2067
rect 6053 -2086 6137 -2077
tri 6053 -2105 6072 -2086 ne
rect 6072 -2105 6137 -2086
rect 5954 -2131 6014 -2109
rect 6136 -2109 6137 -2105
rect 6154 -2109 6196 -2077
rect 6136 -2131 6196 -2109
rect 6042 -2147 6059 -2133
rect 6091 -2147 6108 -2133
rect 6235 -2147 6250 -1992
tri 6250 -1999 6263 -1986 nw
rect 6336 -2067 6351 -1839
rect 6336 -2147 6351 -2109
rect 6379 1984 6394 2174
tri 6459 2138 6481 2160 se
rect 6481 2153 6496 2174
tri 6481 2138 6496 2153 nw
rect 6815 2153 6830 2174
tri 6453 2132 6459 2138 se
rect 6459 2132 6468 2138
rect 6453 2116 6468 2132
tri 6468 2125 6481 2138 nw
rect 6622 2130 6639 2144
rect 6671 2130 6688 2144
tri 6815 2138 6830 2153 ne
tri 6830 2138 6852 2160 sw
rect 6453 2080 6468 2088
rect 6534 2116 6594 2130
rect 6549 2106 6594 2116
rect 6549 2088 6577 2106
tri 6453 2065 6468 2080 ne
tri 6468 2065 6490 2087 sw
rect 6534 2078 6577 2088
rect 6592 2102 6594 2106
rect 6716 2116 6776 2130
tri 6830 2125 6843 2138 ne
rect 6843 2132 6852 2138
tri 6852 2132 6858 2138 sw
rect 6716 2106 6761 2116
rect 6592 2078 6666 2102
rect 6534 2074 6666 2078
tri 6666 2074 6694 2102 sw
rect 6716 2092 6718 2106
tri 6716 2090 6718 2092 ne
rect 6730 2088 6761 2106
rect 6730 2078 6776 2088
rect 6843 2117 6858 2132
tri 6468 2053 6480 2065 ne
rect 6480 2060 6490 2065
tri 6490 2060 6495 2065 sw
rect 6379 1714 6394 1942
rect 6480 1904 6495 2060
rect 6534 2018 6562 2074
tri 6654 2056 6672 2074 ne
rect 6672 2054 6694 2074
tri 6694 2054 6714 2074 sw
tri 6730 2060 6748 2078 ne
rect 6553 1984 6562 2018
rect 6596 2045 6638 2046
rect 6596 2011 6601 2045
rect 6631 2011 6638 2045
rect 6596 2002 6638 2011
rect 6672 2045 6714 2054
rect 6672 2011 6679 2045
rect 6709 2011 6714 2045
rect 6672 2006 6714 2011
rect 6748 2018 6776 2078
tri 6821 2065 6843 2087 se
rect 6843 2080 6858 2088
tri 6843 2065 6858 2080 nw
tri 6815 2059 6821 2065 se
rect 6821 2059 6830 2065
rect 6534 1974 6562 1984
tri 6562 1974 6586 1998 sw
rect 6534 1942 6576 1974
tri 6593 1966 6594 1967 sw
rect 6593 1942 6594 1966
tri 6596 1965 6633 2002 ne
rect 6633 1974 6638 2002
tri 6638 1974 6664 2000 sw
rect 6748 1984 6757 2018
rect 6748 1974 6776 1984
rect 6633 1965 6717 1974
tri 6633 1946 6652 1965 ne
rect 6652 1946 6717 1965
rect 6534 1920 6594 1942
rect 6716 1942 6717 1946
rect 6734 1942 6776 1974
rect 6716 1920 6776 1942
rect 6622 1904 6639 1918
rect 6671 1904 6688 1918
tri 6459 1868 6481 1890 se
rect 6481 1883 6496 1904
tri 6481 1868 6496 1883 nw
rect 6815 1883 6830 2059
tri 6830 2052 6843 2065 nw
rect 6916 1984 6931 2174
tri 6453 1862 6459 1868 se
rect 6459 1862 6468 1868
rect 6453 1846 6468 1862
tri 6468 1855 6481 1868 nw
rect 6622 1860 6639 1874
rect 6671 1860 6688 1874
tri 6815 1868 6830 1883 ne
tri 6830 1868 6852 1890 sw
rect 6453 1810 6468 1818
rect 6534 1846 6594 1860
rect 6549 1836 6594 1846
rect 6549 1818 6577 1836
tri 6453 1795 6468 1810 ne
tri 6468 1795 6490 1817 sw
rect 6534 1808 6577 1818
rect 6592 1832 6594 1836
rect 6716 1846 6776 1860
tri 6830 1855 6843 1868 ne
rect 6843 1862 6852 1868
tri 6852 1862 6858 1868 sw
rect 6716 1836 6761 1846
rect 6592 1808 6666 1832
rect 6534 1804 6666 1808
tri 6666 1804 6694 1832 sw
rect 6716 1822 6718 1836
tri 6716 1820 6718 1822 ne
rect 6730 1818 6761 1836
rect 6730 1808 6776 1818
rect 6843 1847 6858 1862
tri 6468 1783 6480 1795 ne
rect 6480 1790 6490 1795
tri 6490 1790 6495 1795 sw
rect 6379 1444 6394 1672
rect 6480 1682 6495 1790
rect 6534 1748 6562 1804
tri 6654 1786 6672 1804 ne
rect 6672 1784 6694 1804
tri 6694 1784 6714 1804 sw
tri 6730 1790 6748 1808 ne
rect 6553 1714 6562 1748
rect 6596 1775 6638 1776
rect 6596 1741 6601 1775
rect 6631 1741 6638 1775
rect 6596 1732 6638 1741
rect 6672 1775 6714 1784
rect 6672 1741 6679 1775
rect 6709 1741 6714 1775
rect 6672 1736 6714 1741
rect 6748 1748 6776 1808
tri 6821 1795 6843 1817 se
rect 6843 1810 6858 1818
tri 6843 1795 6858 1810 nw
tri 6815 1789 6821 1795 se
rect 6821 1789 6830 1795
rect 6534 1704 6562 1714
tri 6562 1704 6586 1728 sw
rect 6480 1634 6496 1682
rect 6534 1672 6576 1704
tri 6593 1696 6594 1697 sw
rect 6593 1672 6594 1696
tri 6596 1695 6633 1732 ne
rect 6633 1704 6638 1732
tri 6638 1704 6664 1730 sw
rect 6748 1714 6757 1748
rect 6748 1704 6776 1714
rect 6633 1695 6717 1704
tri 6633 1676 6652 1695 ne
rect 6652 1676 6717 1695
rect 6534 1650 6594 1672
rect 6716 1672 6717 1676
rect 6734 1672 6776 1704
rect 6716 1650 6776 1672
rect 6622 1634 6639 1648
rect 6671 1634 6688 1648
tri 6459 1598 6481 1620 se
rect 6481 1613 6496 1634
tri 6481 1598 6496 1613 nw
rect 6815 1613 6830 1789
tri 6830 1782 6843 1795 nw
rect 6916 1714 6931 1942
tri 6453 1592 6459 1598 se
rect 6459 1592 6468 1598
rect 6453 1576 6468 1592
tri 6468 1585 6481 1598 nw
rect 6622 1590 6639 1604
rect 6671 1590 6688 1604
tri 6815 1598 6830 1613 ne
tri 6830 1598 6852 1620 sw
rect 6453 1540 6468 1548
rect 6534 1576 6594 1590
rect 6549 1566 6594 1576
rect 6549 1548 6577 1566
tri 6453 1525 6468 1540 ne
tri 6468 1525 6490 1547 sw
rect 6534 1538 6577 1548
rect 6592 1562 6594 1566
rect 6716 1576 6776 1590
tri 6830 1585 6843 1598 ne
rect 6843 1592 6852 1598
tri 6852 1592 6858 1598 sw
rect 6716 1566 6761 1576
rect 6592 1538 6666 1562
rect 6534 1534 6666 1538
tri 6666 1534 6694 1562 sw
rect 6716 1552 6718 1566
tri 6716 1550 6718 1552 ne
rect 6730 1548 6761 1566
rect 6730 1538 6776 1548
rect 6843 1577 6858 1592
tri 6468 1513 6480 1525 ne
rect 6480 1520 6490 1525
tri 6490 1520 6495 1525 sw
rect 6379 1174 6394 1402
rect 6480 1364 6495 1520
rect 6534 1478 6562 1534
tri 6654 1516 6672 1534 ne
rect 6672 1514 6694 1534
tri 6694 1514 6714 1534 sw
tri 6730 1520 6748 1538 ne
rect 6553 1444 6562 1478
rect 6596 1505 6638 1506
rect 6596 1471 6601 1505
rect 6631 1471 6638 1505
rect 6596 1462 6638 1471
rect 6672 1505 6714 1514
rect 6672 1471 6679 1505
rect 6709 1471 6714 1505
rect 6672 1466 6714 1471
rect 6748 1478 6776 1538
tri 6821 1525 6843 1547 se
rect 6843 1540 6858 1548
tri 6843 1525 6858 1540 nw
tri 6815 1519 6821 1525 se
rect 6821 1519 6830 1525
rect 6534 1434 6562 1444
tri 6562 1434 6586 1458 sw
rect 6534 1402 6576 1434
tri 6593 1426 6594 1427 sw
rect 6593 1402 6594 1426
tri 6596 1425 6633 1462 ne
rect 6633 1434 6638 1462
tri 6638 1434 6664 1460 sw
rect 6748 1444 6757 1478
rect 6748 1434 6776 1444
rect 6633 1425 6717 1434
tri 6633 1406 6652 1425 ne
rect 6652 1406 6717 1425
rect 6534 1380 6594 1402
rect 6716 1402 6717 1406
rect 6734 1402 6776 1434
rect 6716 1380 6776 1402
rect 6622 1364 6639 1378
rect 6671 1364 6688 1378
tri 6459 1328 6481 1350 se
rect 6481 1343 6496 1364
tri 6481 1328 6496 1343 nw
rect 6815 1343 6830 1519
tri 6830 1512 6843 1525 nw
rect 6916 1444 6931 1672
tri 6453 1322 6459 1328 se
rect 6459 1322 6468 1328
rect 6453 1306 6468 1322
tri 6468 1315 6481 1328 nw
rect 6622 1320 6639 1334
rect 6671 1320 6688 1334
tri 6815 1328 6830 1343 ne
tri 6830 1328 6852 1350 sw
rect 6453 1270 6468 1278
rect 6534 1306 6594 1320
rect 6549 1296 6594 1306
rect 6549 1278 6577 1296
tri 6453 1255 6468 1270 ne
tri 6468 1255 6490 1277 sw
rect 6534 1268 6577 1278
rect 6592 1292 6594 1296
rect 6716 1306 6776 1320
tri 6830 1315 6843 1328 ne
rect 6843 1322 6852 1328
tri 6852 1322 6858 1328 sw
rect 6716 1296 6761 1306
rect 6592 1268 6666 1292
rect 6534 1264 6666 1268
tri 6666 1264 6694 1292 sw
rect 6716 1282 6718 1296
tri 6716 1280 6718 1282 ne
rect 6730 1278 6761 1296
rect 6730 1268 6776 1278
rect 6843 1307 6858 1322
tri 6468 1243 6480 1255 ne
rect 6480 1250 6490 1255
tri 6490 1250 6495 1255 sw
rect 6379 903 6394 1132
rect 6480 1141 6495 1250
rect 6534 1208 6562 1264
tri 6654 1246 6672 1264 ne
rect 6672 1244 6694 1264
tri 6694 1244 6714 1264 sw
tri 6730 1250 6748 1268 ne
rect 6553 1174 6562 1208
rect 6596 1235 6638 1236
rect 6596 1201 6601 1235
rect 6631 1201 6638 1235
rect 6596 1192 6638 1201
rect 6672 1235 6714 1244
rect 6672 1201 6679 1235
rect 6709 1201 6714 1235
rect 6672 1196 6714 1201
rect 6748 1208 6776 1268
tri 6821 1255 6843 1277 se
rect 6843 1270 6858 1278
tri 6843 1255 6858 1270 nw
tri 6815 1249 6821 1255 se
rect 6821 1249 6830 1255
rect 6534 1164 6562 1174
tri 6562 1164 6586 1188 sw
rect 6480 1094 6496 1141
rect 6534 1132 6576 1164
tri 6593 1156 6594 1157 sw
rect 6593 1132 6594 1156
tri 6596 1155 6633 1192 ne
rect 6633 1164 6638 1192
tri 6638 1164 6664 1190 sw
rect 6748 1174 6757 1208
rect 6748 1164 6776 1174
rect 6633 1155 6717 1164
tri 6633 1136 6652 1155 ne
rect 6652 1136 6717 1155
rect 6534 1110 6594 1132
rect 6716 1132 6717 1136
rect 6734 1132 6776 1164
rect 6716 1110 6776 1132
rect 6622 1094 6639 1108
rect 6671 1094 6688 1108
tri 6459 1057 6481 1079 se
rect 6481 1072 6496 1094
tri 6481 1057 6496 1072 nw
rect 6815 1072 6830 1249
tri 6830 1242 6843 1255 nw
rect 6916 1174 6931 1402
tri 6453 1051 6459 1057 se
rect 6459 1051 6468 1057
rect 6453 1035 6468 1051
tri 6468 1044 6481 1057 nw
rect 6622 1049 6639 1063
rect 6671 1049 6688 1063
tri 6815 1057 6830 1072 ne
tri 6830 1057 6852 1079 sw
rect 6453 999 6468 1007
rect 6534 1035 6594 1049
rect 6549 1025 6594 1035
rect 6549 1007 6577 1025
tri 6453 984 6468 999 ne
tri 6468 984 6490 1006 sw
rect 6534 997 6577 1007
rect 6592 1021 6594 1025
rect 6716 1035 6776 1049
tri 6830 1044 6843 1057 ne
rect 6843 1051 6852 1057
tri 6852 1051 6858 1057 sw
rect 6716 1025 6761 1035
rect 6592 997 6666 1021
rect 6534 993 6666 997
tri 6666 993 6694 1021 sw
rect 6716 1011 6718 1025
tri 6716 1009 6718 1011 ne
rect 6730 1007 6761 1025
rect 6730 997 6776 1007
rect 6843 1036 6858 1051
tri 6468 972 6480 984 ne
rect 6480 979 6490 984
tri 6490 979 6495 984 sw
rect 6379 633 6394 861
rect 6480 823 6495 979
rect 6534 937 6562 993
tri 6654 975 6672 993 ne
rect 6672 973 6694 993
tri 6694 973 6714 993 sw
tri 6730 979 6748 997 ne
rect 6553 903 6562 937
rect 6596 964 6638 965
rect 6596 930 6601 964
rect 6631 930 6638 964
rect 6596 921 6638 930
rect 6672 964 6714 973
rect 6672 930 6679 964
rect 6709 930 6714 964
rect 6672 925 6714 930
rect 6748 937 6776 997
tri 6821 984 6843 1006 se
rect 6843 999 6858 1007
tri 6843 984 6858 999 nw
tri 6815 978 6821 984 se
rect 6821 978 6830 984
rect 6534 893 6562 903
tri 6562 893 6586 917 sw
rect 6534 861 6576 893
tri 6593 885 6594 886 sw
rect 6593 861 6594 885
tri 6596 884 6633 921 ne
rect 6633 893 6638 921
tri 6638 893 6664 919 sw
rect 6748 903 6757 937
rect 6748 893 6776 903
rect 6633 884 6717 893
tri 6633 865 6652 884 ne
rect 6652 865 6717 884
rect 6534 839 6594 861
rect 6716 861 6717 865
rect 6734 861 6776 893
rect 6716 839 6776 861
rect 6622 823 6639 837
rect 6671 823 6688 837
tri 6459 787 6481 809 se
rect 6481 802 6496 823
tri 6481 787 6496 802 nw
rect 6815 802 6830 978
tri 6830 971 6843 984 nw
rect 6916 903 6931 1132
tri 6453 781 6459 787 se
rect 6459 781 6468 787
rect 6453 765 6468 781
tri 6468 774 6481 787 nw
rect 6622 779 6639 793
rect 6671 779 6688 793
tri 6815 787 6830 802 ne
tri 6830 787 6852 809 sw
rect 6453 729 6468 737
rect 6534 765 6594 779
rect 6549 755 6594 765
rect 6549 737 6577 755
tri 6453 714 6468 729 ne
tri 6468 714 6490 736 sw
rect 6534 727 6577 737
rect 6592 751 6594 755
rect 6716 765 6776 779
tri 6830 774 6843 787 ne
rect 6843 781 6852 787
tri 6852 781 6858 787 sw
rect 6716 755 6761 765
rect 6592 727 6666 751
rect 6534 723 6666 727
tri 6666 723 6694 751 sw
rect 6716 741 6718 755
tri 6716 739 6718 741 ne
rect 6730 737 6761 755
rect 6730 727 6776 737
rect 6843 766 6858 781
tri 6468 702 6480 714 ne
rect 6480 709 6490 714
tri 6490 709 6495 714 sw
rect 6379 363 6394 591
rect 6480 601 6495 709
rect 6534 667 6562 723
tri 6654 705 6672 723 ne
rect 6672 703 6694 723
tri 6694 703 6714 723 sw
tri 6730 709 6748 727 ne
rect 6553 633 6562 667
rect 6596 694 6638 695
rect 6596 660 6601 694
rect 6631 660 6638 694
rect 6596 651 6638 660
rect 6672 694 6714 703
rect 6672 660 6679 694
rect 6709 660 6714 694
rect 6672 655 6714 660
rect 6748 667 6776 727
tri 6821 714 6843 736 se
rect 6843 729 6858 737
tri 6843 714 6858 729 nw
tri 6815 708 6821 714 se
rect 6821 708 6830 714
rect 6534 623 6562 633
tri 6562 623 6586 647 sw
rect 6480 553 6496 601
rect 6534 591 6576 623
tri 6593 615 6594 616 sw
rect 6593 591 6594 615
tri 6596 614 6633 651 ne
rect 6633 623 6638 651
tri 6638 623 6664 649 sw
rect 6748 633 6757 667
rect 6748 623 6776 633
rect 6633 614 6717 623
tri 6633 595 6652 614 ne
rect 6652 595 6717 614
rect 6534 569 6594 591
rect 6716 591 6717 595
rect 6734 591 6776 623
rect 6716 569 6776 591
rect 6622 553 6639 567
rect 6671 553 6688 567
tri 6459 517 6481 539 se
rect 6481 532 6496 553
tri 6481 517 6496 532 nw
rect 6815 532 6830 708
tri 6830 701 6843 714 nw
rect 6916 633 6931 861
tri 6453 511 6459 517 se
rect 6459 511 6468 517
rect 6453 495 6468 511
tri 6468 504 6481 517 nw
rect 6622 509 6639 523
rect 6671 509 6688 523
tri 6815 517 6830 532 ne
tri 6830 517 6852 539 sw
rect 6453 459 6468 467
rect 6534 495 6594 509
rect 6549 485 6594 495
rect 6549 467 6577 485
tri 6453 444 6468 459 ne
tri 6468 444 6490 466 sw
rect 6534 457 6577 467
rect 6592 481 6594 485
rect 6716 495 6776 509
tri 6830 504 6843 517 ne
rect 6843 511 6852 517
tri 6852 511 6858 517 sw
rect 6716 485 6761 495
rect 6592 457 6666 481
rect 6534 453 6666 457
tri 6666 453 6694 481 sw
rect 6716 471 6718 485
tri 6716 469 6718 471 ne
rect 6730 467 6761 485
rect 6730 457 6776 467
rect 6843 496 6858 511
tri 6468 432 6480 444 ne
rect 6480 439 6490 444
tri 6490 439 6495 444 sw
rect 6379 93 6394 321
rect 6480 283 6495 439
rect 6534 397 6562 453
tri 6654 435 6672 453 ne
rect 6672 433 6694 453
tri 6694 433 6714 453 sw
tri 6730 439 6748 457 ne
rect 6553 363 6562 397
rect 6596 424 6638 425
rect 6596 390 6601 424
rect 6631 390 6638 424
rect 6596 381 6638 390
rect 6672 424 6714 433
rect 6672 390 6679 424
rect 6709 390 6714 424
rect 6672 385 6714 390
rect 6748 397 6776 457
tri 6821 444 6843 466 se
rect 6843 459 6858 467
tri 6843 444 6858 459 nw
tri 6815 438 6821 444 se
rect 6821 438 6830 444
rect 6534 353 6562 363
tri 6562 353 6586 377 sw
rect 6534 321 6576 353
tri 6593 345 6594 346 sw
rect 6593 321 6594 345
tri 6596 344 6633 381 ne
rect 6633 353 6638 381
tri 6638 353 6664 379 sw
rect 6748 363 6757 397
rect 6748 353 6776 363
rect 6633 344 6717 353
tri 6633 325 6652 344 ne
rect 6652 325 6717 344
rect 6534 299 6594 321
rect 6716 321 6717 325
rect 6734 321 6776 353
rect 6716 299 6776 321
rect 6622 283 6639 297
rect 6671 283 6688 297
tri 6459 247 6481 269 se
rect 6481 262 6496 283
tri 6481 247 6496 262 nw
rect 6815 262 6830 438
tri 6830 431 6843 444 nw
rect 6916 363 6931 591
tri 6453 241 6459 247 se
rect 6459 241 6468 247
rect 6453 225 6468 241
tri 6468 234 6481 247 nw
rect 6622 239 6639 253
rect 6671 239 6688 253
tri 6815 247 6830 262 ne
tri 6830 247 6852 269 sw
rect 6453 189 6468 197
rect 6534 225 6594 239
rect 6549 215 6594 225
rect 6549 197 6577 215
tri 6453 174 6468 189 ne
tri 6468 174 6490 196 sw
rect 6534 187 6577 197
rect 6592 211 6594 215
rect 6716 225 6776 239
tri 6830 234 6843 247 ne
rect 6843 241 6852 247
tri 6852 241 6858 247 sw
rect 6716 215 6761 225
rect 6592 187 6666 211
rect 6534 183 6666 187
tri 6666 183 6694 211 sw
rect 6716 201 6718 215
tri 6716 199 6718 201 ne
rect 6730 197 6761 215
rect 6730 187 6776 197
rect 6843 226 6858 241
tri 6468 162 6480 174 ne
rect 6480 169 6490 174
tri 6490 169 6495 174 sw
rect 6379 -177 6394 51
rect 6480 61 6495 169
rect 6534 127 6562 183
tri 6654 165 6672 183 ne
rect 6672 163 6694 183
tri 6694 163 6714 183 sw
tri 6730 169 6748 187 ne
rect 6553 93 6562 127
rect 6596 154 6638 155
rect 6596 120 6601 154
rect 6631 120 6638 154
rect 6596 111 6638 120
rect 6672 154 6714 163
rect 6672 120 6679 154
rect 6709 120 6714 154
rect 6672 115 6714 120
rect 6748 127 6776 187
tri 6821 174 6843 196 se
rect 6843 189 6858 197
tri 6843 174 6858 189 nw
tri 6815 168 6821 174 se
rect 6821 168 6830 174
rect 6534 83 6562 93
tri 6562 83 6586 107 sw
rect 6480 13 6496 61
rect 6534 51 6576 83
tri 6593 75 6594 76 sw
rect 6593 51 6594 75
tri 6596 74 6633 111 ne
rect 6633 83 6638 111
tri 6638 83 6664 109 sw
rect 6748 93 6757 127
rect 6748 83 6776 93
rect 6633 74 6717 83
tri 6633 55 6652 74 ne
rect 6652 55 6717 74
rect 6534 29 6594 51
rect 6716 51 6717 55
rect 6734 51 6776 83
rect 6716 29 6776 51
rect 6622 13 6639 27
rect 6671 13 6688 27
tri 6459 -23 6481 -1 se
rect 6481 -8 6496 13
tri 6481 -23 6496 -8 nw
rect 6815 -8 6830 168
tri 6830 161 6843 174 nw
rect 6916 93 6931 321
tri 6453 -29 6459 -23 se
rect 6459 -29 6468 -23
rect 6453 -45 6468 -29
tri 6468 -36 6481 -23 nw
rect 6622 -31 6639 -17
rect 6671 -31 6688 -17
tri 6815 -23 6830 -8 ne
tri 6830 -23 6852 -1 sw
rect 6453 -81 6468 -73
rect 6534 -45 6594 -31
rect 6549 -55 6594 -45
rect 6549 -73 6577 -55
tri 6453 -96 6468 -81 ne
tri 6468 -96 6490 -74 sw
rect 6534 -83 6577 -73
rect 6592 -59 6594 -55
rect 6716 -45 6776 -31
tri 6830 -36 6843 -23 ne
rect 6843 -29 6852 -23
tri 6852 -29 6858 -23 sw
rect 6716 -55 6761 -45
rect 6592 -83 6666 -59
rect 6534 -87 6666 -83
tri 6666 -87 6694 -59 sw
rect 6716 -69 6718 -55
tri 6716 -71 6718 -69 ne
rect 6730 -73 6761 -55
rect 6730 -83 6776 -73
rect 6843 -44 6858 -29
tri 6468 -108 6480 -96 ne
rect 6480 -101 6490 -96
tri 6490 -101 6495 -96 sw
rect 6379 -447 6394 -219
rect 6480 -257 6495 -101
rect 6534 -143 6562 -87
tri 6654 -105 6672 -87 ne
rect 6672 -107 6694 -87
tri 6694 -107 6714 -87 sw
tri 6730 -101 6748 -83 ne
rect 6553 -177 6562 -143
rect 6596 -116 6638 -115
rect 6596 -150 6601 -116
rect 6631 -150 6638 -116
rect 6596 -159 6638 -150
rect 6672 -116 6714 -107
rect 6672 -150 6679 -116
rect 6709 -150 6714 -116
rect 6672 -155 6714 -150
rect 6748 -143 6776 -83
tri 6821 -96 6843 -74 se
rect 6843 -81 6858 -73
tri 6843 -96 6858 -81 nw
tri 6815 -102 6821 -96 se
rect 6821 -102 6830 -96
rect 6534 -187 6562 -177
tri 6562 -187 6586 -163 sw
rect 6534 -219 6576 -187
tri 6593 -195 6594 -194 sw
rect 6593 -219 6594 -195
tri 6596 -196 6633 -159 ne
rect 6633 -187 6638 -159
tri 6638 -187 6664 -161 sw
rect 6748 -177 6757 -143
rect 6748 -187 6776 -177
rect 6633 -196 6717 -187
tri 6633 -215 6652 -196 ne
rect 6652 -215 6717 -196
rect 6534 -241 6594 -219
rect 6716 -219 6717 -215
rect 6734 -219 6776 -187
rect 6716 -241 6776 -219
rect 6622 -257 6639 -243
rect 6671 -257 6688 -243
tri 6459 -293 6481 -271 se
rect 6481 -278 6496 -257
tri 6481 -293 6496 -278 nw
rect 6815 -278 6830 -102
tri 6830 -109 6843 -96 nw
rect 6916 -177 6931 51
tri 6453 -299 6459 -293 se
rect 6459 -299 6468 -293
rect 6453 -315 6468 -299
tri 6468 -306 6481 -293 nw
rect 6622 -301 6639 -287
rect 6671 -301 6688 -287
tri 6815 -293 6830 -278 ne
tri 6830 -293 6852 -271 sw
rect 6453 -351 6468 -343
rect 6534 -315 6594 -301
rect 6549 -325 6594 -315
rect 6549 -343 6577 -325
tri 6453 -366 6468 -351 ne
tri 6468 -366 6490 -344 sw
rect 6534 -353 6577 -343
rect 6592 -329 6594 -325
rect 6716 -315 6776 -301
tri 6830 -306 6843 -293 ne
rect 6843 -299 6852 -293
tri 6852 -299 6858 -293 sw
rect 6716 -325 6761 -315
rect 6592 -353 6666 -329
rect 6534 -357 6666 -353
tri 6666 -357 6694 -329 sw
rect 6716 -339 6718 -325
tri 6716 -341 6718 -339 ne
rect 6730 -343 6761 -325
rect 6730 -353 6776 -343
rect 6843 -314 6858 -299
tri 6468 -378 6480 -366 ne
rect 6480 -371 6490 -366
tri 6490 -371 6495 -366 sw
rect 6379 -717 6394 -489
rect 6480 -479 6495 -371
rect 6534 -413 6562 -357
tri 6654 -375 6672 -357 ne
rect 6672 -377 6694 -357
tri 6694 -377 6714 -357 sw
tri 6730 -371 6748 -353 ne
rect 6553 -447 6562 -413
rect 6596 -386 6638 -385
rect 6596 -420 6601 -386
rect 6631 -420 6638 -386
rect 6596 -429 6638 -420
rect 6672 -386 6714 -377
rect 6672 -420 6679 -386
rect 6709 -420 6714 -386
rect 6672 -425 6714 -420
rect 6748 -413 6776 -353
tri 6821 -366 6843 -344 se
rect 6843 -351 6858 -343
tri 6843 -366 6858 -351 nw
tri 6815 -372 6821 -366 se
rect 6821 -372 6830 -366
rect 6534 -457 6562 -447
tri 6562 -457 6586 -433 sw
rect 6480 -527 6496 -479
rect 6534 -489 6576 -457
tri 6593 -465 6594 -464 sw
rect 6593 -489 6594 -465
tri 6596 -466 6633 -429 ne
rect 6633 -457 6638 -429
tri 6638 -457 6664 -431 sw
rect 6748 -447 6757 -413
rect 6748 -457 6776 -447
rect 6633 -466 6717 -457
tri 6633 -485 6652 -466 ne
rect 6652 -485 6717 -466
rect 6534 -511 6594 -489
rect 6716 -489 6717 -485
rect 6734 -489 6776 -457
rect 6716 -511 6776 -489
rect 6622 -527 6639 -513
rect 6671 -527 6688 -513
tri 6459 -563 6481 -541 se
rect 6481 -548 6496 -527
tri 6481 -563 6496 -548 nw
rect 6815 -548 6830 -372
tri 6830 -379 6843 -366 nw
rect 6916 -447 6931 -219
tri 6453 -569 6459 -563 se
rect 6459 -569 6468 -563
rect 6453 -585 6468 -569
tri 6468 -576 6481 -563 nw
rect 6622 -571 6639 -557
rect 6671 -571 6688 -557
tri 6815 -563 6830 -548 ne
tri 6830 -563 6852 -541 sw
rect 6453 -621 6468 -613
rect 6534 -585 6594 -571
rect 6549 -595 6594 -585
rect 6549 -613 6577 -595
tri 6453 -636 6468 -621 ne
tri 6468 -636 6490 -614 sw
rect 6534 -623 6577 -613
rect 6592 -599 6594 -595
rect 6716 -585 6776 -571
tri 6830 -576 6843 -563 ne
rect 6843 -569 6852 -563
tri 6852 -569 6858 -563 sw
rect 6716 -595 6761 -585
rect 6592 -623 6666 -599
rect 6534 -627 6666 -623
tri 6666 -627 6694 -599 sw
rect 6716 -609 6718 -595
tri 6716 -611 6718 -609 ne
rect 6730 -613 6761 -595
rect 6730 -623 6776 -613
rect 6843 -584 6858 -569
tri 6468 -648 6480 -636 ne
rect 6480 -641 6490 -636
tri 6490 -641 6495 -636 sw
rect 6379 -987 6394 -759
rect 6480 -797 6495 -641
rect 6534 -683 6562 -627
tri 6654 -645 6672 -627 ne
rect 6672 -647 6694 -627
tri 6694 -647 6714 -627 sw
tri 6730 -641 6748 -623 ne
rect 6553 -717 6562 -683
rect 6596 -656 6638 -655
rect 6596 -690 6601 -656
rect 6631 -690 6638 -656
rect 6596 -699 6638 -690
rect 6672 -656 6714 -647
rect 6672 -690 6679 -656
rect 6709 -690 6714 -656
rect 6672 -695 6714 -690
rect 6748 -683 6776 -623
tri 6821 -636 6843 -614 se
rect 6843 -621 6858 -613
tri 6843 -636 6858 -621 nw
tri 6815 -642 6821 -636 se
rect 6821 -642 6830 -636
rect 6534 -727 6562 -717
tri 6562 -727 6586 -703 sw
rect 6534 -759 6576 -727
tri 6593 -735 6594 -734 sw
rect 6593 -759 6594 -735
tri 6596 -736 6633 -699 ne
rect 6633 -727 6638 -699
tri 6638 -727 6664 -701 sw
rect 6748 -717 6757 -683
rect 6748 -727 6776 -717
rect 6633 -736 6717 -727
tri 6633 -755 6652 -736 ne
rect 6652 -755 6717 -736
rect 6534 -781 6594 -759
rect 6716 -759 6717 -755
rect 6734 -759 6776 -727
rect 6716 -781 6776 -759
rect 6622 -797 6639 -783
rect 6671 -797 6688 -783
tri 6459 -833 6481 -811 se
rect 6481 -818 6496 -797
tri 6481 -833 6496 -818 nw
rect 6815 -818 6830 -642
tri 6830 -649 6843 -636 nw
rect 6916 -717 6931 -489
tri 6453 -839 6459 -833 se
rect 6459 -839 6468 -833
rect 6453 -855 6468 -839
tri 6468 -846 6481 -833 nw
rect 6622 -841 6639 -827
rect 6671 -841 6688 -827
tri 6815 -833 6830 -818 ne
tri 6830 -833 6852 -811 sw
rect 6453 -891 6468 -883
rect 6534 -855 6594 -841
rect 6549 -865 6594 -855
rect 6549 -883 6577 -865
tri 6453 -906 6468 -891 ne
tri 6468 -906 6490 -884 sw
rect 6534 -893 6577 -883
rect 6592 -869 6594 -865
rect 6716 -855 6776 -841
tri 6830 -846 6843 -833 ne
rect 6843 -839 6852 -833
tri 6852 -839 6858 -833 sw
rect 6716 -865 6761 -855
rect 6592 -893 6666 -869
rect 6534 -897 6666 -893
tri 6666 -897 6694 -869 sw
rect 6716 -879 6718 -865
tri 6716 -881 6718 -879 ne
rect 6730 -883 6761 -865
rect 6730 -893 6776 -883
rect 6843 -854 6858 -839
tri 6468 -918 6480 -906 ne
rect 6480 -911 6490 -906
tri 6490 -911 6495 -906 sw
rect 6379 -1257 6394 -1029
rect 6480 -1019 6495 -911
rect 6534 -953 6562 -897
tri 6654 -915 6672 -897 ne
rect 6672 -917 6694 -897
tri 6694 -917 6714 -897 sw
tri 6730 -911 6748 -893 ne
rect 6553 -987 6562 -953
rect 6596 -926 6638 -925
rect 6596 -960 6601 -926
rect 6631 -960 6638 -926
rect 6596 -969 6638 -960
rect 6672 -926 6714 -917
rect 6672 -960 6679 -926
rect 6709 -960 6714 -926
rect 6672 -965 6714 -960
rect 6748 -953 6776 -893
tri 6821 -906 6843 -884 se
rect 6843 -891 6858 -883
tri 6843 -906 6858 -891 nw
tri 6815 -912 6821 -906 se
rect 6821 -912 6830 -906
rect 6534 -997 6562 -987
tri 6562 -997 6586 -973 sw
rect 6480 -1067 6496 -1019
rect 6534 -1029 6576 -997
tri 6593 -1005 6594 -1004 sw
rect 6593 -1029 6594 -1005
tri 6596 -1006 6633 -969 ne
rect 6633 -997 6638 -969
tri 6638 -997 6664 -971 sw
rect 6748 -987 6757 -953
rect 6748 -997 6776 -987
rect 6633 -1006 6717 -997
tri 6633 -1025 6652 -1006 ne
rect 6652 -1025 6717 -1006
rect 6534 -1051 6594 -1029
rect 6716 -1029 6717 -1025
rect 6734 -1029 6776 -997
rect 6716 -1051 6776 -1029
rect 6622 -1067 6639 -1053
rect 6671 -1067 6688 -1053
tri 6459 -1103 6481 -1081 se
rect 6481 -1088 6496 -1067
tri 6481 -1103 6496 -1088 nw
rect 6815 -1088 6830 -912
tri 6830 -919 6843 -906 nw
rect 6916 -987 6931 -759
tri 6453 -1109 6459 -1103 se
rect 6459 -1109 6468 -1103
rect 6453 -1125 6468 -1109
tri 6468 -1116 6481 -1103 nw
rect 6622 -1111 6639 -1097
rect 6671 -1111 6688 -1097
tri 6815 -1103 6830 -1088 ne
tri 6830 -1103 6852 -1081 sw
rect 6453 -1161 6468 -1153
rect 6534 -1125 6594 -1111
rect 6549 -1135 6594 -1125
rect 6549 -1153 6577 -1135
tri 6453 -1176 6468 -1161 ne
tri 6468 -1176 6490 -1154 sw
rect 6534 -1163 6577 -1153
rect 6592 -1139 6594 -1135
rect 6716 -1125 6776 -1111
tri 6830 -1116 6843 -1103 ne
rect 6843 -1109 6852 -1103
tri 6852 -1109 6858 -1103 sw
rect 6716 -1135 6761 -1125
rect 6592 -1163 6666 -1139
rect 6534 -1167 6666 -1163
tri 6666 -1167 6694 -1139 sw
rect 6716 -1149 6718 -1135
tri 6716 -1151 6718 -1149 ne
rect 6730 -1153 6761 -1135
rect 6730 -1163 6776 -1153
rect 6843 -1124 6858 -1109
tri 6468 -1188 6480 -1176 ne
rect 6480 -1181 6490 -1176
tri 6490 -1181 6495 -1176 sw
rect 6379 -1527 6394 -1299
rect 6480 -1337 6495 -1181
rect 6534 -1223 6562 -1167
tri 6654 -1185 6672 -1167 ne
rect 6672 -1187 6694 -1167
tri 6694 -1187 6714 -1167 sw
tri 6730 -1181 6748 -1163 ne
rect 6553 -1257 6562 -1223
rect 6596 -1196 6638 -1195
rect 6596 -1230 6601 -1196
rect 6631 -1230 6638 -1196
rect 6596 -1239 6638 -1230
rect 6672 -1196 6714 -1187
rect 6672 -1230 6679 -1196
rect 6709 -1230 6714 -1196
rect 6672 -1235 6714 -1230
rect 6748 -1223 6776 -1163
tri 6821 -1176 6843 -1154 se
rect 6843 -1161 6858 -1153
tri 6843 -1176 6858 -1161 nw
tri 6815 -1182 6821 -1176 se
rect 6821 -1182 6830 -1176
rect 6534 -1267 6562 -1257
tri 6562 -1267 6586 -1243 sw
rect 6534 -1299 6576 -1267
tri 6593 -1275 6594 -1274 sw
rect 6593 -1299 6594 -1275
tri 6596 -1276 6633 -1239 ne
rect 6633 -1267 6638 -1239
tri 6638 -1267 6664 -1241 sw
rect 6748 -1257 6757 -1223
rect 6748 -1267 6776 -1257
rect 6633 -1276 6717 -1267
tri 6633 -1295 6652 -1276 ne
rect 6652 -1295 6717 -1276
rect 6534 -1321 6594 -1299
rect 6716 -1299 6717 -1295
rect 6734 -1299 6776 -1267
rect 6716 -1321 6776 -1299
rect 6622 -1337 6639 -1323
rect 6671 -1337 6688 -1323
tri 6459 -1373 6481 -1351 se
rect 6481 -1358 6496 -1337
tri 6481 -1373 6496 -1358 nw
rect 6815 -1358 6830 -1182
tri 6830 -1189 6843 -1176 nw
rect 6916 -1257 6931 -1029
tri 6453 -1379 6459 -1373 se
rect 6459 -1379 6468 -1373
rect 6453 -1395 6468 -1379
tri 6468 -1386 6481 -1373 nw
rect 6622 -1381 6639 -1367
rect 6671 -1381 6688 -1367
tri 6815 -1373 6830 -1358 ne
tri 6830 -1373 6852 -1351 sw
rect 6453 -1431 6468 -1423
rect 6534 -1395 6594 -1381
rect 6549 -1405 6594 -1395
rect 6549 -1423 6577 -1405
tri 6453 -1446 6468 -1431 ne
tri 6468 -1446 6490 -1424 sw
rect 6534 -1433 6577 -1423
rect 6592 -1409 6594 -1405
rect 6716 -1395 6776 -1381
tri 6830 -1386 6843 -1373 ne
rect 6843 -1379 6852 -1373
tri 6852 -1379 6858 -1373 sw
rect 6716 -1405 6761 -1395
rect 6592 -1433 6666 -1409
rect 6534 -1437 6666 -1433
tri 6666 -1437 6694 -1409 sw
rect 6716 -1419 6718 -1405
tri 6716 -1421 6718 -1419 ne
rect 6730 -1423 6761 -1405
rect 6730 -1433 6776 -1423
rect 6843 -1394 6858 -1379
tri 6468 -1458 6480 -1446 ne
rect 6480 -1451 6490 -1446
tri 6490 -1451 6495 -1446 sw
rect 6379 -1797 6394 -1569
rect 6480 -1559 6495 -1451
rect 6534 -1493 6562 -1437
tri 6654 -1455 6672 -1437 ne
rect 6672 -1457 6694 -1437
tri 6694 -1457 6714 -1437 sw
tri 6730 -1451 6748 -1433 ne
rect 6553 -1527 6562 -1493
rect 6596 -1466 6638 -1465
rect 6596 -1500 6601 -1466
rect 6631 -1500 6638 -1466
rect 6596 -1509 6638 -1500
rect 6672 -1466 6714 -1457
rect 6672 -1500 6679 -1466
rect 6709 -1500 6714 -1466
rect 6672 -1505 6714 -1500
rect 6748 -1493 6776 -1433
tri 6821 -1446 6843 -1424 se
rect 6843 -1431 6858 -1423
tri 6843 -1446 6858 -1431 nw
tri 6815 -1452 6821 -1446 se
rect 6821 -1452 6830 -1446
rect 6534 -1537 6562 -1527
tri 6562 -1537 6586 -1513 sw
rect 6480 -1607 6496 -1559
rect 6534 -1569 6576 -1537
tri 6593 -1545 6594 -1544 sw
rect 6593 -1569 6594 -1545
tri 6596 -1546 6633 -1509 ne
rect 6633 -1537 6638 -1509
tri 6638 -1537 6664 -1511 sw
rect 6748 -1527 6757 -1493
rect 6748 -1537 6776 -1527
rect 6633 -1546 6717 -1537
tri 6633 -1565 6652 -1546 ne
rect 6652 -1565 6717 -1546
rect 6534 -1591 6594 -1569
rect 6716 -1569 6717 -1565
rect 6734 -1569 6776 -1537
rect 6716 -1591 6776 -1569
rect 6622 -1607 6639 -1593
rect 6671 -1607 6688 -1593
tri 6459 -1643 6481 -1621 se
rect 6481 -1628 6496 -1607
tri 6481 -1643 6496 -1628 nw
rect 6815 -1628 6830 -1452
tri 6830 -1459 6843 -1446 nw
rect 6916 -1527 6931 -1299
tri 6453 -1649 6459 -1643 se
rect 6459 -1649 6468 -1643
rect 6453 -1665 6468 -1649
tri 6468 -1656 6481 -1643 nw
rect 6622 -1651 6639 -1637
rect 6671 -1651 6688 -1637
tri 6815 -1643 6830 -1628 ne
tri 6830 -1643 6852 -1621 sw
rect 6453 -1701 6468 -1693
rect 6534 -1665 6594 -1651
rect 6549 -1675 6594 -1665
rect 6549 -1693 6577 -1675
tri 6453 -1716 6468 -1701 ne
tri 6468 -1716 6490 -1694 sw
rect 6534 -1703 6577 -1693
rect 6592 -1679 6594 -1675
rect 6716 -1665 6776 -1651
tri 6830 -1656 6843 -1643 ne
rect 6843 -1649 6852 -1643
tri 6852 -1649 6858 -1643 sw
rect 6716 -1675 6761 -1665
rect 6592 -1703 6666 -1679
rect 6534 -1707 6666 -1703
tri 6666 -1707 6694 -1679 sw
rect 6716 -1689 6718 -1675
tri 6716 -1691 6718 -1689 ne
rect 6730 -1693 6761 -1675
rect 6730 -1703 6776 -1693
rect 6843 -1664 6858 -1649
tri 6468 -1728 6480 -1716 ne
rect 6480 -1721 6490 -1716
tri 6490 -1721 6495 -1716 sw
rect 6379 -2067 6394 -1839
rect 6480 -1877 6495 -1721
rect 6534 -1763 6562 -1707
tri 6654 -1725 6672 -1707 ne
rect 6672 -1727 6694 -1707
tri 6694 -1727 6714 -1707 sw
tri 6730 -1721 6748 -1703 ne
rect 6553 -1797 6562 -1763
rect 6596 -1736 6638 -1735
rect 6596 -1770 6601 -1736
rect 6631 -1770 6638 -1736
rect 6596 -1779 6638 -1770
rect 6672 -1736 6714 -1727
rect 6672 -1770 6679 -1736
rect 6709 -1770 6714 -1736
rect 6672 -1775 6714 -1770
rect 6748 -1763 6776 -1703
tri 6821 -1716 6843 -1694 se
rect 6843 -1701 6858 -1693
tri 6843 -1716 6858 -1701 nw
tri 6815 -1722 6821 -1716 se
rect 6821 -1722 6830 -1716
rect 6534 -1807 6562 -1797
tri 6562 -1807 6586 -1783 sw
rect 6534 -1839 6576 -1807
tri 6593 -1815 6594 -1814 sw
rect 6593 -1839 6594 -1815
tri 6596 -1816 6633 -1779 ne
rect 6633 -1807 6638 -1779
tri 6638 -1807 6664 -1781 sw
rect 6748 -1797 6757 -1763
rect 6748 -1807 6776 -1797
rect 6633 -1816 6717 -1807
tri 6633 -1835 6652 -1816 ne
rect 6652 -1835 6717 -1816
rect 6534 -1861 6594 -1839
rect 6716 -1839 6717 -1835
rect 6734 -1839 6776 -1807
rect 6716 -1861 6776 -1839
rect 6622 -1877 6639 -1863
rect 6671 -1877 6688 -1863
tri 6459 -1913 6481 -1891 se
rect 6481 -1898 6496 -1877
tri 6481 -1913 6496 -1898 nw
rect 6815 -1898 6830 -1722
tri 6830 -1729 6843 -1716 nw
rect 6916 -1797 6931 -1569
tri 6453 -1919 6459 -1913 se
rect 6459 -1919 6468 -1913
rect 6453 -1935 6468 -1919
tri 6468 -1926 6481 -1913 nw
rect 6622 -1921 6639 -1907
rect 6671 -1921 6688 -1907
tri 6815 -1913 6830 -1898 ne
tri 6830 -1913 6852 -1891 sw
rect 6453 -1971 6468 -1963
rect 6534 -1935 6594 -1921
rect 6549 -1945 6594 -1935
rect 6549 -1963 6577 -1945
tri 6453 -1986 6468 -1971 ne
tri 6468 -1986 6490 -1964 sw
rect 6534 -1973 6577 -1963
rect 6592 -1949 6594 -1945
rect 6716 -1935 6776 -1921
tri 6830 -1926 6843 -1913 ne
rect 6843 -1919 6852 -1913
tri 6852 -1919 6858 -1913 sw
rect 6716 -1945 6761 -1935
rect 6592 -1973 6666 -1949
rect 6534 -1977 6666 -1973
tri 6666 -1977 6694 -1949 sw
rect 6716 -1959 6718 -1945
tri 6716 -1961 6718 -1959 ne
rect 6730 -1963 6761 -1945
rect 6730 -1973 6776 -1963
rect 6843 -1934 6858 -1919
tri 6468 -1998 6480 -1986 ne
rect 6480 -1991 6490 -1986
tri 6490 -1991 6495 -1986 sw
rect 6379 -2147 6394 -2109
rect 6480 -2147 6495 -1991
rect 6534 -2033 6562 -1977
tri 6654 -1995 6672 -1977 ne
rect 6672 -1997 6694 -1977
tri 6694 -1997 6714 -1977 sw
tri 6730 -1991 6748 -1973 ne
rect 6553 -2067 6562 -2033
rect 6596 -2006 6638 -2005
rect 6596 -2040 6601 -2006
rect 6631 -2040 6638 -2006
rect 6596 -2049 6638 -2040
rect 6672 -2006 6714 -1997
rect 6672 -2040 6679 -2006
rect 6709 -2040 6714 -2006
rect 6672 -2045 6714 -2040
rect 6748 -2033 6776 -1973
tri 6821 -1986 6843 -1964 se
rect 6843 -1971 6858 -1963
tri 6843 -1986 6858 -1971 nw
tri 6815 -1992 6821 -1986 se
rect 6821 -1992 6830 -1986
rect 6534 -2077 6562 -2067
tri 6562 -2077 6586 -2053 sw
rect 6534 -2109 6576 -2077
tri 6593 -2085 6594 -2084 sw
rect 6593 -2109 6594 -2085
tri 6596 -2086 6633 -2049 ne
rect 6633 -2077 6638 -2049
tri 6638 -2077 6664 -2051 sw
rect 6748 -2067 6757 -2033
rect 6748 -2077 6776 -2067
rect 6633 -2086 6717 -2077
tri 6633 -2105 6652 -2086 ne
rect 6652 -2105 6717 -2086
rect 6534 -2131 6594 -2109
rect 6716 -2109 6717 -2105
rect 6734 -2109 6776 -2077
rect 6716 -2131 6776 -2109
rect 6622 -2147 6639 -2133
rect 6671 -2147 6688 -2133
rect 6815 -2147 6830 -1992
tri 6830 -1999 6843 -1986 nw
rect 6916 -2067 6931 -1839
rect 6916 -2147 6931 -2109
<< viali >>
rect 259 2130 291 2144
rect 42 2006 72 2040
rect 259 1904 291 1918
rect 478 2006 508 2040
rect 259 1860 291 1874
rect 42 1736 72 1770
rect 259 1634 291 1648
rect 478 1736 508 1770
rect 259 1590 291 1604
rect 42 1466 72 1500
rect 259 1364 291 1378
rect 478 1466 508 1500
rect 259 1320 291 1334
rect 42 1196 72 1230
rect 259 1094 291 1108
rect 478 1196 508 1230
rect 259 1050 291 1064
rect 42 926 72 960
rect 259 824 291 838
rect 478 926 508 960
rect 259 780 291 794
rect 42 656 72 690
rect 259 554 291 568
rect 478 656 508 690
rect 259 510 291 524
rect 42 386 72 420
rect 259 284 291 298
rect 478 386 508 420
rect 259 240 291 254
rect 42 116 72 150
rect 259 14 291 28
rect 478 116 508 150
rect 259 -30 291 -16
rect 42 -154 72 -120
rect 259 -256 291 -242
rect 478 -154 508 -120
rect 259 -300 291 -286
rect 42 -424 72 -390
rect 259 -526 291 -512
rect 478 -424 508 -390
rect 259 -570 291 -556
rect 42 -694 72 -660
rect 259 -796 291 -782
rect 478 -694 508 -660
rect 259 -840 291 -826
rect 42 -964 72 -930
rect 259 -1066 291 -1052
rect 478 -964 508 -930
rect 259 -1110 291 -1096
rect 42 -1234 72 -1200
rect 259 -1336 291 -1322
rect 478 -1234 508 -1200
rect 259 -1380 291 -1366
rect 42 -1504 72 -1470
rect 259 -1606 291 -1592
rect 478 -1504 508 -1470
rect 259 -1650 291 -1636
rect 42 -1774 72 -1740
rect 259 -1876 291 -1862
rect 478 -1774 508 -1740
rect 259 -1920 291 -1906
rect 42 -2044 72 -2010
rect 259 -2146 291 -2132
rect 478 -2044 508 -2010
rect 839 2130 871 2144
rect 622 2006 652 2040
rect 839 1904 871 1918
rect 1058 2006 1088 2040
rect 839 1860 871 1874
rect 622 1736 652 1770
rect 839 1634 871 1648
rect 1058 1736 1088 1770
rect 839 1590 871 1604
rect 622 1466 652 1500
rect 839 1364 871 1378
rect 1058 1466 1088 1500
rect 839 1320 871 1334
rect 622 1196 652 1230
rect 839 1094 871 1108
rect 1058 1196 1088 1230
rect 839 1050 871 1064
rect 622 926 652 960
rect 839 824 871 838
rect 1058 926 1088 960
rect 839 780 871 794
rect 622 656 652 690
rect 839 554 871 568
rect 1058 656 1088 690
rect 839 510 871 524
rect 622 386 652 420
rect 839 284 871 298
rect 1058 386 1088 420
rect 839 240 871 254
rect 622 116 652 150
rect 839 14 871 28
rect 1058 116 1088 150
rect 839 -30 871 -16
rect 622 -154 652 -120
rect 839 -256 871 -242
rect 1058 -154 1088 -120
rect 839 -300 871 -286
rect 622 -424 652 -390
rect 839 -526 871 -512
rect 1058 -424 1088 -390
rect 839 -570 871 -556
rect 622 -694 652 -660
rect 839 -796 871 -782
rect 1058 -694 1088 -660
rect 839 -840 871 -826
rect 622 -964 652 -930
rect 839 -1066 871 -1052
rect 1058 -964 1088 -930
rect 839 -1110 871 -1096
rect 622 -1234 652 -1200
rect 839 -1336 871 -1322
rect 1058 -1234 1088 -1200
rect 839 -1380 871 -1366
rect 622 -1504 652 -1470
rect 839 -1606 871 -1592
rect 1058 -1504 1088 -1470
rect 839 -1650 871 -1636
rect 622 -1774 652 -1740
rect 839 -1876 871 -1862
rect 1058 -1774 1088 -1740
rect 839 -1920 871 -1906
rect 622 -2044 652 -2010
rect 839 -2146 871 -2132
rect 1058 -2044 1088 -2010
rect 1419 2130 1451 2144
rect 1202 2006 1232 2040
rect 1419 1904 1451 1918
rect 1638 2006 1668 2040
rect 1419 1860 1451 1874
rect 1202 1736 1232 1770
rect 1419 1634 1451 1648
rect 1638 1736 1668 1770
rect 1419 1590 1451 1604
rect 1202 1466 1232 1500
rect 1419 1364 1451 1378
rect 1638 1466 1668 1500
rect 1419 1320 1451 1334
rect 1202 1196 1232 1230
rect 1419 1094 1451 1108
rect 1638 1196 1668 1230
rect 1419 1050 1451 1064
rect 1202 926 1232 960
rect 1419 824 1451 838
rect 1638 926 1668 960
rect 1419 780 1451 794
rect 1202 656 1232 690
rect 1419 554 1451 568
rect 1638 656 1668 690
rect 1419 510 1451 524
rect 1202 386 1232 420
rect 1419 284 1451 298
rect 1638 386 1668 420
rect 1419 240 1451 254
rect 1202 116 1232 150
rect 1419 14 1451 28
rect 1638 116 1668 150
rect 1419 -30 1451 -16
rect 1202 -154 1232 -120
rect 1419 -256 1451 -242
rect 1638 -154 1668 -120
rect 1419 -300 1451 -286
rect 1202 -424 1232 -390
rect 1419 -526 1451 -512
rect 1638 -424 1668 -390
rect 1419 -570 1451 -556
rect 1202 -694 1232 -660
rect 1419 -796 1451 -782
rect 1638 -694 1668 -660
rect 1419 -840 1451 -826
rect 1202 -964 1232 -930
rect 1419 -1066 1451 -1052
rect 1638 -964 1668 -930
rect 1419 -1110 1451 -1096
rect 1202 -1234 1232 -1200
rect 1419 -1336 1451 -1322
rect 1638 -1234 1668 -1200
rect 1419 -1380 1451 -1366
rect 1202 -1504 1232 -1470
rect 1419 -1606 1451 -1592
rect 1638 -1504 1668 -1470
rect 1419 -1650 1451 -1636
rect 1202 -1774 1232 -1740
rect 1419 -1876 1451 -1862
rect 1638 -1774 1668 -1740
rect 1419 -1920 1451 -1906
rect 1202 -2044 1232 -2010
rect 1419 -2146 1451 -2132
rect 1638 -2044 1668 -2010
rect 1999 2130 2031 2144
rect 1782 2006 1812 2040
rect 1999 1904 2031 1918
rect 2218 2006 2248 2040
rect 1999 1860 2031 1874
rect 1782 1736 1812 1770
rect 1999 1634 2031 1648
rect 2218 1736 2248 1770
rect 1999 1590 2031 1604
rect 1782 1466 1812 1500
rect 1999 1364 2031 1378
rect 2218 1466 2248 1500
rect 1999 1320 2031 1334
rect 1782 1196 1812 1230
rect 1999 1094 2031 1108
rect 2218 1196 2248 1230
rect 1999 1050 2031 1064
rect 1782 926 1812 960
rect 1999 824 2031 838
rect 2218 926 2248 960
rect 1999 780 2031 794
rect 1782 656 1812 690
rect 1999 554 2031 568
rect 2218 656 2248 690
rect 1999 510 2031 524
rect 1782 386 1812 420
rect 1999 284 2031 298
rect 2218 386 2248 420
rect 1999 240 2031 254
rect 1782 116 1812 150
rect 1999 14 2031 28
rect 2218 116 2248 150
rect 1999 -30 2031 -16
rect 1782 -154 1812 -120
rect 1999 -256 2031 -242
rect 2218 -154 2248 -120
rect 1999 -300 2031 -286
rect 1782 -424 1812 -390
rect 1999 -526 2031 -512
rect 2218 -424 2248 -390
rect 1999 -570 2031 -556
rect 1782 -694 1812 -660
rect 1999 -796 2031 -782
rect 2218 -694 2248 -660
rect 1999 -840 2031 -826
rect 1782 -964 1812 -930
rect 1999 -1066 2031 -1052
rect 2218 -964 2248 -930
rect 1999 -1110 2031 -1096
rect 1782 -1234 1812 -1200
rect 1999 -1336 2031 -1322
rect 2218 -1234 2248 -1200
rect 1999 -1380 2031 -1366
rect 1782 -1504 1812 -1470
rect 1999 -1606 2031 -1592
rect 2218 -1504 2248 -1470
rect 1999 -1650 2031 -1636
rect 1782 -1774 1812 -1740
rect 1999 -1876 2031 -1862
rect 2218 -1774 2248 -1740
rect 1999 -1920 2031 -1906
rect 1782 -2044 1812 -2010
rect 1999 -2146 2031 -2132
rect 2218 -2044 2248 -2010
rect 2579 2130 2611 2144
rect 2362 2006 2392 2040
rect 2579 1904 2611 1918
rect 2798 2006 2828 2040
rect 2579 1860 2611 1874
rect 2362 1736 2392 1770
rect 2579 1634 2611 1648
rect 2798 1736 2828 1770
rect 2579 1590 2611 1604
rect 2362 1466 2392 1500
rect 2579 1364 2611 1378
rect 2798 1466 2828 1500
rect 2579 1320 2611 1334
rect 2362 1196 2392 1230
rect 2579 1094 2611 1108
rect 2798 1196 2828 1230
rect 2579 1050 2611 1064
rect 2362 926 2392 960
rect 2579 824 2611 838
rect 2798 926 2828 960
rect 2579 780 2611 794
rect 2362 656 2392 690
rect 2579 554 2611 568
rect 2798 656 2828 690
rect 2579 510 2611 524
rect 2362 386 2392 420
rect 2579 284 2611 298
rect 2798 386 2828 420
rect 2579 240 2611 254
rect 2362 116 2392 150
rect 2579 14 2611 28
rect 2798 116 2828 150
rect 2579 -30 2611 -16
rect 2362 -154 2392 -120
rect 2579 -256 2611 -242
rect 2798 -154 2828 -120
rect 2579 -300 2611 -286
rect 2362 -424 2392 -390
rect 2579 -526 2611 -512
rect 2798 -424 2828 -390
rect 2579 -570 2611 -556
rect 2362 -694 2392 -660
rect 2579 -796 2611 -782
rect 2798 -694 2828 -660
rect 2579 -840 2611 -826
rect 2362 -964 2392 -930
rect 2579 -1066 2611 -1052
rect 2798 -964 2828 -930
rect 2579 -1110 2611 -1096
rect 2362 -1234 2392 -1200
rect 2579 -1336 2611 -1322
rect 2798 -1234 2828 -1200
rect 2579 -1380 2611 -1366
rect 2362 -1504 2392 -1470
rect 2579 -1606 2611 -1592
rect 2798 -1504 2828 -1470
rect 2579 -1650 2611 -1636
rect 2362 -1774 2392 -1740
rect 2579 -1876 2611 -1862
rect 2798 -1774 2828 -1740
rect 2579 -1920 2611 -1906
rect 2362 -2044 2392 -2010
rect 2579 -2146 2611 -2132
rect 2798 -2044 2828 -2010
rect 3159 2130 3191 2144
rect 2942 2006 2972 2040
rect 3159 1904 3191 1918
rect 3378 2006 3408 2040
rect 3159 1860 3191 1874
rect 2942 1736 2972 1770
rect 3159 1634 3191 1648
rect 3378 1736 3408 1770
rect 3159 1590 3191 1604
rect 2942 1466 2972 1500
rect 3159 1364 3191 1378
rect 3378 1466 3408 1500
rect 3159 1320 3191 1334
rect 2942 1196 2972 1230
rect 3159 1094 3191 1108
rect 3378 1196 3408 1230
rect 3159 1050 3191 1064
rect 2942 926 2972 960
rect 3159 824 3191 838
rect 3378 926 3408 960
rect 3159 780 3191 794
rect 2942 656 2972 690
rect 3159 554 3191 568
rect 3378 656 3408 690
rect 3159 510 3191 524
rect 2942 386 2972 420
rect 3159 284 3191 298
rect 3378 386 3408 420
rect 3159 240 3191 254
rect 2942 116 2972 150
rect 3159 14 3191 28
rect 3378 116 3408 150
rect 3159 -30 3191 -16
rect 2942 -154 2972 -120
rect 3159 -256 3191 -242
rect 3378 -154 3408 -120
rect 3159 -300 3191 -286
rect 2942 -424 2972 -390
rect 3159 -526 3191 -512
rect 3378 -424 3408 -390
rect 3159 -570 3191 -556
rect 2942 -694 2972 -660
rect 3159 -796 3191 -782
rect 3378 -694 3408 -660
rect 3159 -840 3191 -826
rect 2942 -964 2972 -930
rect 3159 -1066 3191 -1052
rect 3378 -964 3408 -930
rect 3159 -1110 3191 -1096
rect 2942 -1234 2972 -1200
rect 3159 -1336 3191 -1322
rect 3378 -1234 3408 -1200
rect 3159 -1380 3191 -1366
rect 2942 -1504 2972 -1470
rect 3159 -1606 3191 -1592
rect 3378 -1504 3408 -1470
rect 3159 -1650 3191 -1636
rect 2942 -1774 2972 -1740
rect 3159 -1876 3191 -1862
rect 3378 -1774 3408 -1740
rect 3159 -1920 3191 -1906
rect 2942 -2044 2972 -2010
rect 3159 -2146 3191 -2132
rect 3378 -2044 3408 -2010
rect 3739 2130 3771 2144
rect 3522 2006 3552 2040
rect 3739 1904 3771 1918
rect 3958 2006 3988 2040
rect 3739 1860 3771 1874
rect 3522 1736 3552 1770
rect 3739 1634 3771 1648
rect 3958 1736 3988 1770
rect 3739 1590 3771 1604
rect 3522 1466 3552 1500
rect 3739 1364 3771 1378
rect 3958 1466 3988 1500
rect 3739 1320 3771 1334
rect 3522 1196 3552 1230
rect 3739 1094 3771 1108
rect 3958 1196 3988 1230
rect 3739 1050 3771 1064
rect 3522 926 3552 960
rect 3739 824 3771 838
rect 3958 926 3988 960
rect 3739 780 3771 794
rect 3522 656 3552 690
rect 3739 554 3771 568
rect 3958 656 3988 690
rect 3739 510 3771 524
rect 3522 386 3552 420
rect 3739 284 3771 298
rect 3958 386 3988 420
rect 3739 240 3771 254
rect 3522 116 3552 150
rect 3739 14 3771 28
rect 3958 116 3988 150
rect 3739 -30 3771 -16
rect 3522 -154 3552 -120
rect 3739 -256 3771 -242
rect 3958 -154 3988 -120
rect 3739 -300 3771 -286
rect 3522 -424 3552 -390
rect 3739 -526 3771 -512
rect 3958 -424 3988 -390
rect 3739 -570 3771 -556
rect 3522 -694 3552 -660
rect 3739 -796 3771 -782
rect 3958 -694 3988 -660
rect 3739 -840 3771 -826
rect 3522 -964 3552 -930
rect 3739 -1066 3771 -1052
rect 3958 -964 3988 -930
rect 3739 -1110 3771 -1096
rect 3522 -1234 3552 -1200
rect 3739 -1336 3771 -1322
rect 3958 -1234 3988 -1200
rect 3739 -1380 3771 -1366
rect 3522 -1504 3552 -1470
rect 3739 -1606 3771 -1592
rect 3958 -1504 3988 -1470
rect 3739 -1650 3771 -1636
rect 3522 -1774 3552 -1740
rect 3739 -1876 3771 -1862
rect 3958 -1774 3988 -1740
rect 3739 -1920 3771 -1906
rect 3522 -2044 3552 -2010
rect 3739 -2146 3771 -2132
rect 3958 -2044 3988 -2010
rect 4319 2130 4351 2144
rect 4102 2006 4132 2040
rect 4319 1904 4351 1918
rect 4538 2006 4568 2040
rect 4319 1860 4351 1874
rect 4102 1736 4132 1770
rect 4319 1634 4351 1648
rect 4538 1736 4568 1770
rect 4319 1590 4351 1604
rect 4102 1466 4132 1500
rect 4319 1364 4351 1378
rect 4538 1466 4568 1500
rect 4319 1320 4351 1334
rect 4102 1196 4132 1230
rect 4319 1094 4351 1108
rect 4538 1196 4568 1230
rect 4319 1050 4351 1064
rect 4102 926 4132 960
rect 4319 824 4351 838
rect 4538 926 4568 960
rect 4319 780 4351 794
rect 4102 656 4132 690
rect 4319 554 4351 568
rect 4538 656 4568 690
rect 4319 510 4351 524
rect 4102 386 4132 420
rect 4319 284 4351 298
rect 4538 386 4568 420
rect 4319 240 4351 254
rect 4102 116 4132 150
rect 4319 14 4351 28
rect 4538 116 4568 150
rect 4319 -30 4351 -16
rect 4102 -154 4132 -120
rect 4319 -256 4351 -242
rect 4538 -154 4568 -120
rect 4319 -300 4351 -286
rect 4102 -424 4132 -390
rect 4319 -526 4351 -512
rect 4538 -424 4568 -390
rect 4319 -570 4351 -556
rect 4102 -694 4132 -660
rect 4319 -796 4351 -782
rect 4538 -694 4568 -660
rect 4319 -840 4351 -826
rect 4102 -964 4132 -930
rect 4319 -1066 4351 -1052
rect 4538 -964 4568 -930
rect 4319 -1110 4351 -1096
rect 4102 -1234 4132 -1200
rect 4319 -1336 4351 -1322
rect 4538 -1234 4568 -1200
rect 4319 -1380 4351 -1366
rect 4102 -1504 4132 -1470
rect 4319 -1606 4351 -1592
rect 4538 -1504 4568 -1470
rect 4319 -1650 4351 -1636
rect 4102 -1774 4132 -1740
rect 4319 -1876 4351 -1862
rect 4538 -1774 4568 -1740
rect 4319 -1920 4351 -1906
rect 4102 -2044 4132 -2010
rect 4319 -2146 4351 -2132
rect 4538 -2044 4568 -2010
rect 4899 2130 4931 2144
rect 4682 2006 4712 2040
rect 4899 1904 4931 1918
rect 5118 2006 5148 2040
rect 4899 1860 4931 1874
rect 4682 1736 4712 1770
rect 4899 1634 4931 1648
rect 5118 1736 5148 1770
rect 4899 1590 4931 1604
rect 4682 1466 4712 1500
rect 4899 1364 4931 1378
rect 5118 1466 5148 1500
rect 4899 1320 4931 1334
rect 4682 1196 4712 1230
rect 4899 1094 4931 1108
rect 5118 1196 5148 1230
rect 4899 1049 4931 1063
rect 4682 925 4712 959
rect 4899 823 4931 837
rect 5118 925 5148 959
rect 4899 779 4931 793
rect 4682 655 4712 689
rect 4899 553 4931 567
rect 5118 655 5148 689
rect 4899 509 4931 523
rect 4682 385 4712 419
rect 4899 283 4931 297
rect 5118 385 5148 419
rect 4899 239 4931 253
rect 4682 115 4712 149
rect 4899 13 4931 27
rect 5118 115 5148 149
rect 4899 -31 4931 -17
rect 4682 -155 4712 -121
rect 4899 -257 4931 -243
rect 5118 -155 5148 -121
rect 4899 -301 4931 -287
rect 4682 -425 4712 -391
rect 4899 -527 4931 -513
rect 5118 -425 5148 -391
rect 4899 -571 4931 -557
rect 4682 -695 4712 -661
rect 4899 -797 4931 -783
rect 5118 -695 5148 -661
rect 4899 -841 4931 -827
rect 4682 -965 4712 -931
rect 4899 -1067 4931 -1053
rect 5118 -965 5148 -931
rect 4899 -1111 4931 -1097
rect 4682 -1235 4712 -1201
rect 4899 -1337 4931 -1323
rect 5118 -1235 5148 -1201
rect 4899 -1381 4931 -1367
rect 4682 -1505 4712 -1471
rect 4899 -1607 4931 -1593
rect 5118 -1505 5148 -1471
rect 4899 -1651 4931 -1637
rect 4682 -1775 4712 -1741
rect 4899 -1877 4931 -1863
rect 5118 -1775 5148 -1741
rect 4899 -1921 4931 -1907
rect 4682 -2045 4712 -2011
rect 4899 -2147 4931 -2133
rect 5118 -2045 5148 -2011
rect 5479 2130 5511 2144
rect 5262 2006 5292 2040
rect 5479 1904 5511 1918
rect 5698 2006 5728 2040
rect 5479 1860 5511 1874
rect 5262 1736 5292 1770
rect 5479 1634 5511 1648
rect 5698 1736 5728 1770
rect 5479 1590 5511 1604
rect 5262 1466 5292 1500
rect 5479 1364 5511 1378
rect 5698 1466 5728 1500
rect 5479 1320 5511 1334
rect 5262 1196 5292 1230
rect 5479 1094 5511 1108
rect 5698 1196 5728 1230
rect 5479 1049 5511 1063
rect 5262 925 5292 959
rect 5479 823 5511 837
rect 5698 925 5728 959
rect 5479 779 5511 793
rect 5262 655 5292 689
rect 5479 553 5511 567
rect 5698 655 5728 689
rect 5479 509 5511 523
rect 5262 385 5292 419
rect 5479 283 5511 297
rect 5698 385 5728 419
rect 5479 239 5511 253
rect 5262 115 5292 149
rect 5479 13 5511 27
rect 5698 115 5728 149
rect 5479 -31 5511 -17
rect 5262 -155 5292 -121
rect 5479 -257 5511 -243
rect 5698 -155 5728 -121
rect 5479 -301 5511 -287
rect 5262 -425 5292 -391
rect 5479 -527 5511 -513
rect 5698 -425 5728 -391
rect 5479 -571 5511 -557
rect 5262 -695 5292 -661
rect 5479 -797 5511 -783
rect 5698 -695 5728 -661
rect 5479 -841 5511 -827
rect 5262 -965 5292 -931
rect 5479 -1067 5511 -1053
rect 5698 -965 5728 -931
rect 5479 -1111 5511 -1097
rect 5262 -1235 5292 -1201
rect 5479 -1337 5511 -1323
rect 5698 -1235 5728 -1201
rect 5479 -1381 5511 -1367
rect 5262 -1505 5292 -1471
rect 5479 -1607 5511 -1593
rect 5698 -1505 5728 -1471
rect 5479 -1651 5511 -1637
rect 5262 -1775 5292 -1741
rect 5479 -1877 5511 -1863
rect 5698 -1775 5728 -1741
rect 5479 -1921 5511 -1907
rect 5262 -2045 5292 -2011
rect 5479 -2147 5511 -2133
rect 5698 -2045 5728 -2011
rect 6059 2130 6091 2144
rect 5842 2006 5872 2040
rect 6059 1904 6091 1918
rect 6278 2006 6308 2040
rect 6059 1860 6091 1874
rect 5842 1736 5872 1770
rect 6059 1634 6091 1648
rect 6278 1736 6308 1770
rect 6059 1590 6091 1604
rect 5842 1466 5872 1500
rect 6059 1364 6091 1378
rect 6278 1466 6308 1500
rect 6059 1320 6091 1334
rect 5842 1196 5872 1230
rect 6059 1094 6091 1108
rect 6278 1196 6308 1230
rect 6059 1049 6091 1063
rect 5842 925 5872 959
rect 6059 823 6091 837
rect 6278 925 6308 959
rect 6059 779 6091 793
rect 5842 655 5872 689
rect 6059 553 6091 567
rect 6278 655 6308 689
rect 6059 509 6091 523
rect 5842 385 5872 419
rect 6059 283 6091 297
rect 6278 385 6308 419
rect 6059 239 6091 253
rect 5842 115 5872 149
rect 6059 13 6091 27
rect 6278 115 6308 149
rect 6059 -31 6091 -17
rect 5842 -155 5872 -121
rect 6059 -257 6091 -243
rect 6278 -155 6308 -121
rect 6059 -301 6091 -287
rect 5842 -425 5872 -391
rect 6059 -527 6091 -513
rect 6278 -425 6308 -391
rect 6059 -571 6091 -557
rect 5842 -695 5872 -661
rect 6059 -797 6091 -783
rect 6278 -695 6308 -661
rect 6059 -841 6091 -827
rect 5842 -965 5872 -931
rect 6059 -1067 6091 -1053
rect 6278 -965 6308 -931
rect 6059 -1111 6091 -1097
rect 5842 -1235 5872 -1201
rect 6059 -1337 6091 -1323
rect 6278 -1235 6308 -1201
rect 6059 -1381 6091 -1367
rect 5842 -1505 5872 -1471
rect 6059 -1607 6091 -1593
rect 6278 -1505 6308 -1471
rect 6059 -1651 6091 -1637
rect 5842 -1775 5872 -1741
rect 6059 -1877 6091 -1863
rect 6278 -1775 6308 -1741
rect 6059 -1921 6091 -1907
rect 5842 -2045 5872 -2011
rect 6059 -2147 6091 -2133
rect 6278 -2045 6308 -2011
rect 6639 2130 6671 2144
rect 6422 2006 6452 2040
rect 6639 1904 6671 1918
rect 6858 2006 6888 2040
rect 6639 1860 6671 1874
rect 6422 1736 6452 1770
rect 6639 1634 6671 1648
rect 6858 1736 6888 1770
rect 6639 1590 6671 1604
rect 6422 1466 6452 1500
rect 6639 1364 6671 1378
rect 6858 1466 6888 1500
rect 6639 1320 6671 1334
rect 6422 1196 6452 1230
rect 6639 1094 6671 1108
rect 6858 1196 6888 1230
rect 6639 1049 6671 1063
rect 6422 925 6452 959
rect 6639 823 6671 837
rect 6858 925 6888 959
rect 6639 779 6671 793
rect 6422 655 6452 689
rect 6639 553 6671 567
rect 6858 655 6888 689
rect 6639 509 6671 523
rect 6422 385 6452 419
rect 6639 283 6671 297
rect 6858 385 6888 419
rect 6639 239 6671 253
rect 6422 115 6452 149
rect 6639 13 6671 27
rect 6858 115 6888 149
rect 6639 -31 6671 -17
rect 6422 -155 6452 -121
rect 6639 -257 6671 -243
rect 6858 -155 6888 -121
rect 6639 -301 6671 -287
rect 6422 -425 6452 -391
rect 6639 -527 6671 -513
rect 6858 -425 6888 -391
rect 6639 -571 6671 -557
rect 6422 -695 6452 -661
rect 6639 -797 6671 -783
rect 6858 -695 6888 -661
rect 6639 -841 6671 -827
rect 6422 -965 6452 -931
rect 6639 -1067 6671 -1053
rect 6858 -965 6888 -931
rect 6639 -1111 6671 -1097
rect 6422 -1235 6452 -1201
rect 6639 -1337 6671 -1323
rect 6858 -1235 6888 -1201
rect 6639 -1381 6671 -1367
rect 6422 -1505 6452 -1471
rect 6639 -1607 6671 -1593
rect 6858 -1505 6888 -1471
rect 6639 -1651 6671 -1637
rect 6422 -1775 6452 -1741
rect 6639 -1877 6671 -1863
rect 6858 -1775 6888 -1741
rect 6639 -1921 6671 -1907
rect 6422 -2045 6452 -2011
rect 6639 -2147 6671 -2133
rect 6858 -2045 6888 -2011
<< metal1 >>
rect -1 2130 259 2144
rect 291 2130 839 2144
rect 871 2130 1419 2144
rect 1451 2130 1999 2144
rect 2031 2130 2579 2144
rect 2611 2130 3159 2144
rect 3191 2130 3739 2144
rect 3771 2130 4319 2144
rect 4351 2130 4899 2144
rect 4931 2130 5479 2144
rect 5511 2130 6059 2144
rect 6091 2130 6639 2144
rect 6671 2130 6931 2144
rect -1 2006 42 2040
rect 72 2006 478 2040
rect 508 2006 622 2040
rect 652 2006 1058 2040
rect 1088 2006 1202 2040
rect 1232 2006 1638 2040
rect 1668 2006 1782 2040
rect 1812 2006 2218 2040
rect 2248 2006 2362 2040
rect 2392 2006 2798 2040
rect 2828 2006 2942 2040
rect 2972 2006 3378 2040
rect 3408 2006 3522 2040
rect 3552 2006 3958 2040
rect 3988 2006 4102 2040
rect 4132 2006 4538 2040
rect 4568 2006 4682 2040
rect 4712 2006 5118 2040
rect 5148 2006 5262 2040
rect 5292 2006 5698 2040
rect 5728 2006 5842 2040
rect 5872 2006 6278 2040
rect 6308 2006 6422 2040
rect 6452 2006 6858 2040
rect 6888 2006 6931 2040
rect -1 1904 259 1918
rect 291 1904 839 1918
rect 871 1904 1419 1918
rect 1451 1904 1999 1918
rect 2031 1904 2579 1918
rect 2611 1904 3159 1918
rect 3191 1904 3739 1918
rect 3771 1904 4319 1918
rect 4351 1904 4899 1918
rect 4931 1904 5479 1918
rect 5511 1904 6059 1918
rect 6091 1904 6639 1918
rect 6671 1904 6931 1918
rect -1 1860 259 1874
rect 291 1860 839 1874
rect 871 1860 1419 1874
rect 1451 1860 1999 1874
rect 2031 1860 2579 1874
rect 2611 1860 3159 1874
rect 3191 1860 3739 1874
rect 3771 1860 4319 1874
rect 4351 1860 4899 1874
rect 4931 1860 5479 1874
rect 5511 1860 6059 1874
rect 6091 1860 6639 1874
rect 6671 1860 6931 1874
rect -1 1736 42 1770
rect 72 1736 478 1770
rect 508 1736 622 1770
rect 652 1736 1058 1770
rect 1088 1736 1202 1770
rect 1232 1736 1638 1770
rect 1668 1736 1782 1770
rect 1812 1736 2218 1770
rect 2248 1736 2362 1770
rect 2392 1736 2798 1770
rect 2828 1736 2942 1770
rect 2972 1736 3378 1770
rect 3408 1736 3522 1770
rect 3552 1736 3958 1770
rect 3988 1736 4102 1770
rect 4132 1736 4538 1770
rect 4568 1736 4682 1770
rect 4712 1736 5118 1770
rect 5148 1736 5262 1770
rect 5292 1736 5698 1770
rect 5728 1736 5842 1770
rect 5872 1736 6278 1770
rect 6308 1736 6422 1770
rect 6452 1736 6858 1770
rect 6888 1736 6931 1770
rect -1 1634 259 1648
rect 291 1634 839 1648
rect 871 1634 1419 1648
rect 1451 1634 1999 1648
rect 2031 1634 2579 1648
rect 2611 1634 3159 1648
rect 3191 1634 3739 1648
rect 3771 1634 4319 1648
rect 4351 1634 4899 1648
rect 4931 1634 5479 1648
rect 5511 1634 6059 1648
rect 6091 1634 6639 1648
rect 6671 1634 6931 1648
rect -1 1590 259 1604
rect 291 1590 839 1604
rect 871 1590 1419 1604
rect 1451 1590 1999 1604
rect 2031 1590 2579 1604
rect 2611 1590 3159 1604
rect 3191 1590 3739 1604
rect 3771 1590 4319 1604
rect 4351 1590 4899 1604
rect 4931 1590 5479 1604
rect 5511 1590 6059 1604
rect 6091 1590 6639 1604
rect 6671 1590 6931 1604
rect -1 1466 42 1500
rect 72 1466 478 1500
rect 508 1466 622 1500
rect 652 1466 1058 1500
rect 1088 1466 1202 1500
rect 1232 1466 1638 1500
rect 1668 1466 1782 1500
rect 1812 1466 2218 1500
rect 2248 1466 2362 1500
rect 2392 1466 2798 1500
rect 2828 1466 2942 1500
rect 2972 1466 3378 1500
rect 3408 1466 3522 1500
rect 3552 1466 3958 1500
rect 3988 1466 4102 1500
rect 4132 1466 4538 1500
rect 4591 1466 4682 1500
rect 4712 1466 5118 1500
rect 5148 1466 5262 1500
rect 5292 1466 5698 1500
rect 5728 1466 5842 1500
rect 5872 1466 6278 1500
rect 6308 1466 6422 1500
rect 6452 1466 6858 1500
rect 6888 1466 6931 1500
rect -1 1364 259 1378
rect 291 1364 839 1378
rect 871 1364 1419 1378
rect 1451 1364 1999 1378
rect 2031 1364 2579 1378
rect 2611 1364 3159 1378
rect 3191 1364 3739 1378
rect 3771 1364 4319 1378
rect 4351 1364 4899 1378
rect 4931 1364 5479 1378
rect 5511 1364 6059 1378
rect 6091 1364 6639 1378
rect 6671 1364 6931 1378
rect -1 1320 259 1334
rect 291 1320 839 1334
rect 871 1320 1419 1334
rect 1451 1320 1999 1334
rect 2031 1320 2579 1334
rect 2611 1320 3159 1334
rect 3191 1320 3739 1334
rect 3771 1320 4319 1334
rect 4351 1320 4899 1334
rect 4931 1320 5479 1334
rect 5511 1320 6059 1334
rect 6091 1320 6639 1334
rect 6671 1320 6931 1334
rect -1 1196 42 1230
rect 72 1196 478 1230
rect 508 1196 622 1230
rect 652 1196 1058 1230
rect 1088 1196 1202 1230
rect 1232 1196 1638 1230
rect 1668 1196 1782 1230
rect 1812 1196 2218 1230
rect 2248 1196 2362 1230
rect 2392 1196 2798 1230
rect 2828 1196 2942 1230
rect 2972 1196 3378 1230
rect 3408 1196 3522 1230
rect 3552 1196 3958 1230
rect 3988 1196 4102 1230
rect 4132 1196 4538 1230
rect 4591 1196 4682 1230
rect 4712 1196 5118 1230
rect 5148 1196 5262 1230
rect 5292 1196 5698 1230
rect 5728 1196 5842 1230
rect 5872 1196 6278 1230
rect 6308 1196 6422 1230
rect 6452 1196 6858 1230
rect 6888 1196 6931 1230
rect -1 1094 259 1108
rect 291 1094 839 1108
rect 871 1094 1419 1108
rect 1451 1094 1999 1108
rect 2031 1094 2579 1108
rect 2611 1094 3159 1108
rect 3191 1094 3739 1108
rect 3771 1094 4319 1108
rect 4351 1094 4899 1108
rect 4931 1094 5479 1108
rect 5511 1094 6059 1108
rect 6091 1094 6639 1108
rect 6671 1094 6931 1108
rect -1 1050 259 1064
rect 291 1050 839 1064
rect 871 1050 1419 1064
rect 1451 1050 1999 1064
rect 2031 1050 2579 1064
rect 2611 1050 3159 1064
rect 3191 1050 3739 1064
rect 3771 1050 4319 1064
rect 4351 1063 4611 1064
rect 4351 1050 4899 1063
rect 4591 1049 4899 1050
rect 4931 1049 5479 1063
rect 5511 1049 6059 1063
rect 6091 1049 6639 1063
rect 6671 1049 6931 1063
rect -1 926 42 960
rect 72 926 478 960
rect 508 926 622 960
rect 652 926 1058 960
rect 1088 926 1202 960
rect 1232 926 1638 960
rect 1668 926 1782 960
rect 1812 926 2218 960
rect 2248 926 2362 960
rect 2392 926 2798 960
rect 2828 926 2942 960
rect 2972 926 3378 960
rect 3408 926 3522 960
rect 3552 926 3958 960
rect 3988 926 4102 960
rect 4132 926 4538 960
rect 4591 925 4682 959
rect 4712 925 5118 959
rect 5148 925 5262 959
rect 5292 925 5698 959
rect 5728 925 5842 959
rect 5872 925 6278 959
rect 6308 925 6422 959
rect 6452 925 6858 959
rect 6888 925 6931 959
rect -1 824 259 838
rect 291 824 839 838
rect 871 824 1419 838
rect 1451 824 1999 838
rect 2031 824 2579 838
rect 2611 824 3159 838
rect 3191 824 3739 838
rect 3771 824 4319 838
rect 4351 837 4611 838
rect 4351 824 4899 837
rect 4591 823 4899 824
rect 4931 823 5479 837
rect 5511 823 6059 837
rect 6091 823 6639 837
rect 6671 823 6931 837
rect -1 780 259 794
rect 291 780 839 794
rect 871 780 1419 794
rect 1451 780 1999 794
rect 2031 780 2579 794
rect 2611 780 3159 794
rect 3191 780 3739 794
rect 3771 780 4319 794
rect 4351 793 4611 794
rect 4351 780 4899 793
rect 4591 779 4899 780
rect 4931 779 5479 793
rect 5511 779 6059 793
rect 6091 779 6639 793
rect 6671 779 6931 793
rect -1 656 42 690
rect 72 656 478 690
rect 508 656 622 690
rect 652 656 1058 690
rect 1088 656 1202 690
rect 1232 656 1638 690
rect 1668 656 1782 690
rect 1812 656 2218 690
rect 2248 656 2362 690
rect 2392 656 2798 690
rect 2828 656 2942 690
rect 2972 656 3378 690
rect 3408 656 3522 690
rect 3552 656 3958 690
rect 3988 656 4102 690
rect 4132 656 4538 690
rect 4591 655 4682 689
rect 4712 655 5118 689
rect 5148 655 5262 689
rect 5292 655 5698 689
rect 5728 655 5842 689
rect 5872 655 6278 689
rect 6308 655 6422 689
rect 6452 655 6858 689
rect 6888 655 6931 689
rect -1 554 259 568
rect 291 554 839 568
rect 871 554 1419 568
rect 1451 554 1999 568
rect 2031 554 2579 568
rect 2611 554 3159 568
rect 3191 554 3739 568
rect 3771 554 4319 568
rect 4351 567 4611 568
rect 4351 554 4899 567
rect 4591 553 4899 554
rect 4931 553 5479 567
rect 5511 553 6059 567
rect 6091 553 6639 567
rect 6671 553 6931 567
rect -1 510 259 524
rect 291 510 839 524
rect 871 510 1419 524
rect 1451 510 1999 524
rect 2031 510 2579 524
rect 2611 510 3159 524
rect 3191 510 3739 524
rect 3771 510 4319 524
rect 4351 523 4611 524
rect 4351 510 4899 523
rect 4591 509 4899 510
rect 4931 509 5479 523
rect 5511 509 6059 523
rect 6091 509 6639 523
rect 6671 509 6931 523
rect -1 386 42 420
rect 72 386 478 420
rect 508 386 622 420
rect 652 386 1058 420
rect 1088 386 1202 420
rect 1232 386 1638 420
rect 1668 386 1782 420
rect 1812 386 2218 420
rect 2248 386 2362 420
rect 2392 386 2798 420
rect 2828 386 2942 420
rect 2972 386 3378 420
rect 3408 386 3522 420
rect 3552 386 3958 420
rect 3988 386 4102 420
rect 4132 386 4538 420
rect 4591 385 4682 419
rect 4712 385 5118 419
rect 5148 385 5262 419
rect 5292 385 5698 419
rect 5728 385 5842 419
rect 5872 385 6278 419
rect 6308 385 6422 419
rect 6452 385 6858 419
rect 6888 385 6931 419
rect -1 284 259 298
rect 291 284 839 298
rect 871 284 1419 298
rect 1451 284 1999 298
rect 2031 284 2579 298
rect 2611 284 3159 298
rect 3191 284 3739 298
rect 3771 284 4319 298
rect 4351 297 4611 298
rect 4351 284 4899 297
rect 4591 283 4899 284
rect 4931 283 5479 297
rect 5511 283 6059 297
rect 6091 283 6639 297
rect 6671 283 6931 297
rect -1 240 259 254
rect 291 240 839 254
rect 871 240 1419 254
rect 1451 240 1999 254
rect 2031 240 2579 254
rect 2611 240 3159 254
rect 3191 240 3739 254
rect 3771 240 4319 254
rect 4351 253 4611 254
rect 4351 240 4899 253
rect 4591 239 4899 240
rect 4931 239 5479 253
rect 5511 239 6059 253
rect 6091 239 6639 253
rect 6671 239 6931 253
rect -1 116 42 150
rect 72 116 478 150
rect 508 116 622 150
rect 652 116 1058 150
rect 1088 116 1202 150
rect 1232 116 1638 150
rect 1668 116 1782 150
rect 1812 116 2218 150
rect 2248 116 2362 150
rect 2392 116 2798 150
rect 2828 116 2942 150
rect 2972 116 3378 150
rect 3408 116 3522 150
rect 3552 116 3958 150
rect 3988 116 4102 150
rect 4132 116 4538 150
rect 4591 115 4682 149
rect 4712 115 5118 149
rect 5148 115 5262 149
rect 5292 115 5698 149
rect 5728 115 5842 149
rect 5872 115 6278 149
rect 6308 115 6422 149
rect 6452 115 6858 149
rect 6888 115 6931 149
rect -1 14 259 28
rect 291 14 839 28
rect 871 14 1419 28
rect 1451 14 1999 28
rect 2031 14 2579 28
rect 2611 14 3159 28
rect 3191 14 3739 28
rect 3771 14 4319 28
rect 4351 27 4611 28
rect 4351 14 4899 27
rect 4591 13 4899 14
rect 4931 13 5479 27
rect 5511 13 6059 27
rect 6091 13 6639 27
rect 6671 13 6931 27
rect -1 -30 259 -16
rect 291 -30 839 -16
rect 871 -30 1419 -16
rect 1451 -30 1999 -16
rect 2031 -30 2579 -16
rect 2611 -30 3159 -16
rect 3191 -30 3739 -16
rect 3771 -30 4319 -16
rect 4351 -17 4611 -16
rect 4351 -30 4899 -17
rect 4591 -31 4899 -30
rect 4931 -31 5479 -17
rect 5511 -31 6059 -17
rect 6091 -31 6639 -17
rect 6671 -31 6931 -17
rect -1 -154 42 -120
rect 72 -154 478 -120
rect 508 -154 622 -120
rect 652 -154 1058 -120
rect 1088 -154 1202 -120
rect 1232 -154 1638 -120
rect 1668 -154 1782 -120
rect 1812 -154 2218 -120
rect 2248 -154 2362 -120
rect 2392 -154 2798 -120
rect 2828 -154 2942 -120
rect 2972 -154 3378 -120
rect 3408 -154 3522 -120
rect 3552 -154 3958 -120
rect 3988 -154 4102 -120
rect 4132 -154 4538 -120
rect 4591 -155 4682 -121
rect 4712 -155 5118 -121
rect 5148 -155 5262 -121
rect 5292 -155 5698 -121
rect 5728 -155 5842 -121
rect 5872 -155 6278 -121
rect 6308 -155 6422 -121
rect 6452 -155 6858 -121
rect 6888 -155 6931 -121
rect -1 -256 259 -242
rect 291 -256 839 -242
rect 871 -256 1419 -242
rect 1451 -256 1999 -242
rect 2031 -256 2579 -242
rect 2611 -256 3159 -242
rect 3191 -256 3739 -242
rect 3771 -256 4319 -242
rect 4351 -243 4611 -242
rect 4351 -256 4899 -243
rect 4591 -257 4899 -256
rect 4931 -257 5479 -243
rect 5511 -257 6059 -243
rect 6091 -257 6639 -243
rect 6671 -257 6931 -243
rect -1 -300 259 -286
rect 291 -300 839 -286
rect 871 -300 1419 -286
rect 1451 -300 1999 -286
rect 2031 -300 2579 -286
rect 2611 -300 3159 -286
rect 3191 -300 3739 -286
rect 3771 -300 4319 -286
rect 4351 -287 4611 -286
rect 4351 -300 4899 -287
rect 4591 -301 4899 -300
rect 4931 -301 5479 -287
rect 5511 -301 6059 -287
rect 6091 -301 6639 -287
rect 6671 -301 6931 -287
rect -1 -424 42 -390
rect 72 -424 478 -390
rect 508 -424 622 -390
rect 652 -424 1058 -390
rect 1088 -424 1202 -390
rect 1232 -424 1638 -390
rect 1668 -424 1782 -390
rect 1812 -424 2218 -390
rect 2248 -424 2362 -390
rect 2392 -424 2798 -390
rect 2828 -424 2942 -390
rect 2972 -424 3378 -390
rect 3408 -424 3522 -390
rect 3552 -424 3958 -390
rect 3988 -424 4102 -390
rect 4132 -424 4538 -390
rect 4591 -425 4682 -391
rect 4712 -425 5118 -391
rect 5148 -425 5262 -391
rect 5292 -425 5698 -391
rect 5728 -425 5842 -391
rect 5872 -425 6278 -391
rect 6308 -425 6422 -391
rect 6452 -425 6858 -391
rect 6888 -425 6931 -391
rect -1 -526 259 -512
rect 291 -526 839 -512
rect 871 -526 1419 -512
rect 1451 -526 1999 -512
rect 2031 -526 2579 -512
rect 2611 -526 3159 -512
rect 3191 -526 3739 -512
rect 3771 -526 4319 -512
rect 4351 -513 4611 -512
rect 4351 -526 4899 -513
rect 4591 -527 4899 -526
rect 4931 -527 5479 -513
rect 5511 -527 6059 -513
rect 6091 -527 6639 -513
rect 6671 -527 6931 -513
rect -1 -570 259 -556
rect 291 -570 839 -556
rect 871 -570 1419 -556
rect 1451 -570 1999 -556
rect 2031 -570 2579 -556
rect 2611 -570 3159 -556
rect 3191 -570 3739 -556
rect 3771 -570 4319 -556
rect 4351 -557 4611 -556
rect 4351 -570 4899 -557
rect 4591 -571 4899 -570
rect 4931 -571 5479 -557
rect 5511 -571 6059 -557
rect 6091 -571 6639 -557
rect 6671 -571 6931 -557
rect -1 -694 42 -660
rect 72 -694 478 -660
rect 508 -694 622 -660
rect 652 -694 1058 -660
rect 1088 -694 1202 -660
rect 1232 -694 1638 -660
rect 1668 -694 1782 -660
rect 1812 -694 2218 -660
rect 2248 -694 2362 -660
rect 2392 -694 2798 -660
rect 2828 -694 2942 -660
rect 2972 -694 3378 -660
rect 3408 -694 3522 -660
rect 3552 -694 3958 -660
rect 3988 -694 4102 -660
rect 4132 -694 4538 -660
rect 4591 -695 4682 -661
rect 4712 -695 5118 -661
rect 5148 -695 5262 -661
rect 5292 -695 5698 -661
rect 5728 -695 5842 -661
rect 5872 -695 6278 -661
rect 6308 -695 6422 -661
rect 6452 -695 6858 -661
rect 6888 -695 6931 -661
rect -1 -796 259 -782
rect 291 -796 839 -782
rect 871 -796 1419 -782
rect 1451 -796 1999 -782
rect 2031 -796 2579 -782
rect 2611 -796 3159 -782
rect 3191 -796 3739 -782
rect 3771 -796 4319 -782
rect 4351 -783 4611 -782
rect 4351 -796 4899 -783
rect 4591 -797 4899 -796
rect 4931 -797 5479 -783
rect 5511 -797 6059 -783
rect 6091 -797 6639 -783
rect 6671 -797 6931 -783
rect -1 -840 259 -826
rect 291 -840 839 -826
rect 871 -840 1419 -826
rect 1451 -840 1999 -826
rect 2031 -840 2579 -826
rect 2611 -840 3159 -826
rect 3191 -840 3739 -826
rect 3771 -840 4319 -826
rect 4351 -827 4611 -826
rect 4351 -840 4899 -827
rect 4591 -841 4899 -840
rect 4931 -841 5479 -827
rect 5511 -841 6059 -827
rect 6091 -841 6639 -827
rect 6671 -841 6931 -827
rect -1 -964 42 -930
rect 72 -964 478 -930
rect 508 -964 622 -930
rect 652 -964 1058 -930
rect 1088 -964 1202 -930
rect 1232 -964 1638 -930
rect 1668 -964 1782 -930
rect 1812 -964 2218 -930
rect 2248 -964 2362 -930
rect 2392 -964 2798 -930
rect 2828 -964 2942 -930
rect 2972 -964 3378 -930
rect 3408 -964 3522 -930
rect 3552 -964 3958 -930
rect 3988 -964 4102 -930
rect 4132 -964 4538 -930
rect 4591 -965 4682 -931
rect 4712 -965 5118 -931
rect 5148 -965 5262 -931
rect 5292 -965 5698 -931
rect 5728 -965 5842 -931
rect 5872 -965 6278 -931
rect 6308 -965 6422 -931
rect 6452 -965 6858 -931
rect 6888 -965 6931 -931
rect -1 -1066 259 -1052
rect 291 -1066 839 -1052
rect 871 -1066 1419 -1052
rect 1451 -1066 1999 -1052
rect 2031 -1066 2579 -1052
rect 2611 -1066 3159 -1052
rect 3191 -1066 3739 -1052
rect 3771 -1066 4319 -1052
rect 4351 -1053 4611 -1052
rect 4351 -1066 4899 -1053
rect 4591 -1067 4899 -1066
rect 4931 -1067 5479 -1053
rect 5511 -1067 6059 -1053
rect 6091 -1067 6639 -1053
rect 6671 -1067 6931 -1053
rect -1 -1110 259 -1096
rect 291 -1110 839 -1096
rect 871 -1110 1419 -1096
rect 1451 -1110 1999 -1096
rect 2031 -1110 2579 -1096
rect 2611 -1110 3159 -1096
rect 3191 -1110 3739 -1096
rect 3771 -1110 4319 -1096
rect 4351 -1097 4611 -1096
rect 4351 -1110 4899 -1097
rect 4591 -1111 4899 -1110
rect 4931 -1111 5479 -1097
rect 5511 -1111 6059 -1097
rect 6091 -1111 6639 -1097
rect 6671 -1111 6931 -1097
rect -1 -1234 42 -1200
rect 72 -1234 478 -1200
rect 508 -1234 622 -1200
rect 652 -1234 1058 -1200
rect 1088 -1234 1202 -1200
rect 1232 -1234 1638 -1200
rect 1668 -1234 1782 -1200
rect 1812 -1234 2218 -1200
rect 2248 -1234 2362 -1200
rect 2392 -1234 2798 -1200
rect 2828 -1234 2942 -1200
rect 2972 -1234 3378 -1200
rect 3408 -1234 3522 -1200
rect 3552 -1234 3958 -1200
rect 3988 -1234 4102 -1200
rect 4132 -1234 4538 -1200
rect 4591 -1235 4682 -1201
rect 4712 -1235 5118 -1201
rect 5148 -1235 5262 -1201
rect 5292 -1235 5698 -1201
rect 5728 -1235 5842 -1201
rect 5872 -1235 6278 -1201
rect 6308 -1235 6422 -1201
rect 6452 -1235 6858 -1201
rect 6888 -1235 6931 -1201
rect -1 -1336 259 -1322
rect 291 -1336 839 -1322
rect 871 -1336 1419 -1322
rect 1451 -1336 1999 -1322
rect 2031 -1336 2579 -1322
rect 2611 -1336 3159 -1322
rect 3191 -1336 3739 -1322
rect 3771 -1336 4319 -1322
rect 4351 -1323 4611 -1322
rect 4351 -1336 4899 -1323
rect 4591 -1337 4899 -1336
rect 4931 -1337 5479 -1323
rect 5511 -1337 6059 -1323
rect 6091 -1337 6639 -1323
rect 6671 -1337 6931 -1323
rect -1 -1380 259 -1366
rect 291 -1380 839 -1366
rect 871 -1380 1419 -1366
rect 1451 -1380 1999 -1366
rect 2031 -1380 2579 -1366
rect 2611 -1380 3159 -1366
rect 3191 -1380 3739 -1366
rect 3771 -1380 4319 -1366
rect 4351 -1367 4611 -1366
rect 4351 -1380 4899 -1367
rect 4591 -1381 4899 -1380
rect 4931 -1381 5479 -1367
rect 5511 -1381 6059 -1367
rect 6091 -1381 6639 -1367
rect 6671 -1381 6931 -1367
rect -1 -1504 42 -1470
rect 72 -1504 478 -1470
rect 508 -1504 622 -1470
rect 652 -1504 1058 -1470
rect 1088 -1504 1202 -1470
rect 1232 -1504 1638 -1470
rect 1668 -1504 1782 -1470
rect 1812 -1504 2218 -1470
rect 2248 -1504 2362 -1470
rect 2392 -1504 2798 -1470
rect 2828 -1504 2942 -1470
rect 2972 -1504 3378 -1470
rect 3408 -1504 3522 -1470
rect 3552 -1504 3958 -1470
rect 3988 -1504 4102 -1470
rect 4132 -1504 4538 -1470
rect 4591 -1505 4682 -1471
rect 4712 -1505 5118 -1471
rect 5148 -1505 5262 -1471
rect 5292 -1505 5698 -1471
rect 5728 -1505 5842 -1471
rect 5872 -1505 6278 -1471
rect 6308 -1505 6422 -1471
rect 6452 -1505 6858 -1471
rect 6888 -1505 6931 -1471
rect -1 -1606 259 -1592
rect 291 -1606 839 -1592
rect 871 -1606 1419 -1592
rect 1451 -1606 1999 -1592
rect 2031 -1606 2579 -1592
rect 2611 -1606 3159 -1592
rect 3191 -1606 3739 -1592
rect 3771 -1606 4319 -1592
rect 4351 -1593 4611 -1592
rect 4351 -1606 4899 -1593
rect 4591 -1607 4899 -1606
rect 4931 -1607 5479 -1593
rect 5511 -1607 6059 -1593
rect 6091 -1607 6639 -1593
rect 6671 -1607 6931 -1593
rect -1 -1650 259 -1636
rect 291 -1650 839 -1636
rect 871 -1650 1419 -1636
rect 1451 -1650 1999 -1636
rect 2031 -1650 2579 -1636
rect 2611 -1650 3159 -1636
rect 3191 -1650 3739 -1636
rect 3771 -1650 4319 -1636
rect 4351 -1637 4611 -1636
rect 4351 -1650 4899 -1637
rect 4591 -1651 4899 -1650
rect 4931 -1651 5479 -1637
rect 5511 -1651 6059 -1637
rect 6091 -1651 6639 -1637
rect 6671 -1651 6931 -1637
rect -1 -1774 42 -1740
rect 72 -1774 478 -1740
rect 508 -1774 622 -1740
rect 652 -1774 1058 -1740
rect 1088 -1774 1202 -1740
rect 1232 -1774 1638 -1740
rect 1668 -1774 1782 -1740
rect 1812 -1774 2218 -1740
rect 2248 -1774 2362 -1740
rect 2392 -1774 2798 -1740
rect 2828 -1774 2942 -1740
rect 2972 -1774 3378 -1740
rect 3408 -1774 3522 -1740
rect 3552 -1774 3958 -1740
rect 3988 -1774 4102 -1740
rect 4132 -1774 4538 -1740
rect 4591 -1775 4682 -1741
rect 4712 -1775 5118 -1741
rect 5148 -1775 5262 -1741
rect 5292 -1775 5698 -1741
rect 5728 -1775 5842 -1741
rect 5872 -1775 6278 -1741
rect 6308 -1775 6422 -1741
rect 6452 -1775 6858 -1741
rect 6888 -1775 6931 -1741
rect -1 -1876 259 -1862
rect 291 -1876 839 -1862
rect 871 -1876 1419 -1862
rect 1451 -1876 1999 -1862
rect 2031 -1876 2579 -1862
rect 2611 -1876 3159 -1862
rect 3191 -1876 3739 -1862
rect 3771 -1876 4319 -1862
rect 4351 -1863 4611 -1862
rect 4351 -1876 4899 -1863
rect 4591 -1877 4899 -1876
rect 4931 -1877 5479 -1863
rect 5511 -1877 6059 -1863
rect 6091 -1877 6639 -1863
rect 6671 -1877 6931 -1863
rect -1 -1920 259 -1906
rect 291 -1920 839 -1906
rect 871 -1920 1419 -1906
rect 1451 -1920 1999 -1906
rect 2031 -1920 2579 -1906
rect 2611 -1920 3159 -1906
rect 3191 -1920 3739 -1906
rect 3771 -1920 4319 -1906
rect 4351 -1907 4611 -1906
rect 4351 -1920 4899 -1907
rect 4591 -1921 4899 -1920
rect 4931 -1921 5479 -1907
rect 5511 -1921 6059 -1907
rect 6091 -1921 6639 -1907
rect 6671 -1921 6931 -1907
rect -1 -2044 42 -2010
rect 72 -2044 478 -2010
rect 508 -2044 622 -2010
rect 652 -2044 1058 -2010
rect 1088 -2044 1202 -2010
rect 1232 -2044 1638 -2010
rect 1668 -2044 1782 -2010
rect 1812 -2044 2218 -2010
rect 2248 -2044 2362 -2010
rect 2392 -2044 2798 -2010
rect 2828 -2044 2942 -2010
rect 2972 -2044 3378 -2010
rect 3408 -2044 3522 -2010
rect 3552 -2044 3958 -2010
rect 3988 -2044 4102 -2010
rect 4132 -2044 4538 -2010
rect 4591 -2045 4682 -2011
rect 4712 -2045 5118 -2011
rect 5148 -2045 5262 -2011
rect 5292 -2045 5698 -2011
rect 5728 -2045 5842 -2011
rect 5872 -2045 6278 -2011
rect 6308 -2045 6422 -2011
rect 6452 -2045 6858 -2011
rect 6888 -2045 6931 -2011
rect -1 -2146 259 -2132
rect 291 -2146 839 -2132
rect 871 -2146 1419 -2132
rect 1451 -2146 1999 -2132
rect 2031 -2146 2579 -2132
rect 2611 -2146 3159 -2132
rect 3191 -2146 3739 -2132
rect 3771 -2146 4319 -2132
rect 4351 -2133 4611 -2132
rect 4351 -2146 4899 -2133
rect 4591 -2147 4899 -2146
rect 4931 -2147 5479 -2133
rect 5511 -2147 6059 -2133
rect 6091 -2147 6639 -2133
rect 6671 -2147 6931 -2133
<< labels >>
rlabel poly 4591 523 4621 553 1 10T_4x4_magic_3/WWL_0
rlabel poly 4591 253 4621 283 1 10T_4x4_magic_3/WWL_1
rlabel metal1 4591 509 4621 523 1 10T_4x4_magic_3/VDD
rlabel metal1 4591 239 4621 253 1 10T_4x4_magic_3/VDD
rlabel metal1 4591 283 4621 297 1 10T_4x4_magic_3/GND
rlabel metal1 4591 13 4621 27 1 10T_4x4_magic_3/GND
rlabel corelocali 4639 -35 4654 -5 1 10T_4x4_magic_3/RBL1_0
rlabel corelocali 5176 -35 5191 -5 1 10T_4x4_magic_3/RBL0_0
rlabel corelocali 5219 -35 5234 -5 1 10T_4x4_magic_3/RBL1_1
rlabel corelocali 5756 -35 5771 -5 1 10T_4x4_magic_3/RBL0_1
rlabel metal1 4591 115 4621 149 1 10T_4x4_magic_3/RWL_1
rlabel metal1 4591 385 4621 419 1 10T_4x4_magic_3/RWL_0
rlabel poly 5219 253 5771 283 1 10T_4x4_magic_3/10T_toy_magic_3/WWL
rlabel locali 5698 115 5728 149 1 10T_4x4_magic_3/10T_toy_magic_3/RWL
rlabel locali 5262 115 5292 149 1 10T_4x4_magic_3/10T_toy_magic_3/RWL
rlabel locali 5683 197 5698 226 1 10T_4x4_magic_3/10T_toy_magic_3/WBL
rlabel locali 5293 197 5308 225 1 10T_4x4_magic_3/10T_toy_magic_3/WBLb
rlabel locali 5756 51 5771 93 1 10T_4x4_magic_3/10T_toy_magic_3/RBL0
rlabel locali 5219 51 5234 93 1 10T_4x4_magic_3/10T_toy_magic_3/RBL1
rlabel metal1 5479 239 5511 253 1 10T_4x4_magic_3/10T_toy_magic_3/VDD
rlabel metal1 5479 13 5511 27 7 10T_4x4_magic_3/10T_toy_magic_3/GND
rlabel polycont 5441 120 5471 154 1 10T_4x4_magic_3/10T_toy_magic_3/junc0
rlabel polycont 5519 120 5549 154 1 10T_4x4_magic_3/10T_toy_magic_3/junc1
rlabel ndiff 5292 51 5348 79 1 10T_4x4_magic_3/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 51 5698 79 1 10T_4x4_magic_3/10T_toy_magic_3/RWL0_junc
rlabel poly 4639 253 5191 283 1 10T_4x4_magic_3/10T_toy_magic_2/WWL
rlabel locali 5118 115 5148 149 1 10T_4x4_magic_3/10T_toy_magic_2/RWL
rlabel locali 4682 115 4712 149 1 10T_4x4_magic_3/10T_toy_magic_2/RWL
rlabel locali 5103 197 5118 226 1 10T_4x4_magic_3/10T_toy_magic_2/WBL
rlabel locali 4713 197 4728 225 1 10T_4x4_magic_3/10T_toy_magic_2/WBLb
rlabel locali 5176 51 5191 93 1 10T_4x4_magic_3/10T_toy_magic_2/RBL0
rlabel locali 4639 51 4654 93 1 10T_4x4_magic_3/10T_toy_magic_2/RBL1
rlabel metal1 4899 239 4931 253 1 10T_4x4_magic_3/10T_toy_magic_2/VDD
rlabel metal1 4899 13 4931 27 7 10T_4x4_magic_3/10T_toy_magic_2/GND
rlabel polycont 4861 120 4891 154 1 10T_4x4_magic_3/10T_toy_magic_2/junc0
rlabel polycont 4939 120 4969 154 1 10T_4x4_magic_3/10T_toy_magic_2/junc1
rlabel ndiff 4712 51 4768 79 1 10T_4x4_magic_3/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 51 5118 79 1 10T_4x4_magic_3/10T_toy_magic_2/RWL0_junc
rlabel poly 5219 523 5771 553 1 10T_4x4_magic_3/10T_toy_magic_1/WWL
rlabel locali 5698 385 5728 419 1 10T_4x4_magic_3/10T_toy_magic_1/RWL
rlabel locali 5262 385 5292 419 1 10T_4x4_magic_3/10T_toy_magic_1/RWL
rlabel locali 5683 467 5698 496 1 10T_4x4_magic_3/10T_toy_magic_1/WBL
rlabel locali 5293 467 5308 495 1 10T_4x4_magic_3/10T_toy_magic_1/WBLb
rlabel locali 5756 321 5771 363 1 10T_4x4_magic_3/10T_toy_magic_1/RBL0
rlabel locali 5219 321 5234 363 1 10T_4x4_magic_3/10T_toy_magic_1/RBL1
rlabel metal1 5479 509 5511 523 1 10T_4x4_magic_3/10T_toy_magic_1/VDD
rlabel metal1 5479 283 5511 297 7 10T_4x4_magic_3/10T_toy_magic_1/GND
rlabel polycont 5441 390 5471 424 1 10T_4x4_magic_3/10T_toy_magic_1/junc0
rlabel polycont 5519 390 5549 424 1 10T_4x4_magic_3/10T_toy_magic_1/junc1
rlabel ndiff 5292 321 5348 349 1 10T_4x4_magic_3/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 321 5698 349 1 10T_4x4_magic_3/10T_toy_magic_1/RWL0_junc
rlabel poly 4639 523 5191 553 1 10T_4x4_magic_3/10T_toy_magic_0/WWL
rlabel locali 5118 385 5148 419 1 10T_4x4_magic_3/10T_toy_magic_0/RWL
rlabel locali 4682 385 4712 419 1 10T_4x4_magic_3/10T_toy_magic_0/RWL
rlabel locali 5103 467 5118 496 1 10T_4x4_magic_3/10T_toy_magic_0/WBL
rlabel locali 4713 467 4728 495 1 10T_4x4_magic_3/10T_toy_magic_0/WBLb
rlabel locali 5176 321 5191 363 1 10T_4x4_magic_3/10T_toy_magic_0/RBL0
rlabel locali 4639 321 4654 363 1 10T_4x4_magic_3/10T_toy_magic_0/RBL1
rlabel metal1 4899 509 4931 523 1 10T_4x4_magic_3/10T_toy_magic_0/VDD
rlabel metal1 4899 283 4931 297 7 10T_4x4_magic_3/10T_toy_magic_0/GND
rlabel polycont 4861 390 4891 424 1 10T_4x4_magic_3/10T_toy_magic_0/junc0
rlabel polycont 4939 390 4969 424 1 10T_4x4_magic_3/10T_toy_magic_0/junc1
rlabel ndiff 4712 321 4768 349 1 10T_4x4_magic_3/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 321 5118 349 1 10T_4x4_magic_3/10T_toy_magic_0/RWL0_junc
rlabel poly 4591 -17 4621 13 1 10T_4x4_magic_4/WWL_0
rlabel poly 4591 -287 4621 -257 1 10T_4x4_magic_4/WWL_1
rlabel metal1 4591 -31 4621 -17 1 10T_4x4_magic_4/VDD
rlabel metal1 4591 -301 4621 -287 1 10T_4x4_magic_4/VDD
rlabel metal1 4591 -257 4621 -243 1 10T_4x4_magic_4/GND
rlabel metal1 4591 -527 4621 -513 1 10T_4x4_magic_4/GND
rlabel corelocali 4639 -575 4654 -545 1 10T_4x4_magic_4/RBL1_0
rlabel corelocali 5176 -575 5191 -545 1 10T_4x4_magic_4/RBL0_0
rlabel corelocali 5219 -575 5234 -545 1 10T_4x4_magic_4/RBL1_1
rlabel corelocali 5756 -575 5771 -545 1 10T_4x4_magic_4/RBL0_1
rlabel metal1 4591 -425 4621 -391 1 10T_4x4_magic_4/RWL_1
rlabel metal1 4591 -155 4621 -121 1 10T_4x4_magic_4/RWL_0
rlabel poly 5219 -287 5771 -257 1 10T_4x4_magic_4/10T_toy_magic_3/WWL
rlabel locali 5698 -425 5728 -391 1 10T_4x4_magic_4/10T_toy_magic_3/RWL
rlabel locali 5262 -425 5292 -391 1 10T_4x4_magic_4/10T_toy_magic_3/RWL
rlabel locali 5683 -343 5698 -314 1 10T_4x4_magic_4/10T_toy_magic_3/WBL
rlabel locali 5293 -343 5308 -315 1 10T_4x4_magic_4/10T_toy_magic_3/WBLb
rlabel locali 5756 -489 5771 -447 1 10T_4x4_magic_4/10T_toy_magic_3/RBL0
rlabel locali 5219 -489 5234 -447 1 10T_4x4_magic_4/10T_toy_magic_3/RBL1
rlabel metal1 5479 -301 5511 -287 1 10T_4x4_magic_4/10T_toy_magic_3/VDD
rlabel metal1 5479 -527 5511 -513 7 10T_4x4_magic_4/10T_toy_magic_3/GND
rlabel polycont 5441 -420 5471 -386 1 10T_4x4_magic_4/10T_toy_magic_3/junc0
rlabel polycont 5519 -420 5549 -386 1 10T_4x4_magic_4/10T_toy_magic_3/junc1
rlabel ndiff 5292 -489 5348 -461 1 10T_4x4_magic_4/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 -489 5698 -461 1 10T_4x4_magic_4/10T_toy_magic_3/RWL0_junc
rlabel poly 4639 -287 5191 -257 1 10T_4x4_magic_4/10T_toy_magic_2/WWL
rlabel locali 5118 -425 5148 -391 1 10T_4x4_magic_4/10T_toy_magic_2/RWL
rlabel locali 4682 -425 4712 -391 1 10T_4x4_magic_4/10T_toy_magic_2/RWL
rlabel locali 5103 -343 5118 -314 1 10T_4x4_magic_4/10T_toy_magic_2/WBL
rlabel locali 4713 -343 4728 -315 1 10T_4x4_magic_4/10T_toy_magic_2/WBLb
rlabel locali 5176 -489 5191 -447 1 10T_4x4_magic_4/10T_toy_magic_2/RBL0
rlabel locali 4639 -489 4654 -447 1 10T_4x4_magic_4/10T_toy_magic_2/RBL1
rlabel metal1 4899 -301 4931 -287 1 10T_4x4_magic_4/10T_toy_magic_2/VDD
rlabel metal1 4899 -527 4931 -513 7 10T_4x4_magic_4/10T_toy_magic_2/GND
rlabel polycont 4861 -420 4891 -386 1 10T_4x4_magic_4/10T_toy_magic_2/junc0
rlabel polycont 4939 -420 4969 -386 1 10T_4x4_magic_4/10T_toy_magic_2/junc1
rlabel ndiff 4712 -489 4768 -461 1 10T_4x4_magic_4/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 -489 5118 -461 1 10T_4x4_magic_4/10T_toy_magic_2/RWL0_junc
rlabel poly 5219 -17 5771 13 1 10T_4x4_magic_4/10T_toy_magic_1/WWL
rlabel locali 5698 -155 5728 -121 1 10T_4x4_magic_4/10T_toy_magic_1/RWL
rlabel locali 5262 -155 5292 -121 1 10T_4x4_magic_4/10T_toy_magic_1/RWL
rlabel locali 5683 -73 5698 -44 1 10T_4x4_magic_4/10T_toy_magic_1/WBL
rlabel locali 5293 -73 5308 -45 1 10T_4x4_magic_4/10T_toy_magic_1/WBLb
rlabel locali 5756 -219 5771 -177 1 10T_4x4_magic_4/10T_toy_magic_1/RBL0
rlabel locali 5219 -219 5234 -177 1 10T_4x4_magic_4/10T_toy_magic_1/RBL1
rlabel metal1 5479 -31 5511 -17 1 10T_4x4_magic_4/10T_toy_magic_1/VDD
rlabel metal1 5479 -257 5511 -243 7 10T_4x4_magic_4/10T_toy_magic_1/GND
rlabel polycont 5441 -150 5471 -116 1 10T_4x4_magic_4/10T_toy_magic_1/junc0
rlabel polycont 5519 -150 5549 -116 1 10T_4x4_magic_4/10T_toy_magic_1/junc1
rlabel ndiff 5292 -219 5348 -191 1 10T_4x4_magic_4/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 -219 5698 -191 1 10T_4x4_magic_4/10T_toy_magic_1/RWL0_junc
rlabel poly 4639 -17 5191 13 1 10T_4x4_magic_4/10T_toy_magic_0/WWL
rlabel locali 5118 -155 5148 -121 1 10T_4x4_magic_4/10T_toy_magic_0/RWL
rlabel locali 4682 -155 4712 -121 1 10T_4x4_magic_4/10T_toy_magic_0/RWL
rlabel locali 5103 -73 5118 -44 1 10T_4x4_magic_4/10T_toy_magic_0/WBL
rlabel locali 4713 -73 4728 -45 1 10T_4x4_magic_4/10T_toy_magic_0/WBLb
rlabel locali 5176 -219 5191 -177 1 10T_4x4_magic_4/10T_toy_magic_0/RBL0
rlabel locali 4639 -219 4654 -177 1 10T_4x4_magic_4/10T_toy_magic_0/RBL1
rlabel metal1 4899 -31 4931 -17 1 10T_4x4_magic_4/10T_toy_magic_0/VDD
rlabel metal1 4899 -257 4931 -243 7 10T_4x4_magic_4/10T_toy_magic_0/GND
rlabel polycont 4861 -150 4891 -116 1 10T_4x4_magic_4/10T_toy_magic_0/junc0
rlabel polycont 4939 -150 4969 -116 1 10T_4x4_magic_4/10T_toy_magic_0/junc1
rlabel ndiff 4712 -219 4768 -191 1 10T_4x4_magic_4/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 -219 5118 -191 1 10T_4x4_magic_4/10T_toy_magic_0/RWL0_junc
rlabel poly 4591 -557 4621 -527 1 10T_4x4_magic_5/WWL_0
rlabel poly 4591 -827 4621 -797 1 10T_4x4_magic_5/WWL_1
rlabel metal1 4591 -571 4621 -557 1 10T_4x4_magic_5/VDD
rlabel metal1 4591 -841 4621 -827 1 10T_4x4_magic_5/VDD
rlabel metal1 4591 -797 4621 -783 1 10T_4x4_magic_5/GND
rlabel metal1 4591 -1067 4621 -1053 1 10T_4x4_magic_5/GND
rlabel corelocali 4639 -1115 4654 -1085 1 10T_4x4_magic_5/RBL1_0
rlabel corelocali 5176 -1115 5191 -1085 1 10T_4x4_magic_5/RBL0_0
rlabel corelocali 5219 -1115 5234 -1085 1 10T_4x4_magic_5/RBL1_1
rlabel corelocali 5756 -1115 5771 -1085 1 10T_4x4_magic_5/RBL0_1
rlabel metal1 4591 -965 4621 -931 1 10T_4x4_magic_5/RWL_1
rlabel metal1 4591 -695 4621 -661 1 10T_4x4_magic_5/RWL_0
rlabel poly 5219 -827 5771 -797 1 10T_4x4_magic_5/10T_toy_magic_3/WWL
rlabel locali 5698 -965 5728 -931 1 10T_4x4_magic_5/10T_toy_magic_3/RWL
rlabel locali 5262 -965 5292 -931 1 10T_4x4_magic_5/10T_toy_magic_3/RWL
rlabel locali 5683 -883 5698 -854 1 10T_4x4_magic_5/10T_toy_magic_3/WBL
rlabel locali 5293 -883 5308 -855 1 10T_4x4_magic_5/10T_toy_magic_3/WBLb
rlabel locali 5756 -1029 5771 -987 1 10T_4x4_magic_5/10T_toy_magic_3/RBL0
rlabel locali 5219 -1029 5234 -987 1 10T_4x4_magic_5/10T_toy_magic_3/RBL1
rlabel metal1 5479 -841 5511 -827 1 10T_4x4_magic_5/10T_toy_magic_3/VDD
rlabel metal1 5479 -1067 5511 -1053 7 10T_4x4_magic_5/10T_toy_magic_3/GND
rlabel polycont 5441 -960 5471 -926 1 10T_4x4_magic_5/10T_toy_magic_3/junc0
rlabel polycont 5519 -960 5549 -926 1 10T_4x4_magic_5/10T_toy_magic_3/junc1
rlabel ndiff 5292 -1029 5348 -1001 1 10T_4x4_magic_5/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 -1029 5698 -1001 1 10T_4x4_magic_5/10T_toy_magic_3/RWL0_junc
rlabel poly 4639 -827 5191 -797 1 10T_4x4_magic_5/10T_toy_magic_2/WWL
rlabel locali 5118 -965 5148 -931 1 10T_4x4_magic_5/10T_toy_magic_2/RWL
rlabel locali 4682 -965 4712 -931 1 10T_4x4_magic_5/10T_toy_magic_2/RWL
rlabel locali 5103 -883 5118 -854 1 10T_4x4_magic_5/10T_toy_magic_2/WBL
rlabel locali 4713 -883 4728 -855 1 10T_4x4_magic_5/10T_toy_magic_2/WBLb
rlabel locali 5176 -1029 5191 -987 1 10T_4x4_magic_5/10T_toy_magic_2/RBL0
rlabel locali 4639 -1029 4654 -987 1 10T_4x4_magic_5/10T_toy_magic_2/RBL1
rlabel metal1 4899 -841 4931 -827 1 10T_4x4_magic_5/10T_toy_magic_2/VDD
rlabel metal1 4899 -1067 4931 -1053 7 10T_4x4_magic_5/10T_toy_magic_2/GND
rlabel polycont 4861 -960 4891 -926 1 10T_4x4_magic_5/10T_toy_magic_2/junc0
rlabel polycont 4939 -960 4969 -926 1 10T_4x4_magic_5/10T_toy_magic_2/junc1
rlabel ndiff 4712 -1029 4768 -1001 1 10T_4x4_magic_5/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 -1029 5118 -1001 1 10T_4x4_magic_5/10T_toy_magic_2/RWL0_junc
rlabel poly 5219 -557 5771 -527 1 10T_4x4_magic_5/10T_toy_magic_1/WWL
rlabel locali 5698 -695 5728 -661 1 10T_4x4_magic_5/10T_toy_magic_1/RWL
rlabel locali 5262 -695 5292 -661 1 10T_4x4_magic_5/10T_toy_magic_1/RWL
rlabel locali 5683 -613 5698 -584 1 10T_4x4_magic_5/10T_toy_magic_1/WBL
rlabel locali 5293 -613 5308 -585 1 10T_4x4_magic_5/10T_toy_magic_1/WBLb
rlabel locali 5756 -759 5771 -717 1 10T_4x4_magic_5/10T_toy_magic_1/RBL0
rlabel locali 5219 -759 5234 -717 1 10T_4x4_magic_5/10T_toy_magic_1/RBL1
rlabel metal1 5479 -571 5511 -557 1 10T_4x4_magic_5/10T_toy_magic_1/VDD
rlabel metal1 5479 -797 5511 -783 7 10T_4x4_magic_5/10T_toy_magic_1/GND
rlabel polycont 5441 -690 5471 -656 1 10T_4x4_magic_5/10T_toy_magic_1/junc0
rlabel polycont 5519 -690 5549 -656 1 10T_4x4_magic_5/10T_toy_magic_1/junc1
rlabel ndiff 5292 -759 5348 -731 1 10T_4x4_magic_5/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 -759 5698 -731 1 10T_4x4_magic_5/10T_toy_magic_1/RWL0_junc
rlabel poly 4639 -557 5191 -527 1 10T_4x4_magic_5/10T_toy_magic_0/WWL
rlabel locali 5118 -695 5148 -661 1 10T_4x4_magic_5/10T_toy_magic_0/RWL
rlabel locali 4682 -695 4712 -661 1 10T_4x4_magic_5/10T_toy_magic_0/RWL
rlabel locali 5103 -613 5118 -584 1 10T_4x4_magic_5/10T_toy_magic_0/WBL
rlabel locali 4713 -613 4728 -585 1 10T_4x4_magic_5/10T_toy_magic_0/WBLb
rlabel locali 5176 -759 5191 -717 1 10T_4x4_magic_5/10T_toy_magic_0/RBL0
rlabel locali 4639 -759 4654 -717 1 10T_4x4_magic_5/10T_toy_magic_0/RBL1
rlabel metal1 4899 -571 4931 -557 1 10T_4x4_magic_5/10T_toy_magic_0/VDD
rlabel metal1 4899 -797 4931 -783 7 10T_4x4_magic_5/10T_toy_magic_0/GND
rlabel polycont 4861 -690 4891 -656 1 10T_4x4_magic_5/10T_toy_magic_0/junc0
rlabel polycont 4939 -690 4969 -656 1 10T_4x4_magic_5/10T_toy_magic_0/junc1
rlabel ndiff 4712 -759 4768 -731 1 10T_4x4_magic_5/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 -759 5118 -731 1 10T_4x4_magic_5/10T_toy_magic_0/RWL0_junc
rlabel poly 4591 -1097 4621 -1067 1 10T_4x4_magic_6/WWL_0
rlabel poly 4591 -1367 4621 -1337 1 10T_4x4_magic_6/WWL_1
rlabel metal1 4591 -1111 4621 -1097 1 10T_4x4_magic_6/VDD
rlabel metal1 4591 -1381 4621 -1367 1 10T_4x4_magic_6/VDD
rlabel metal1 4591 -1337 4621 -1323 1 10T_4x4_magic_6/GND
rlabel metal1 4591 -1607 4621 -1593 1 10T_4x4_magic_6/GND
rlabel corelocali 4639 -1655 4654 -1625 1 10T_4x4_magic_6/RBL1_0
rlabel corelocali 5176 -1655 5191 -1625 1 10T_4x4_magic_6/RBL0_0
rlabel corelocali 5219 -1655 5234 -1625 1 10T_4x4_magic_6/RBL1_1
rlabel corelocali 5756 -1655 5771 -1625 1 10T_4x4_magic_6/RBL0_1
rlabel metal1 4591 -1505 4621 -1471 1 10T_4x4_magic_6/RWL_1
rlabel metal1 4591 -1235 4621 -1201 1 10T_4x4_magic_6/RWL_0
rlabel poly 5219 -1367 5771 -1337 1 10T_4x4_magic_6/10T_toy_magic_3/WWL
rlabel locali 5698 -1505 5728 -1471 1 10T_4x4_magic_6/10T_toy_magic_3/RWL
rlabel locali 5262 -1505 5292 -1471 1 10T_4x4_magic_6/10T_toy_magic_3/RWL
rlabel locali 5683 -1423 5698 -1394 1 10T_4x4_magic_6/10T_toy_magic_3/WBL
rlabel locali 5293 -1423 5308 -1395 1 10T_4x4_magic_6/10T_toy_magic_3/WBLb
rlabel locali 5756 -1569 5771 -1527 1 10T_4x4_magic_6/10T_toy_magic_3/RBL0
rlabel locali 5219 -1569 5234 -1527 1 10T_4x4_magic_6/10T_toy_magic_3/RBL1
rlabel metal1 5479 -1381 5511 -1367 1 10T_4x4_magic_6/10T_toy_magic_3/VDD
rlabel metal1 5479 -1607 5511 -1593 7 10T_4x4_magic_6/10T_toy_magic_3/GND
rlabel polycont 5441 -1500 5471 -1466 1 10T_4x4_magic_6/10T_toy_magic_3/junc0
rlabel polycont 5519 -1500 5549 -1466 1 10T_4x4_magic_6/10T_toy_magic_3/junc1
rlabel ndiff 5292 -1569 5348 -1541 1 10T_4x4_magic_6/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 -1569 5698 -1541 1 10T_4x4_magic_6/10T_toy_magic_3/RWL0_junc
rlabel poly 4639 -1367 5191 -1337 1 10T_4x4_magic_6/10T_toy_magic_2/WWL
rlabel locali 5118 -1505 5148 -1471 1 10T_4x4_magic_6/10T_toy_magic_2/RWL
rlabel locali 4682 -1505 4712 -1471 1 10T_4x4_magic_6/10T_toy_magic_2/RWL
rlabel locali 5103 -1423 5118 -1394 1 10T_4x4_magic_6/10T_toy_magic_2/WBL
rlabel locali 4713 -1423 4728 -1395 1 10T_4x4_magic_6/10T_toy_magic_2/WBLb
rlabel locali 5176 -1569 5191 -1527 1 10T_4x4_magic_6/10T_toy_magic_2/RBL0
rlabel locali 4639 -1569 4654 -1527 1 10T_4x4_magic_6/10T_toy_magic_2/RBL1
rlabel metal1 4899 -1381 4931 -1367 1 10T_4x4_magic_6/10T_toy_magic_2/VDD
rlabel metal1 4899 -1607 4931 -1593 7 10T_4x4_magic_6/10T_toy_magic_2/GND
rlabel polycont 4861 -1500 4891 -1466 1 10T_4x4_magic_6/10T_toy_magic_2/junc0
rlabel polycont 4939 -1500 4969 -1466 1 10T_4x4_magic_6/10T_toy_magic_2/junc1
rlabel ndiff 4712 -1569 4768 -1541 1 10T_4x4_magic_6/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 -1569 5118 -1541 1 10T_4x4_magic_6/10T_toy_magic_2/RWL0_junc
rlabel poly 5219 -1097 5771 -1067 1 10T_4x4_magic_6/10T_toy_magic_1/WWL
rlabel locali 5698 -1235 5728 -1201 1 10T_4x4_magic_6/10T_toy_magic_1/RWL
rlabel locali 5262 -1235 5292 -1201 1 10T_4x4_magic_6/10T_toy_magic_1/RWL
rlabel locali 5683 -1153 5698 -1124 1 10T_4x4_magic_6/10T_toy_magic_1/WBL
rlabel locali 5293 -1153 5308 -1125 1 10T_4x4_magic_6/10T_toy_magic_1/WBLb
rlabel locali 5756 -1299 5771 -1257 1 10T_4x4_magic_6/10T_toy_magic_1/RBL0
rlabel locali 5219 -1299 5234 -1257 1 10T_4x4_magic_6/10T_toy_magic_1/RBL1
rlabel metal1 5479 -1111 5511 -1097 1 10T_4x4_magic_6/10T_toy_magic_1/VDD
rlabel metal1 5479 -1337 5511 -1323 7 10T_4x4_magic_6/10T_toy_magic_1/GND
rlabel polycont 5441 -1230 5471 -1196 1 10T_4x4_magic_6/10T_toy_magic_1/junc0
rlabel polycont 5519 -1230 5549 -1196 1 10T_4x4_magic_6/10T_toy_magic_1/junc1
rlabel ndiff 5292 -1299 5348 -1271 1 10T_4x4_magic_6/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 -1299 5698 -1271 1 10T_4x4_magic_6/10T_toy_magic_1/RWL0_junc
rlabel poly 4639 -1097 5191 -1067 1 10T_4x4_magic_6/10T_toy_magic_0/WWL
rlabel locali 5118 -1235 5148 -1201 1 10T_4x4_magic_6/10T_toy_magic_0/RWL
rlabel locali 4682 -1235 4712 -1201 1 10T_4x4_magic_6/10T_toy_magic_0/RWL
rlabel locali 5103 -1153 5118 -1124 1 10T_4x4_magic_6/10T_toy_magic_0/WBL
rlabel locali 4713 -1153 4728 -1125 1 10T_4x4_magic_6/10T_toy_magic_0/WBLb
rlabel locali 5176 -1299 5191 -1257 1 10T_4x4_magic_6/10T_toy_magic_0/RBL0
rlabel locali 4639 -1299 4654 -1257 1 10T_4x4_magic_6/10T_toy_magic_0/RBL1
rlabel metal1 4899 -1111 4931 -1097 1 10T_4x4_magic_6/10T_toy_magic_0/VDD
rlabel metal1 4899 -1337 4931 -1323 7 10T_4x4_magic_6/10T_toy_magic_0/GND
rlabel polycont 4861 -1230 4891 -1196 1 10T_4x4_magic_6/10T_toy_magic_0/junc0
rlabel polycont 4939 -1230 4969 -1196 1 10T_4x4_magic_6/10T_toy_magic_0/junc1
rlabel ndiff 4712 -1299 4768 -1271 1 10T_4x4_magic_6/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 -1299 5118 -1271 1 10T_4x4_magic_6/10T_toy_magic_0/RWL0_junc
rlabel poly 4591 -1637 4621 -1607 1 10T_4x4_magic_7/WWL_0
rlabel poly 4591 -1907 4621 -1877 1 10T_4x4_magic_7/WWL_1
rlabel metal1 4591 -1651 4621 -1637 1 10T_4x4_magic_7/VDD
rlabel metal1 4591 -1921 4621 -1907 1 10T_4x4_magic_7/VDD
rlabel metal1 4591 -1877 4621 -1863 1 10T_4x4_magic_7/GND
rlabel metal1 4591 -2147 4621 -2133 1 10T_4x4_magic_7/GND
rlabel metal1 4591 -2045 4621 -2011 1 10T_4x4_magic_7/RWL_1
rlabel metal1 4591 -1775 4621 -1741 1 10T_4x4_magic_7/RWL_0
rlabel poly 5219 -1907 5771 -1877 1 10T_4x4_magic_7/10T_toy_magic_3/WWL
rlabel locali 5698 -2045 5728 -2011 1 10T_4x4_magic_7/10T_toy_magic_3/RWL
rlabel locali 5262 -2045 5292 -2011 1 10T_4x4_magic_7/10T_toy_magic_3/RWL
rlabel locali 5683 -1963 5698 -1934 1 10T_4x4_magic_7/10T_toy_magic_3/WBL
rlabel locali 5293 -1963 5308 -1935 1 10T_4x4_magic_7/10T_toy_magic_3/WBLb
rlabel locali 5756 -2109 5771 -2067 1 10T_4x4_magic_7/10T_toy_magic_3/RBL0
rlabel locali 5219 -2109 5234 -2067 1 10T_4x4_magic_7/10T_toy_magic_3/RBL1
rlabel metal1 5479 -1921 5511 -1907 1 10T_4x4_magic_7/10T_toy_magic_3/VDD
rlabel metal1 5479 -2147 5511 -2133 7 10T_4x4_magic_7/10T_toy_magic_3/GND
rlabel polycont 5441 -2040 5471 -2006 1 10T_4x4_magic_7/10T_toy_magic_3/junc0
rlabel polycont 5519 -2040 5549 -2006 1 10T_4x4_magic_7/10T_toy_magic_3/junc1
rlabel ndiff 5292 -2109 5348 -2081 1 10T_4x4_magic_7/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 -2109 5698 -2081 1 10T_4x4_magic_7/10T_toy_magic_3/RWL0_junc
rlabel poly 4639 -1907 5191 -1877 1 10T_4x4_magic_7/10T_toy_magic_2/WWL
rlabel locali 5118 -2045 5148 -2011 1 10T_4x4_magic_7/10T_toy_magic_2/RWL
rlabel locali 4682 -2045 4712 -2011 1 10T_4x4_magic_7/10T_toy_magic_2/RWL
rlabel locali 5103 -1963 5118 -1934 1 10T_4x4_magic_7/10T_toy_magic_2/WBL
rlabel locali 4713 -1963 4728 -1935 1 10T_4x4_magic_7/10T_toy_magic_2/WBLb
rlabel locali 5176 -2109 5191 -2067 1 10T_4x4_magic_7/10T_toy_magic_2/RBL0
rlabel locali 4639 -2109 4654 -2067 1 10T_4x4_magic_7/10T_toy_magic_2/RBL1
rlabel metal1 4899 -1921 4931 -1907 1 10T_4x4_magic_7/10T_toy_magic_2/VDD
rlabel metal1 4899 -2147 4931 -2133 7 10T_4x4_magic_7/10T_toy_magic_2/GND
rlabel polycont 4861 -2040 4891 -2006 1 10T_4x4_magic_7/10T_toy_magic_2/junc0
rlabel polycont 4939 -2040 4969 -2006 1 10T_4x4_magic_7/10T_toy_magic_2/junc1
rlabel ndiff 4712 -2109 4768 -2081 1 10T_4x4_magic_7/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 -2109 5118 -2081 1 10T_4x4_magic_7/10T_toy_magic_2/RWL0_junc
rlabel poly 5219 -1637 5771 -1607 1 10T_4x4_magic_7/10T_toy_magic_1/WWL
rlabel locali 5698 -1775 5728 -1741 1 10T_4x4_magic_7/10T_toy_magic_1/RWL
rlabel locali 5262 -1775 5292 -1741 1 10T_4x4_magic_7/10T_toy_magic_1/RWL
rlabel locali 5683 -1693 5698 -1664 1 10T_4x4_magic_7/10T_toy_magic_1/WBL
rlabel locali 5293 -1693 5308 -1665 1 10T_4x4_magic_7/10T_toy_magic_1/WBLb
rlabel locali 5756 -1839 5771 -1797 1 10T_4x4_magic_7/10T_toy_magic_1/RBL0
rlabel locali 5219 -1839 5234 -1797 1 10T_4x4_magic_7/10T_toy_magic_1/RBL1
rlabel metal1 5479 -1651 5511 -1637 1 10T_4x4_magic_7/10T_toy_magic_1/VDD
rlabel metal1 5479 -1877 5511 -1863 7 10T_4x4_magic_7/10T_toy_magic_1/GND
rlabel polycont 5441 -1770 5471 -1736 1 10T_4x4_magic_7/10T_toy_magic_1/junc0
rlabel polycont 5519 -1770 5549 -1736 1 10T_4x4_magic_7/10T_toy_magic_1/junc1
rlabel ndiff 5292 -1839 5348 -1811 1 10T_4x4_magic_7/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 -1839 5698 -1811 1 10T_4x4_magic_7/10T_toy_magic_1/RWL0_junc
rlabel poly 4639 -1637 5191 -1607 1 10T_4x4_magic_7/10T_toy_magic_0/WWL
rlabel locali 5118 -1775 5148 -1741 1 10T_4x4_magic_7/10T_toy_magic_0/RWL
rlabel locali 4682 -1775 4712 -1741 1 10T_4x4_magic_7/10T_toy_magic_0/RWL
rlabel locali 5103 -1693 5118 -1664 1 10T_4x4_magic_7/10T_toy_magic_0/WBL
rlabel locali 4713 -1693 4728 -1665 1 10T_4x4_magic_7/10T_toy_magic_0/WBLb
rlabel locali 5176 -1839 5191 -1797 1 10T_4x4_magic_7/10T_toy_magic_0/RBL0
rlabel locali 4639 -1839 4654 -1797 1 10T_4x4_magic_7/10T_toy_magic_0/RBL1
rlabel metal1 4899 -1651 4931 -1637 1 10T_4x4_magic_7/10T_toy_magic_0/VDD
rlabel metal1 4899 -1877 4931 -1863 7 10T_4x4_magic_7/10T_toy_magic_0/GND
rlabel polycont 4861 -1770 4891 -1736 1 10T_4x4_magic_7/10T_toy_magic_0/junc0
rlabel polycont 4939 -1770 4969 -1736 1 10T_4x4_magic_7/10T_toy_magic_0/junc1
rlabel ndiff 4712 -1839 4768 -1811 1 10T_4x4_magic_7/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 -1839 5118 -1811 1 10T_4x4_magic_7/10T_toy_magic_0/RWL0_junc
rlabel locali -1 52 14 94 1 10T_8x8_magic_0/RBL1_0
rlabel locali 536 52 551 94 1 10T_8x8_magic_0/RBL0_0
rlabel locali 579 52 594 94 1 10T_8x8_magic_0/RBL1_1
rlabel locali 1116 52 1131 94 1 10T_8x8_magic_0/RBL0_1
rlabel locali 1159 52 1174 94 1 10T_8x8_magic_0/RBL1_2
rlabel locali 1696 52 1711 94 1 10T_8x8_magic_0/RBL0_2
rlabel locali 1739 52 1754 94 1 10T_8x8_magic_0/RBL1_3
rlabel locali 2276 52 2291 94 1 10T_8x8_magic_0/RBL0_3
rlabel locali 2319 52 2334 94 1 10T_8x8_magic_0/RBL1_4
rlabel locali 2856 52 2871 94 1 10T_8x8_magic_0/RBL0_4
rlabel locali 2899 52 2914 94 1 10T_8x8_magic_0/RBL1_5
rlabel locali 3436 52 3451 94 1 10T_8x8_magic_0/RBL0_5
rlabel locali 3479 52 3494 94 1 10T_8x8_magic_0/RBL1_6
rlabel locali 4016 52 4031 94 1 10T_8x8_magic_0/RBL0_6
rlabel locali 4059 52 4074 94 1 10T_8x8_magic_0/RBL1_7
rlabel locali 4596 52 4611 94 1 10T_8x8_magic_0/RBL0_7
rlabel locali 463 198 478 227 1 10T_8x8_magic_0/WBL_0
rlabel locali 73 198 88 226 1 10T_8x8_magic_0/WBLb_0
rlabel locali 1043 198 1058 227 1 10T_8x8_magic_0/WBL_1
rlabel locali 653 198 668 226 1 10T_8x8_magic_0/WBLb_1
rlabel locali 1623 198 1638 227 1 10T_8x8_magic_0/WBL_2
rlabel locali 1233 198 1248 226 1 10T_8x8_magic_0/WBLb_2
rlabel locali 2203 198 2218 227 1 10T_8x8_magic_0/WBL_3
rlabel locali 1813 198 1828 226 1 10T_8x8_magic_0/WBLb_3
rlabel locali 2783 198 2798 227 1 10T_8x8_magic_0/WBL_4
rlabel locali 2393 198 2408 226 1 10T_8x8_magic_0/WBLb_4
rlabel locali 3363 198 3378 227 1 10T_8x8_magic_0/WBL_5
rlabel locali 2973 198 2988 226 1 10T_8x8_magic_0/WBLb_5
rlabel locali 3943 198 3958 227 1 10T_8x8_magic_0/WBL_6
rlabel locali 3553 198 3568 226 1 10T_8x8_magic_0/WBLb_6
rlabel locali 4523 198 4538 227 1 10T_8x8_magic_0/WBL_7
rlabel locali 4133 198 4148 226 1 10T_8x8_magic_0/WBLb_7
rlabel metal1 -1 1736 14 1770 1 10T_8x8_magic_0/RWL_1
rlabel metal1 -1 1466 14 1500 1 10T_8x8_magic_0/RWL_2
rlabel metal1 -1 1196 14 1230 1 10T_8x8_magic_0/RWL_3
rlabel metal1 -1 926 14 960 1 10T_8x8_magic_0/RWL_4
rlabel metal1 -1 656 14 690 1 10T_8x8_magic_0/RWL_5
rlabel poly -1 524 29 554 1 10T_8x8_magic_0/WWL_6
rlabel metal1 -1 386 14 420 1 10T_8x8_magic_0/RWL_6
rlabel poly -1 254 29 284 1 10T_8x8_magic_0/WWL_7
rlabel metal1 -1 116 14 150 1 10T_8x8_magic_0/RWL_7
rlabel metal1 -1 1590 14 1604 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 1320 14 1334 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 1860 14 1874 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 1050 14 1064 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 510 14 524 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 240 14 254 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 780 14 794 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 1094 14 1108 1 10T_8x8_magic_0/GND
rlabel metal1 -1 1364 14 1378 1 10T_8x8_magic_0/GND
rlabel metal1 -1 1634 14 1648 1 10T_8x8_magic_0/GND
rlabel metal1 -1 824 14 838 1 10T_8x8_magic_0/GND
rlabel metal1 -1 14 14 28 1 10T_8x8_magic_0/GND
rlabel metal1 -1 284 14 298 1 10T_8x8_magic_0/GND
rlabel metal1 -1 554 14 568 1 10T_8x8_magic_0/GND
rlabel metal1 -1 656 14 690 1 10T_8x8_magic_0/10T_1x8_magic_7/RWL
rlabel corelocali 73 738 88 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_0
rlabel corelocali 463 738 478 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_0
rlabel corelocali -1 592 14 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_0
rlabel corelocali 536 592 551 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_0
rlabel corelocali 653 738 668 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_1
rlabel corelocali 1043 738 1058 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_1
rlabel corelocali 579 592 594 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_1
rlabel corelocali 1116 592 1131 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_1
rlabel corelocali 1233 738 1248 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_2
rlabel corelocali 1623 738 1638 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_2
rlabel corelocali 1159 592 1174 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_2
rlabel corelocali 1696 592 1711 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_2
rlabel corelocali 1813 738 1828 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_3
rlabel corelocali 2203 738 2218 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_3
rlabel corelocali 1739 592 1754 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_3
rlabel corelocali 2276 592 2291 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_3
rlabel corelocali 2393 738 2408 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_4
rlabel corelocali 2783 738 2798 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_4
rlabel corelocali 2319 592 2334 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_4
rlabel corelocali 2856 592 2871 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_4
rlabel corelocali 2973 738 2988 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_5
rlabel corelocali 3363 738 3378 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_5
rlabel corelocali 2899 592 2914 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_5
rlabel corelocali 3436 592 3451 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_5
rlabel corelocali 3553 738 3568 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_6
rlabel corelocali 3943 738 3958 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_6
rlabel corelocali 3479 592 3494 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_6
rlabel corelocali 4016 592 4031 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_6
rlabel corelocali 4133 738 4148 766 1 10T_8x8_magic_0/10T_1x8_magic_7/WBLb_7
rlabel corelocali 4523 738 4538 767 1 10T_8x8_magic_0/10T_1x8_magic_7/WBL_7
rlabel corelocali 4059 592 4074 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL1_7
rlabel corelocali 4596 592 4611 634 1 10T_8x8_magic_0/10T_1x8_magic_7/RBL0_7
rlabel metal1 -1 780 14 794 1 10T_8x8_magic_0/10T_1x8_magic_7/VDD
rlabel metal1 -1 554 14 568 1 10T_8x8_magic_0/10T_1x8_magic_7/GND
rlabel locali 478 656 508 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/RWL
rlabel locali 42 656 72 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/RWL
rlabel locali 463 738 478 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/WBL
rlabel locali 73 738 88 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/WBLb
rlabel locali 536 592 551 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/RBL0
rlabel locali -1 592 14 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/RBL1
rlabel metal1 259 780 291 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/VDD
rlabel metal1 259 554 291 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/GND
rlabel polycont 221 661 251 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/junc0
rlabel polycont 299 661 329 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/junc1
rlabel ndiff 72 592 128 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 592 478 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_7/RWL0_junc
rlabel locali 1058 656 1088 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/RWL
rlabel locali 622 656 652 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/RWL
rlabel locali 1043 738 1058 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/WBL
rlabel locali 653 738 668 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/WBLb
rlabel locali 1116 592 1131 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/RBL0
rlabel locali 579 592 594 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/RBL1
rlabel metal1 839 780 871 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/VDD
rlabel metal1 839 554 871 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/GND
rlabel polycont 801 661 831 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/junc0
rlabel polycont 879 661 909 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/junc1
rlabel ndiff 652 592 708 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 592 1058 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_6/RWL0_junc
rlabel locali 1638 656 1668 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/RWL
rlabel locali 1202 656 1232 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/RWL
rlabel locali 1623 738 1638 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/WBL
rlabel locali 1233 738 1248 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/WBLb
rlabel locali 1696 592 1711 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/RBL0
rlabel locali 1159 592 1174 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/RBL1
rlabel metal1 1419 780 1451 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/VDD
rlabel metal1 1419 554 1451 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/GND
rlabel polycont 1381 661 1411 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/junc0
rlabel polycont 1459 661 1489 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/junc1
rlabel ndiff 1232 592 1288 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 592 1638 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_5/RWL0_junc
rlabel locali 2218 656 2248 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/RWL
rlabel locali 1782 656 1812 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/RWL
rlabel locali 2203 738 2218 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/WBL
rlabel locali 1813 738 1828 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/WBLb
rlabel locali 2276 592 2291 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/RBL0
rlabel locali 1739 592 1754 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/RBL1
rlabel metal1 1999 780 2031 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/VDD
rlabel metal1 1999 554 2031 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/GND
rlabel polycont 1961 661 1991 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/junc0
rlabel polycont 2039 661 2069 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/junc1
rlabel ndiff 1812 592 1868 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 592 2218 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_4/RWL0_junc
rlabel locali 2798 656 2828 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/RWL
rlabel locali 2362 656 2392 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/RWL
rlabel locali 2783 738 2798 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/WBL
rlabel locali 2393 738 2408 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/WBLb
rlabel locali 2856 592 2871 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/RBL0
rlabel locali 2319 592 2334 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/RBL1
rlabel metal1 2579 780 2611 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/VDD
rlabel metal1 2579 554 2611 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/GND
rlabel polycont 2541 661 2571 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/junc0
rlabel polycont 2619 661 2649 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/junc1
rlabel ndiff 2392 592 2448 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 592 2798 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_3/RWL0_junc
rlabel locali 3378 656 3408 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/RWL
rlabel locali 2942 656 2972 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/RWL
rlabel locali 3363 738 3378 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/WBL
rlabel locali 2973 738 2988 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/WBLb
rlabel locali 3436 592 3451 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/RBL0
rlabel locali 2899 592 2914 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/RBL1
rlabel metal1 3159 780 3191 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/VDD
rlabel metal1 3159 554 3191 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/GND
rlabel polycont 3121 661 3151 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/junc0
rlabel polycont 3199 661 3229 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/junc1
rlabel ndiff 2972 592 3028 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 592 3378 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_2/RWL0_junc
rlabel locali 4538 656 4568 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/RWL
rlabel locali 4102 656 4132 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/RWL
rlabel locali 4523 738 4538 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/WBL
rlabel locali 4133 738 4148 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/WBLb
rlabel locali 4596 592 4611 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/RBL0
rlabel locali 4059 592 4074 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/RBL1
rlabel metal1 4319 780 4351 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/VDD
rlabel metal1 4319 554 4351 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/GND
rlabel polycont 4281 661 4311 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/junc0
rlabel polycont 4359 661 4389 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/junc1
rlabel ndiff 4132 592 4188 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 592 4538 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_1/RWL0_junc
rlabel locali 3958 656 3988 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/RWL
rlabel locali 3522 656 3552 690 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/RWL
rlabel locali 3943 738 3958 767 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/WBL
rlabel locali 3553 738 3568 766 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/WBLb
rlabel locali 4016 592 4031 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/RBL0
rlabel locali 3479 592 3494 634 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/RBL1
rlabel metal1 3739 780 3771 794 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/VDD
rlabel metal1 3739 554 3771 568 7 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/GND
rlabel polycont 3701 661 3731 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/junc0
rlabel polycont 3779 661 3809 695 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/junc1
rlabel ndiff 3552 592 3608 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 592 3958 620 1 10T_8x8_magic_0/10T_1x8_magic_7/10T_toy_magic_0/RWL0_junc
rlabel metal1 -1 926 14 960 1 10T_8x8_magic_0/10T_1x8_magic_6/RWL
rlabel corelocali 73 1008 88 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_0
rlabel corelocali 463 1008 478 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_0
rlabel corelocali -1 862 14 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_0
rlabel corelocali 536 862 551 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_0
rlabel corelocali 653 1008 668 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_1
rlabel corelocali 1043 1008 1058 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_1
rlabel corelocali 579 862 594 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_1
rlabel corelocali 1116 862 1131 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_1
rlabel corelocali 1233 1008 1248 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_2
rlabel corelocali 1623 1008 1638 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_2
rlabel corelocali 1159 862 1174 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_2
rlabel corelocali 1696 862 1711 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_2
rlabel corelocali 1813 1008 1828 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_3
rlabel corelocali 2203 1008 2218 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_3
rlabel corelocali 1739 862 1754 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_3
rlabel corelocali 2276 862 2291 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_3
rlabel corelocali 2393 1008 2408 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_4
rlabel corelocali 2783 1008 2798 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_4
rlabel corelocali 2319 862 2334 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_4
rlabel corelocali 2856 862 2871 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_4
rlabel corelocali 2973 1008 2988 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_5
rlabel corelocali 3363 1008 3378 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_5
rlabel corelocali 2899 862 2914 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_5
rlabel corelocali 3436 862 3451 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_5
rlabel corelocali 3553 1008 3568 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_6
rlabel corelocali 3943 1008 3958 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_6
rlabel corelocali 3479 862 3494 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_6
rlabel corelocali 4016 862 4031 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_6
rlabel corelocali 4133 1008 4148 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/WBLb_7
rlabel corelocali 4523 1008 4538 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/WBL_7
rlabel corelocali 4059 862 4074 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL1_7
rlabel corelocali 4596 862 4611 904 1 10T_8x8_magic_0/10T_1x8_magic_6/RBL0_7
rlabel metal1 -1 1050 14 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/VDD
rlabel metal1 -1 824 14 838 1 10T_8x8_magic_0/10T_1x8_magic_6/GND
rlabel locali 478 926 508 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/RWL
rlabel locali 42 926 72 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/RWL
rlabel locali 463 1008 478 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/WBL
rlabel locali 73 1008 88 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/WBLb
rlabel locali 536 862 551 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/RBL0
rlabel locali -1 862 14 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/RBL1
rlabel metal1 259 1050 291 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/VDD
rlabel metal1 259 824 291 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/GND
rlabel polycont 221 931 251 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/junc0
rlabel polycont 299 931 329 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/junc1
rlabel ndiff 72 862 128 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 862 478 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_7/RWL0_junc
rlabel locali 1058 926 1088 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/RWL
rlabel locali 622 926 652 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/RWL
rlabel locali 1043 1008 1058 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/WBL
rlabel locali 653 1008 668 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/WBLb
rlabel locali 1116 862 1131 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/RBL0
rlabel locali 579 862 594 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/RBL1
rlabel metal1 839 1050 871 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/VDD
rlabel metal1 839 824 871 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/GND
rlabel polycont 801 931 831 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/junc0
rlabel polycont 879 931 909 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/junc1
rlabel ndiff 652 862 708 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 862 1058 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_6/RWL0_junc
rlabel locali 1638 926 1668 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/RWL
rlabel locali 1202 926 1232 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/RWL
rlabel locali 1623 1008 1638 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/WBL
rlabel locali 1233 1008 1248 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/WBLb
rlabel locali 1696 862 1711 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/RBL0
rlabel locali 1159 862 1174 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/RBL1
rlabel metal1 1419 1050 1451 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/VDD
rlabel metal1 1419 824 1451 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/GND
rlabel polycont 1381 931 1411 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/junc0
rlabel polycont 1459 931 1489 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/junc1
rlabel ndiff 1232 862 1288 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 862 1638 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_5/RWL0_junc
rlabel locali 2218 926 2248 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/RWL
rlabel locali 1782 926 1812 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/RWL
rlabel locali 2203 1008 2218 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/WBL
rlabel locali 1813 1008 1828 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/WBLb
rlabel locali 2276 862 2291 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/RBL0
rlabel locali 1739 862 1754 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/RBL1
rlabel metal1 1999 1050 2031 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/VDD
rlabel metal1 1999 824 2031 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/GND
rlabel polycont 1961 931 1991 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/junc0
rlabel polycont 2039 931 2069 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/junc1
rlabel ndiff 1812 862 1868 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 862 2218 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_4/RWL0_junc
rlabel locali 2798 926 2828 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/RWL
rlabel locali 2362 926 2392 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/RWL
rlabel locali 2783 1008 2798 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/WBL
rlabel locali 2393 1008 2408 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/WBLb
rlabel locali 2856 862 2871 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/RBL0
rlabel locali 2319 862 2334 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/RBL1
rlabel metal1 2579 1050 2611 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/VDD
rlabel metal1 2579 824 2611 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/GND
rlabel polycont 2541 931 2571 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/junc0
rlabel polycont 2619 931 2649 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/junc1
rlabel ndiff 2392 862 2448 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 862 2798 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_3/RWL0_junc
rlabel locali 3378 926 3408 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/RWL
rlabel locali 2942 926 2972 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/RWL
rlabel locali 3363 1008 3378 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/WBL
rlabel locali 2973 1008 2988 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/WBLb
rlabel locali 3436 862 3451 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/RBL0
rlabel locali 2899 862 2914 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/RBL1
rlabel metal1 3159 1050 3191 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/VDD
rlabel metal1 3159 824 3191 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/GND
rlabel polycont 3121 931 3151 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/junc0
rlabel polycont 3199 931 3229 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/junc1
rlabel ndiff 2972 862 3028 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 862 3378 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_2/RWL0_junc
rlabel locali 4538 926 4568 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/RWL
rlabel locali 4102 926 4132 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/RWL
rlabel locali 4523 1008 4538 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/WBL
rlabel locali 4133 1008 4148 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/WBLb
rlabel locali 4596 862 4611 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/RBL0
rlabel locali 4059 862 4074 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/RBL1
rlabel metal1 4319 1050 4351 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/VDD
rlabel metal1 4319 824 4351 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/GND
rlabel polycont 4281 931 4311 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/junc0
rlabel polycont 4359 931 4389 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/junc1
rlabel ndiff 4132 862 4188 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 862 4538 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_1/RWL0_junc
rlabel locali 3958 926 3988 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/RWL
rlabel locali 3522 926 3552 960 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/RWL
rlabel locali 3943 1008 3958 1037 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/WBL
rlabel locali 3553 1008 3568 1036 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/WBLb
rlabel locali 4016 862 4031 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/RBL0
rlabel locali 3479 862 3494 904 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/RBL1
rlabel metal1 3739 1050 3771 1064 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/VDD
rlabel metal1 3739 824 3771 838 7 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/GND
rlabel polycont 3701 931 3731 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/junc0
rlabel polycont 3779 931 3809 965 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/junc1
rlabel ndiff 3552 862 3608 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 862 3958 890 1 10T_8x8_magic_0/10T_1x8_magic_6/10T_toy_magic_0/RWL0_junc
rlabel poly -1 524 29 554 1 10T_8x8_magic_0/10T_1x8_magic_5/WWL
rlabel metal1 -1 386 14 420 1 10T_8x8_magic_0/10T_1x8_magic_5/RWL
rlabel corelocali 73 468 88 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_0
rlabel corelocali 463 468 478 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_0
rlabel corelocali -1 322 14 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_0
rlabel corelocali 536 322 551 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_0
rlabel corelocali 653 468 668 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_1
rlabel corelocali 1043 468 1058 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_1
rlabel corelocali 579 322 594 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_1
rlabel corelocali 1116 322 1131 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_1
rlabel corelocali 1233 468 1248 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_2
rlabel corelocali 1623 468 1638 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_2
rlabel corelocali 1159 322 1174 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_2
rlabel corelocali 1696 322 1711 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_2
rlabel corelocali 1813 468 1828 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_3
rlabel corelocali 2203 468 2218 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_3
rlabel corelocali 1739 322 1754 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_3
rlabel corelocali 2276 322 2291 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_3
rlabel corelocali 2393 468 2408 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_4
rlabel corelocali 2783 468 2798 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_4
rlabel corelocali 2319 322 2334 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_4
rlabel corelocali 2856 322 2871 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_4
rlabel corelocali 2973 468 2988 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_5
rlabel corelocali 3363 468 3378 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_5
rlabel corelocali 2899 322 2914 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_5
rlabel corelocali 3436 322 3451 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_5
rlabel corelocali 3553 468 3568 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_6
rlabel corelocali 3943 468 3958 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_6
rlabel corelocali 3479 322 3494 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_6
rlabel corelocali 4016 322 4031 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_6
rlabel corelocali 4133 468 4148 496 1 10T_8x8_magic_0/10T_1x8_magic_5/WBLb_7
rlabel corelocali 4523 468 4538 497 1 10T_8x8_magic_0/10T_1x8_magic_5/WBL_7
rlabel corelocali 4059 322 4074 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL1_7
rlabel corelocali 4596 322 4611 364 1 10T_8x8_magic_0/10T_1x8_magic_5/RBL0_7
rlabel metal1 -1 510 14 524 1 10T_8x8_magic_0/10T_1x8_magic_5/VDD
rlabel metal1 -1 284 14 298 1 10T_8x8_magic_0/10T_1x8_magic_5/GND
rlabel poly -1 524 551 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/WWL
rlabel locali 478 386 508 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/RWL
rlabel locali 42 386 72 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/RWL
rlabel locali 463 468 478 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/WBL
rlabel locali 73 468 88 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/WBLb
rlabel locali 536 322 551 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/RBL0
rlabel locali -1 322 14 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/RBL1
rlabel metal1 259 510 291 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/VDD
rlabel metal1 259 284 291 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/GND
rlabel polycont 221 391 251 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/junc0
rlabel polycont 299 391 329 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/junc1
rlabel ndiff 72 322 128 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 322 478 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_7/RWL0_junc
rlabel poly 579 524 1131 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/WWL
rlabel locali 1058 386 1088 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/RWL
rlabel locali 622 386 652 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/RWL
rlabel locali 1043 468 1058 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/WBL
rlabel locali 653 468 668 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/WBLb
rlabel locali 1116 322 1131 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/RBL0
rlabel locali 579 322 594 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/RBL1
rlabel metal1 839 510 871 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/VDD
rlabel metal1 839 284 871 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/GND
rlabel polycont 801 391 831 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/junc0
rlabel polycont 879 391 909 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/junc1
rlabel ndiff 652 322 708 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 322 1058 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 524 1711 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/WWL
rlabel locali 1638 386 1668 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/RWL
rlabel locali 1202 386 1232 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/RWL
rlabel locali 1623 468 1638 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/WBL
rlabel locali 1233 468 1248 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/WBLb
rlabel locali 1696 322 1711 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/RBL0
rlabel locali 1159 322 1174 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/RBL1
rlabel metal1 1419 510 1451 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/VDD
rlabel metal1 1419 284 1451 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/GND
rlabel polycont 1381 391 1411 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/junc0
rlabel polycont 1459 391 1489 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/junc1
rlabel ndiff 1232 322 1288 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 322 1638 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 524 2291 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/WWL
rlabel locali 2218 386 2248 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/RWL
rlabel locali 1782 386 1812 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/RWL
rlabel locali 2203 468 2218 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/WBL
rlabel locali 1813 468 1828 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/WBLb
rlabel locali 2276 322 2291 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/RBL0
rlabel locali 1739 322 1754 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/RBL1
rlabel metal1 1999 510 2031 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/VDD
rlabel metal1 1999 284 2031 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/GND
rlabel polycont 1961 391 1991 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/junc0
rlabel polycont 2039 391 2069 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/junc1
rlabel ndiff 1812 322 1868 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 322 2218 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 524 2871 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/WWL
rlabel locali 2798 386 2828 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/RWL
rlabel locali 2362 386 2392 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/RWL
rlabel locali 2783 468 2798 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/WBL
rlabel locali 2393 468 2408 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/WBLb
rlabel locali 2856 322 2871 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/RBL0
rlabel locali 2319 322 2334 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/RBL1
rlabel metal1 2579 510 2611 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/VDD
rlabel metal1 2579 284 2611 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/GND
rlabel polycont 2541 391 2571 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/junc0
rlabel polycont 2619 391 2649 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/junc1
rlabel ndiff 2392 322 2448 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 322 2798 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 524 3451 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/WWL
rlabel locali 3378 386 3408 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/RWL
rlabel locali 2942 386 2972 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/RWL
rlabel locali 3363 468 3378 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/WBL
rlabel locali 2973 468 2988 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/WBLb
rlabel locali 3436 322 3451 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/RBL0
rlabel locali 2899 322 2914 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/RBL1
rlabel metal1 3159 510 3191 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/VDD
rlabel metal1 3159 284 3191 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/GND
rlabel polycont 3121 391 3151 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/junc0
rlabel polycont 3199 391 3229 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/junc1
rlabel ndiff 2972 322 3028 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 322 3378 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 524 4611 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/WWL
rlabel locali 4538 386 4568 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/RWL
rlabel locali 4102 386 4132 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/RWL
rlabel locali 4523 468 4538 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/WBL
rlabel locali 4133 468 4148 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/WBLb
rlabel locali 4596 322 4611 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/RBL0
rlabel locali 4059 322 4074 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/RBL1
rlabel metal1 4319 510 4351 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/VDD
rlabel metal1 4319 284 4351 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/GND
rlabel polycont 4281 391 4311 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/junc0
rlabel polycont 4359 391 4389 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/junc1
rlabel ndiff 4132 322 4188 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 322 4538 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 524 4031 554 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/WWL
rlabel locali 3958 386 3988 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/RWL
rlabel locali 3522 386 3552 420 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/RWL
rlabel locali 3943 468 3958 497 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/WBL
rlabel locali 3553 468 3568 496 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/WBLb
rlabel locali 4016 322 4031 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/RBL0
rlabel locali 3479 322 3494 364 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/RBL1
rlabel metal1 3739 510 3771 524 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/VDD
rlabel metal1 3739 284 3771 298 7 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/GND
rlabel polycont 3701 391 3731 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/junc0
rlabel polycont 3779 391 3809 425 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/junc1
rlabel ndiff 3552 322 3608 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 322 3958 350 1 10T_8x8_magic_0/10T_1x8_magic_5/10T_toy_magic_0/RWL0_junc
rlabel poly -1 254 29 284 1 10T_8x8_magic_0/10T_1x8_magic_4/WWL
rlabel metal1 -1 116 14 150 1 10T_8x8_magic_0/10T_1x8_magic_4/RWL
rlabel corelocali 73 198 88 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_0
rlabel corelocali 463 198 478 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_0
rlabel corelocali -1 52 14 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_0
rlabel corelocali 536 52 551 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_0
rlabel corelocali 653 198 668 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_1
rlabel corelocali 1043 198 1058 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_1
rlabel corelocali 579 52 594 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_1
rlabel corelocali 1116 52 1131 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_1
rlabel corelocali 1233 198 1248 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_2
rlabel corelocali 1623 198 1638 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_2
rlabel corelocali 1159 52 1174 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_2
rlabel corelocali 1696 52 1711 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_2
rlabel corelocali 1813 198 1828 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_3
rlabel corelocali 2203 198 2218 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_3
rlabel corelocali 1739 52 1754 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_3
rlabel corelocali 2276 52 2291 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_3
rlabel corelocali 2393 198 2408 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_4
rlabel corelocali 2783 198 2798 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_4
rlabel corelocali 2319 52 2334 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_4
rlabel corelocali 2856 52 2871 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_4
rlabel corelocali 2973 198 2988 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_5
rlabel corelocali 3363 198 3378 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_5
rlabel corelocali 2899 52 2914 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_5
rlabel corelocali 3436 52 3451 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_5
rlabel corelocali 3553 198 3568 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_6
rlabel corelocali 3943 198 3958 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_6
rlabel corelocali 3479 52 3494 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_6
rlabel corelocali 4016 52 4031 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_6
rlabel corelocali 4133 198 4148 226 1 10T_8x8_magic_0/10T_1x8_magic_4/WBLb_7
rlabel corelocali 4523 198 4538 227 1 10T_8x8_magic_0/10T_1x8_magic_4/WBL_7
rlabel corelocali 4059 52 4074 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL1_7
rlabel corelocali 4596 52 4611 94 1 10T_8x8_magic_0/10T_1x8_magic_4/RBL0_7
rlabel metal1 -1 240 14 254 1 10T_8x8_magic_0/10T_1x8_magic_4/VDD
rlabel metal1 -1 14 14 28 1 10T_8x8_magic_0/10T_1x8_magic_4/GND
rlabel poly -1 254 551 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/WWL
rlabel locali 478 116 508 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/RWL
rlabel locali 42 116 72 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/RWL
rlabel locali 463 198 478 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/WBL
rlabel locali 73 198 88 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/WBLb
rlabel locali 536 52 551 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/RBL0
rlabel locali -1 52 14 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/RBL1
rlabel metal1 259 240 291 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/VDD
rlabel metal1 259 14 291 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/GND
rlabel polycont 221 121 251 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/junc0
rlabel polycont 299 121 329 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/junc1
rlabel ndiff 72 52 128 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 52 478 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_7/RWL0_junc
rlabel poly 579 254 1131 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/WWL
rlabel locali 1058 116 1088 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/RWL
rlabel locali 622 116 652 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/RWL
rlabel locali 1043 198 1058 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/WBL
rlabel locali 653 198 668 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/WBLb
rlabel locali 1116 52 1131 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/RBL0
rlabel locali 579 52 594 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/RBL1
rlabel metal1 839 240 871 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/VDD
rlabel metal1 839 14 871 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/GND
rlabel polycont 801 121 831 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/junc0
rlabel polycont 879 121 909 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/junc1
rlabel ndiff 652 52 708 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 52 1058 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 254 1711 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/WWL
rlabel locali 1638 116 1668 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/RWL
rlabel locali 1202 116 1232 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/RWL
rlabel locali 1623 198 1638 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/WBL
rlabel locali 1233 198 1248 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/WBLb
rlabel locali 1696 52 1711 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/RBL0
rlabel locali 1159 52 1174 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/RBL1
rlabel metal1 1419 240 1451 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/VDD
rlabel metal1 1419 14 1451 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/GND
rlabel polycont 1381 121 1411 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/junc0
rlabel polycont 1459 121 1489 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/junc1
rlabel ndiff 1232 52 1288 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 52 1638 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 254 2291 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/WWL
rlabel locali 2218 116 2248 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/RWL
rlabel locali 1782 116 1812 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/RWL
rlabel locali 2203 198 2218 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/WBL
rlabel locali 1813 198 1828 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/WBLb
rlabel locali 2276 52 2291 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/RBL0
rlabel locali 1739 52 1754 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/RBL1
rlabel metal1 1999 240 2031 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/VDD
rlabel metal1 1999 14 2031 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/GND
rlabel polycont 1961 121 1991 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/junc0
rlabel polycont 2039 121 2069 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/junc1
rlabel ndiff 1812 52 1868 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 52 2218 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 254 2871 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/WWL
rlabel locali 2798 116 2828 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/RWL
rlabel locali 2362 116 2392 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/RWL
rlabel locali 2783 198 2798 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/WBL
rlabel locali 2393 198 2408 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/WBLb
rlabel locali 2856 52 2871 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/RBL0
rlabel locali 2319 52 2334 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/RBL1
rlabel metal1 2579 240 2611 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/VDD
rlabel metal1 2579 14 2611 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/GND
rlabel polycont 2541 121 2571 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/junc0
rlabel polycont 2619 121 2649 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/junc1
rlabel ndiff 2392 52 2448 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 52 2798 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 254 3451 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/WWL
rlabel locali 3378 116 3408 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/RWL
rlabel locali 2942 116 2972 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/RWL
rlabel locali 3363 198 3378 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/WBL
rlabel locali 2973 198 2988 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/WBLb
rlabel locali 3436 52 3451 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/RBL0
rlabel locali 2899 52 2914 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/RBL1
rlabel metal1 3159 240 3191 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/VDD
rlabel metal1 3159 14 3191 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/GND
rlabel polycont 3121 121 3151 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/junc0
rlabel polycont 3199 121 3229 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/junc1
rlabel ndiff 2972 52 3028 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 52 3378 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 254 4611 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/WWL
rlabel locali 4538 116 4568 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/RWL
rlabel locali 4102 116 4132 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/RWL
rlabel locali 4523 198 4538 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/WBL
rlabel locali 4133 198 4148 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/WBLb
rlabel locali 4596 52 4611 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/RBL0
rlabel locali 4059 52 4074 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/RBL1
rlabel metal1 4319 240 4351 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/VDD
rlabel metal1 4319 14 4351 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/GND
rlabel polycont 4281 121 4311 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/junc0
rlabel polycont 4359 121 4389 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/junc1
rlabel ndiff 4132 52 4188 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 52 4538 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 254 4031 284 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/WWL
rlabel locali 3958 116 3988 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/RWL
rlabel locali 3522 116 3552 150 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/RWL
rlabel locali 3943 198 3958 227 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/WBL
rlabel locali 3553 198 3568 226 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/WBLb
rlabel locali 4016 52 4031 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/RBL0
rlabel locali 3479 52 3494 94 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/RBL1
rlabel metal1 3739 240 3771 254 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/VDD
rlabel metal1 3739 14 3771 28 7 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/GND
rlabel polycont 3701 121 3731 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/junc0
rlabel polycont 3779 121 3809 155 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/junc1
rlabel ndiff 3552 52 3608 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 52 3958 80 1 10T_8x8_magic_0/10T_1x8_magic_4/10T_toy_magic_0/RWL0_junc
rlabel metal1 -1 1736 14 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/RWL
rlabel corelocali 73 1818 88 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_0
rlabel corelocali 463 1818 478 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_0
rlabel corelocali -1 1672 14 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_0
rlabel corelocali 536 1672 551 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_0
rlabel corelocali 653 1818 668 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_1
rlabel corelocali 1043 1818 1058 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_1
rlabel corelocali 579 1672 594 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_1
rlabel corelocali 1116 1672 1131 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_1
rlabel corelocali 1233 1818 1248 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_2
rlabel corelocali 1623 1818 1638 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_2
rlabel corelocali 1159 1672 1174 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_2
rlabel corelocali 1696 1672 1711 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_2
rlabel corelocali 1813 1818 1828 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_3
rlabel corelocali 2203 1818 2218 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_3
rlabel corelocali 1739 1672 1754 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_3
rlabel corelocali 2276 1672 2291 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_3
rlabel corelocali 2393 1818 2408 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_4
rlabel corelocali 2783 1818 2798 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_4
rlabel corelocali 2319 1672 2334 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_4
rlabel corelocali 2856 1672 2871 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_4
rlabel corelocali 2973 1818 2988 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_5
rlabel corelocali 3363 1818 3378 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_5
rlabel corelocali 2899 1672 2914 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_5
rlabel corelocali 3436 1672 3451 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_5
rlabel corelocali 3553 1818 3568 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_6
rlabel corelocali 3943 1818 3958 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_6
rlabel corelocali 3479 1672 3494 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_6
rlabel corelocali 4016 1672 4031 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_6
rlabel corelocali 4133 1818 4148 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/WBLb_7
rlabel corelocali 4523 1818 4538 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/WBL_7
rlabel corelocali 4059 1672 4074 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL1_7
rlabel corelocali 4596 1672 4611 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/RBL0_7
rlabel metal1 -1 1860 14 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/VDD
rlabel metal1 -1 1634 14 1648 1 10T_8x8_magic_0/10T_1x8_magic_3/GND
rlabel locali 478 1736 508 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/RWL
rlabel locali 42 1736 72 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/RWL
rlabel locali 463 1818 478 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/WBL
rlabel locali 73 1818 88 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/WBLb
rlabel locali 536 1672 551 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/RBL0
rlabel locali -1 1672 14 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/RBL1
rlabel metal1 259 1860 291 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/VDD
rlabel metal1 259 1634 291 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/GND
rlabel polycont 221 1741 251 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/junc0
rlabel polycont 299 1741 329 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/junc1
rlabel ndiff 72 1672 128 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 1672 478 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_7/RWL0_junc
rlabel locali 1058 1736 1088 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/RWL
rlabel locali 622 1736 652 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/RWL
rlabel locali 1043 1818 1058 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/WBL
rlabel locali 653 1818 668 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/WBLb
rlabel locali 1116 1672 1131 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/RBL0
rlabel locali 579 1672 594 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/RBL1
rlabel metal1 839 1860 871 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/VDD
rlabel metal1 839 1634 871 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/GND
rlabel polycont 801 1741 831 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/junc0
rlabel polycont 879 1741 909 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/junc1
rlabel ndiff 652 1672 708 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 1672 1058 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_6/RWL0_junc
rlabel locali 1638 1736 1668 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/RWL
rlabel locali 1202 1736 1232 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/RWL
rlabel locali 1623 1818 1638 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/WBL
rlabel locali 1233 1818 1248 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/WBLb
rlabel locali 1696 1672 1711 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/RBL0
rlabel locali 1159 1672 1174 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/RBL1
rlabel metal1 1419 1860 1451 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/VDD
rlabel metal1 1419 1634 1451 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/GND
rlabel polycont 1381 1741 1411 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/junc0
rlabel polycont 1459 1741 1489 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/junc1
rlabel ndiff 1232 1672 1288 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 1672 1638 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_5/RWL0_junc
rlabel locali 2218 1736 2248 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/RWL
rlabel locali 1782 1736 1812 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/RWL
rlabel locali 2203 1818 2218 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/WBL
rlabel locali 1813 1818 1828 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/WBLb
rlabel locali 2276 1672 2291 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/RBL0
rlabel locali 1739 1672 1754 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/RBL1
rlabel metal1 1999 1860 2031 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/VDD
rlabel metal1 1999 1634 2031 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/GND
rlabel polycont 1961 1741 1991 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/junc0
rlabel polycont 2039 1741 2069 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/junc1
rlabel ndiff 1812 1672 1868 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 1672 2218 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_4/RWL0_junc
rlabel locali 2798 1736 2828 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/RWL
rlabel locali 2362 1736 2392 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/RWL
rlabel locali 2783 1818 2798 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/WBL
rlabel locali 2393 1818 2408 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/WBLb
rlabel locali 2856 1672 2871 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/RBL0
rlabel locali 2319 1672 2334 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/RBL1
rlabel metal1 2579 1860 2611 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/VDD
rlabel metal1 2579 1634 2611 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/GND
rlabel polycont 2541 1741 2571 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/junc0
rlabel polycont 2619 1741 2649 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/junc1
rlabel ndiff 2392 1672 2448 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 1672 2798 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_3/RWL0_junc
rlabel locali 3378 1736 3408 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/RWL
rlabel locali 2942 1736 2972 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/RWL
rlabel locali 3363 1818 3378 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/WBL
rlabel locali 2973 1818 2988 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/WBLb
rlabel locali 3436 1672 3451 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/RBL0
rlabel locali 2899 1672 2914 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/RBL1
rlabel metal1 3159 1860 3191 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/VDD
rlabel metal1 3159 1634 3191 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/GND
rlabel polycont 3121 1741 3151 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/junc0
rlabel polycont 3199 1741 3229 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/junc1
rlabel ndiff 2972 1672 3028 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 1672 3378 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_2/RWL0_junc
rlabel locali 4538 1736 4568 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/RWL
rlabel locali 4102 1736 4132 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/RWL
rlabel locali 4523 1818 4538 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/WBL
rlabel locali 4133 1818 4148 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/WBLb
rlabel locali 4596 1672 4611 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/RBL0
rlabel locali 4059 1672 4074 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/RBL1
rlabel metal1 4319 1860 4351 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/VDD
rlabel metal1 4319 1634 4351 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/GND
rlabel polycont 4281 1741 4311 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/junc0
rlabel polycont 4359 1741 4389 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/junc1
rlabel ndiff 4132 1672 4188 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 1672 4538 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_1/RWL0_junc
rlabel locali 3958 1736 3988 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/RWL
rlabel locali 3522 1736 3552 1770 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/RWL
rlabel locali 3943 1818 3958 1847 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/WBL
rlabel locali 3553 1818 3568 1846 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/WBLb
rlabel locali 4016 1672 4031 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/RBL0
rlabel locali 3479 1672 3494 1714 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/RBL1
rlabel metal1 3739 1860 3771 1874 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/VDD
rlabel metal1 3739 1634 3771 1648 7 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/GND
rlabel polycont 3701 1741 3731 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/junc0
rlabel polycont 3779 1741 3809 1775 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/junc1
rlabel ndiff 3552 1672 3608 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 1672 3958 1700 1 10T_8x8_magic_0/10T_1x8_magic_3/10T_toy_magic_0/RWL0_junc
rlabel corelocali 653 2088 668 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_1
rlabel corelocali 1043 2088 1058 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_1
rlabel corelocali 1116 1942 1131 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_1
rlabel corelocali 1233 2088 1248 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_2
rlabel corelocali 1623 2088 1638 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_2
rlabel corelocali 1159 1942 1174 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_2
rlabel corelocali 1696 1942 1711 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_2
rlabel corelocali 1813 2088 1828 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_3
rlabel corelocali 2203 2088 2218 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_3
rlabel corelocali 1739 1942 1754 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_3
rlabel corelocali 2276 1942 2291 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_3
rlabel corelocali 2393 2088 2408 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_4
rlabel corelocali 2783 2088 2798 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_4
rlabel corelocali 2319 1942 2334 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_4
rlabel corelocali 2856 1942 2871 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_4
rlabel corelocali 2973 2088 2988 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_5
rlabel corelocali 3363 2088 3378 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_5
rlabel corelocali 2899 1942 2914 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_5
rlabel corelocali 3436 1942 3451 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_5
rlabel corelocali 3553 2088 3568 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_6
rlabel corelocali 3943 2088 3958 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_6
rlabel corelocali 3479 1942 3494 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_6
rlabel corelocali 4016 1942 4031 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_6
rlabel corelocali 4133 2088 4148 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/WBLb_7
rlabel corelocali 4523 2088 4538 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/WBL_7
rlabel corelocali 4059 1942 4074 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_7
rlabel corelocali 4596 1942 4611 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_7
rlabel locali 1058 2006 1088 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/RWL
rlabel locali 622 2006 652 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/RWL
rlabel locali 1043 2088 1058 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/WBL
rlabel locali 653 2088 668 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/WBLb
rlabel locali 1116 1942 1131 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/RBL0
rlabel locali 579 1942 594 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/RBL1
rlabel metal1 839 2130 871 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/VDD
rlabel metal1 839 1904 871 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/GND
rlabel polycont 801 2011 831 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/junc0
rlabel polycont 879 2011 909 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/junc1
rlabel ndiff 652 1942 708 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 1942 1058 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_6/RWL0_junc
rlabel locali 1638 2006 1668 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/RWL
rlabel locali 1202 2006 1232 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/RWL
rlabel locali 1623 2088 1638 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/WBL
rlabel locali 1233 2088 1248 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/WBLb
rlabel locali 1696 1942 1711 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/RBL0
rlabel locali 1159 1942 1174 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/RBL1
rlabel metal1 1419 2130 1451 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/VDD
rlabel metal1 1419 1904 1451 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/GND
rlabel polycont 1381 2011 1411 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/junc0
rlabel polycont 1459 2011 1489 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/junc1
rlabel ndiff 1232 1942 1288 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 1942 1638 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_5/RWL0_junc
rlabel locali 2218 2006 2248 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/RWL
rlabel locali 1782 2006 1812 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/RWL
rlabel locali 2203 2088 2218 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/WBL
rlabel locali 1813 2088 1828 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/WBLb
rlabel locali 2276 1942 2291 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/RBL0
rlabel locali 1739 1942 1754 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/RBL1
rlabel metal1 1999 2130 2031 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/VDD
rlabel metal1 1999 1904 2031 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/GND
rlabel polycont 1961 2011 1991 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/junc0
rlabel polycont 2039 2011 2069 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/junc1
rlabel ndiff 1812 1942 1868 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 1942 2218 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_4/RWL0_junc
rlabel locali 2798 2006 2828 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/RWL
rlabel locali 2362 2006 2392 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/RWL
rlabel locali 2783 2088 2798 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/WBL
rlabel locali 2393 2088 2408 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/WBLb
rlabel locali 2856 1942 2871 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/RBL0
rlabel locali 2319 1942 2334 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/RBL1
rlabel metal1 2579 2130 2611 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/VDD
rlabel metal1 2579 1904 2611 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/GND
rlabel polycont 2541 2011 2571 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/junc0
rlabel polycont 2619 2011 2649 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/junc1
rlabel ndiff 2392 1942 2448 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 1942 2798 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_3/RWL0_junc
rlabel locali 3378 2006 3408 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/RWL
rlabel locali 2942 2006 2972 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/RWL
rlabel locali 3363 2088 3378 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/WBL
rlabel locali 2973 2088 2988 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/WBLb
rlabel locali 3436 1942 3451 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/RBL0
rlabel locali 2899 1942 2914 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/RBL1
rlabel metal1 3159 2130 3191 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/VDD
rlabel metal1 3159 1904 3191 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/GND
rlabel polycont 3121 2011 3151 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/junc0
rlabel polycont 3199 2011 3229 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/junc1
rlabel ndiff 2972 1942 3028 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 1942 3378 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_2/RWL0_junc
rlabel locali 4538 2006 4568 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/RWL
rlabel locali 4102 2006 4132 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/RWL
rlabel locali 4523 2088 4538 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/WBL
rlabel locali 4133 2088 4148 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/WBLb
rlabel locali 4596 1942 4611 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/RBL0
rlabel locali 4059 1942 4074 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/RBL1
rlabel metal1 4319 2130 4351 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/VDD
rlabel metal1 4319 1904 4351 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/GND
rlabel polycont 4281 2011 4311 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/junc0
rlabel polycont 4359 2011 4389 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/junc1
rlabel ndiff 4132 1942 4188 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 1942 4538 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_1/RWL0_junc
rlabel locali 3958 2006 3988 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/RWL
rlabel locali 3522 2006 3552 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/RWL
rlabel locali 3943 2088 3958 2117 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/WBL
rlabel locali 3553 2088 3568 2116 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/WBLb
rlabel locali 4016 1942 4031 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/RBL0
rlabel locali 3479 1942 3494 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/RBL1
rlabel metal1 3739 2130 3771 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/VDD
rlabel metal1 3739 1904 3771 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/GND
rlabel polycont 3701 2011 3731 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/junc0
rlabel polycont 3779 2011 3809 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/junc1
rlabel ndiff 3552 1942 3608 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 1942 3958 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_0/RWL0_junc
rlabel metal1 -1 1196 14 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/RWL
rlabel corelocali 73 1278 88 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_0
rlabel corelocali 463 1278 478 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_0
rlabel corelocali -1 1132 14 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_0
rlabel corelocali 536 1132 551 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_0
rlabel corelocali 653 1278 668 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_1
rlabel corelocali 1043 1278 1058 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_1
rlabel corelocali 579 1132 594 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_1
rlabel corelocali 1116 1132 1131 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_1
rlabel corelocali 1233 1278 1248 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_2
rlabel corelocali 1623 1278 1638 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_2
rlabel corelocali 1159 1132 1174 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_2
rlabel corelocali 1696 1132 1711 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_2
rlabel corelocali 1813 1278 1828 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_3
rlabel corelocali 2203 1278 2218 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_3
rlabel corelocali 1739 1132 1754 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_3
rlabel corelocali 2276 1132 2291 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_3
rlabel corelocali 2393 1278 2408 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_4
rlabel corelocali 2783 1278 2798 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_4
rlabel corelocali 2319 1132 2334 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_4
rlabel corelocali 2856 1132 2871 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_4
rlabel corelocali 2973 1278 2988 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_5
rlabel corelocali 3363 1278 3378 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_5
rlabel corelocali 2899 1132 2914 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_5
rlabel corelocali 3436 1132 3451 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_5
rlabel corelocali 3553 1278 3568 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_6
rlabel corelocali 3943 1278 3958 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_6
rlabel corelocali 3479 1132 3494 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_6
rlabel corelocali 4016 1132 4031 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_6
rlabel corelocali 4133 1278 4148 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/WBLb_7
rlabel corelocali 4523 1278 4538 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/WBL_7
rlabel corelocali 4059 1132 4074 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL1_7
rlabel corelocali 4596 1132 4611 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/RBL0_7
rlabel metal1 -1 1320 14 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/VDD
rlabel metal1 -1 1094 14 1108 1 10T_8x8_magic_0/10T_1x8_magic_1/GND
rlabel locali 478 1196 508 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/RWL
rlabel locali 42 1196 72 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/RWL
rlabel locali 463 1278 478 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/WBL
rlabel locali 73 1278 88 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/WBLb
rlabel locali 536 1132 551 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/RBL0
rlabel locali -1 1132 14 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/RBL1
rlabel metal1 259 1320 291 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/VDD
rlabel metal1 259 1094 291 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/GND
rlabel polycont 221 1201 251 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/junc0
rlabel polycont 299 1201 329 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/junc1
rlabel ndiff 72 1132 128 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 1132 478 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_7/RWL0_junc
rlabel locali 1058 1196 1088 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/RWL
rlabel locali 622 1196 652 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/RWL
rlabel locali 1043 1278 1058 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/WBL
rlabel locali 653 1278 668 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/WBLb
rlabel locali 1116 1132 1131 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/RBL0
rlabel locali 579 1132 594 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/RBL1
rlabel metal1 839 1320 871 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/VDD
rlabel metal1 839 1094 871 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/GND
rlabel polycont 801 1201 831 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/junc0
rlabel polycont 879 1201 909 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/junc1
rlabel ndiff 652 1132 708 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 1132 1058 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_6/RWL0_junc
rlabel locali 1638 1196 1668 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/RWL
rlabel locali 1202 1196 1232 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/RWL
rlabel locali 1623 1278 1638 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/WBL
rlabel locali 1233 1278 1248 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/WBLb
rlabel locali 1696 1132 1711 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/RBL0
rlabel locali 1159 1132 1174 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/RBL1
rlabel metal1 1419 1320 1451 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/VDD
rlabel metal1 1419 1094 1451 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/GND
rlabel polycont 1381 1201 1411 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/junc0
rlabel polycont 1459 1201 1489 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/junc1
rlabel ndiff 1232 1132 1288 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 1132 1638 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_5/RWL0_junc
rlabel locali 2218 1196 2248 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/RWL
rlabel locali 1782 1196 1812 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/RWL
rlabel locali 2203 1278 2218 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/WBL
rlabel locali 1813 1278 1828 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/WBLb
rlabel locali 2276 1132 2291 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/RBL0
rlabel locali 1739 1132 1754 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/RBL1
rlabel metal1 1999 1320 2031 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/VDD
rlabel metal1 1999 1094 2031 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/GND
rlabel polycont 1961 1201 1991 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/junc0
rlabel polycont 2039 1201 2069 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/junc1
rlabel ndiff 1812 1132 1868 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 1132 2218 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_4/RWL0_junc
rlabel locali 2798 1196 2828 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/RWL
rlabel locali 2362 1196 2392 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/RWL
rlabel locali 2783 1278 2798 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/WBL
rlabel locali 2393 1278 2408 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/WBLb
rlabel locali 2856 1132 2871 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/RBL0
rlabel locali 2319 1132 2334 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/RBL1
rlabel metal1 2579 1320 2611 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/VDD
rlabel metal1 2579 1094 2611 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/GND
rlabel polycont 2541 1201 2571 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/junc0
rlabel polycont 2619 1201 2649 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/junc1
rlabel ndiff 2392 1132 2448 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 1132 2798 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_3/RWL0_junc
rlabel locali 3378 1196 3408 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/RWL
rlabel locali 2942 1196 2972 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/RWL
rlabel locali 3363 1278 3378 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/WBL
rlabel locali 2973 1278 2988 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/WBLb
rlabel locali 3436 1132 3451 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/RBL0
rlabel locali 2899 1132 2914 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/RBL1
rlabel metal1 3159 1320 3191 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/VDD
rlabel metal1 3159 1094 3191 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/GND
rlabel polycont 3121 1201 3151 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/junc0
rlabel polycont 3199 1201 3229 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/junc1
rlabel ndiff 2972 1132 3028 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 1132 3378 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_2/RWL0_junc
rlabel locali 4538 1196 4568 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/RWL
rlabel locali 4102 1196 4132 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/RWL
rlabel locali 4523 1278 4538 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/WBL
rlabel locali 4133 1278 4148 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/WBLb
rlabel locali 4596 1132 4611 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/RBL0
rlabel locali 4059 1132 4074 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/RBL1
rlabel metal1 4319 1320 4351 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/VDD
rlabel metal1 4319 1094 4351 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/GND
rlabel polycont 4281 1201 4311 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/junc0
rlabel polycont 4359 1201 4389 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/junc1
rlabel ndiff 4132 1132 4188 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 1132 4538 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_1/RWL0_junc
rlabel locali 3958 1196 3988 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/RWL
rlabel locali 3522 1196 3552 1230 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/RWL
rlabel locali 3943 1278 3958 1307 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/WBL
rlabel locali 3553 1278 3568 1306 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/WBLb
rlabel locali 4016 1132 4031 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/RBL0
rlabel locali 3479 1132 3494 1174 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/RBL1
rlabel metal1 3739 1320 3771 1334 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/VDD
rlabel metal1 3739 1094 3771 1108 7 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/GND
rlabel polycont 3701 1201 3731 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/junc0
rlabel polycont 3779 1201 3809 1235 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/junc1
rlabel ndiff 3552 1132 3608 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 1132 3958 1160 1 10T_8x8_magic_0/10T_1x8_magic_1/10T_toy_magic_0/RWL0_junc
rlabel metal1 -1 1466 14 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/RWL
rlabel corelocali 73 1548 88 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_0
rlabel corelocali 463 1548 478 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_0
rlabel corelocali -1 1402 14 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_0
rlabel corelocali 536 1402 551 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_0
rlabel corelocali 653 1548 668 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_1
rlabel corelocali 1043 1548 1058 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_1
rlabel corelocali 579 1402 594 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_1
rlabel corelocali 1116 1402 1131 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_1
rlabel corelocali 1233 1548 1248 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_2
rlabel corelocali 1623 1548 1638 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_2
rlabel corelocali 1159 1402 1174 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_2
rlabel corelocali 1696 1402 1711 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_2
rlabel corelocali 1813 1548 1828 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_3
rlabel corelocali 2203 1548 2218 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_3
rlabel corelocali 1739 1402 1754 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_3
rlabel corelocali 2276 1402 2291 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_3
rlabel corelocali 2393 1548 2408 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_4
rlabel corelocali 2783 1548 2798 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_4
rlabel corelocali 2319 1402 2334 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_4
rlabel corelocali 2856 1402 2871 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_4
rlabel corelocali 2973 1548 2988 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_5
rlabel corelocali 3363 1548 3378 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_5
rlabel corelocali 2899 1402 2914 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_5
rlabel corelocali 3436 1402 3451 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_5
rlabel corelocali 3553 1548 3568 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_6
rlabel corelocali 3943 1548 3958 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_6
rlabel corelocali 3479 1402 3494 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_6
rlabel corelocali 4016 1402 4031 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_6
rlabel corelocali 4133 1548 4148 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/WBLb_7
rlabel corelocali 4523 1548 4538 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/WBL_7
rlabel corelocali 4059 1402 4074 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL1_7
rlabel corelocali 4596 1402 4611 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/RBL0_7
rlabel metal1 -1 1590 14 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/VDD
rlabel metal1 -1 1364 14 1378 1 10T_8x8_magic_0/10T_1x8_magic_0/GND
rlabel locali 478 1466 508 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/RWL
rlabel locali 42 1466 72 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/RWL
rlabel locali 463 1548 478 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/WBL
rlabel locali 73 1548 88 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/WBLb
rlabel locali 536 1402 551 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/RBL0
rlabel locali -1 1402 14 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/RBL1
rlabel metal1 259 1590 291 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/VDD
rlabel metal1 259 1364 291 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/GND
rlabel polycont 221 1471 251 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/junc0
rlabel polycont 299 1471 329 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/junc1
rlabel ndiff 72 1402 128 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 1402 478 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_7/RWL0_junc
rlabel locali 1058 1466 1088 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/RWL
rlabel locali 622 1466 652 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/RWL
rlabel locali 1043 1548 1058 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/WBL
rlabel locali 653 1548 668 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/WBLb
rlabel locali 1116 1402 1131 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/RBL0
rlabel locali 579 1402 594 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/RBL1
rlabel metal1 839 1590 871 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/VDD
rlabel metal1 839 1364 871 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/GND
rlabel polycont 801 1471 831 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/junc0
rlabel polycont 879 1471 909 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/junc1
rlabel ndiff 652 1402 708 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 1402 1058 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_6/RWL0_junc
rlabel locali 1638 1466 1668 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/RWL
rlabel locali 1202 1466 1232 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/RWL
rlabel locali 1623 1548 1638 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/WBL
rlabel locali 1233 1548 1248 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/WBLb
rlabel locali 1696 1402 1711 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/RBL0
rlabel locali 1159 1402 1174 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/RBL1
rlabel metal1 1419 1590 1451 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/VDD
rlabel metal1 1419 1364 1451 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/GND
rlabel polycont 1381 1471 1411 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/junc0
rlabel polycont 1459 1471 1489 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/junc1
rlabel ndiff 1232 1402 1288 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 1402 1638 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_5/RWL0_junc
rlabel locali 2218 1466 2248 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/RWL
rlabel locali 1782 1466 1812 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/RWL
rlabel locali 2203 1548 2218 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/WBL
rlabel locali 1813 1548 1828 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/WBLb
rlabel locali 2276 1402 2291 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/RBL0
rlabel locali 1739 1402 1754 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/RBL1
rlabel metal1 1999 1590 2031 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/VDD
rlabel metal1 1999 1364 2031 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/GND
rlabel polycont 1961 1471 1991 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/junc0
rlabel polycont 2039 1471 2069 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/junc1
rlabel ndiff 1812 1402 1868 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 1402 2218 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_4/RWL0_junc
rlabel locali 2798 1466 2828 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/RWL
rlabel locali 2362 1466 2392 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/RWL
rlabel locali 2783 1548 2798 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/WBL
rlabel locali 2393 1548 2408 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/WBLb
rlabel locali 2856 1402 2871 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/RBL0
rlabel locali 2319 1402 2334 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/RBL1
rlabel metal1 2579 1590 2611 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/VDD
rlabel metal1 2579 1364 2611 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/GND
rlabel polycont 2541 1471 2571 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/junc0
rlabel polycont 2619 1471 2649 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/junc1
rlabel ndiff 2392 1402 2448 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 1402 2798 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_3/RWL0_junc
rlabel locali 3378 1466 3408 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/RWL
rlabel locali 2942 1466 2972 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/RWL
rlabel locali 3363 1548 3378 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/WBL
rlabel locali 2973 1548 2988 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/WBLb
rlabel locali 3436 1402 3451 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/RBL0
rlabel locali 2899 1402 2914 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/RBL1
rlabel metal1 3159 1590 3191 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/VDD
rlabel metal1 3159 1364 3191 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/GND
rlabel polycont 3121 1471 3151 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/junc0
rlabel polycont 3199 1471 3229 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/junc1
rlabel ndiff 2972 1402 3028 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 1402 3378 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_2/RWL0_junc
rlabel locali 4538 1466 4568 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/RWL
rlabel locali 4102 1466 4132 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/RWL
rlabel locali 4523 1548 4538 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/WBL
rlabel locali 4133 1548 4148 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/WBLb
rlabel locali 4596 1402 4611 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/RBL0
rlabel locali 4059 1402 4074 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/RBL1
rlabel metal1 4319 1590 4351 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/VDD
rlabel metal1 4319 1364 4351 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/GND
rlabel polycont 4281 1471 4311 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/junc0
rlabel polycont 4359 1471 4389 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/junc1
rlabel ndiff 4132 1402 4188 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 1402 4538 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_1/RWL0_junc
rlabel locali 3958 1466 3988 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/RWL
rlabel locali 3522 1466 3552 1500 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/RWL
rlabel locali 3943 1548 3958 1577 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/WBL
rlabel locali 3553 1548 3568 1576 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/WBLb
rlabel locali 4016 1402 4031 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/RBL0
rlabel locali 3479 1402 3494 1444 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/RBL1
rlabel metal1 3739 1590 3771 1604 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/VDD
rlabel metal1 3739 1364 3771 1378 7 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/GND
rlabel polycont 3701 1471 3731 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/junc0
rlabel polycont 3779 1471 3809 1505 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/junc1
rlabel ndiff 3552 1402 3608 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 1402 3958 1430 1 10T_8x8_magic_0/10T_1x8_magic_0/10T_toy_magic_0/RWL0_junc
rlabel locali -1 -2108 14 -2066 1 10T_8x8_magic_1/RBL1_0
rlabel locali 536 -2108 551 -2066 1 10T_8x8_magic_1/RBL0_0
rlabel locali 579 -2108 594 -2066 1 10T_8x8_magic_1/RBL1_1
rlabel locali 1116 -2108 1131 -2066 1 10T_8x8_magic_1/RBL0_1
rlabel locali 1159 -2108 1174 -2066 1 10T_8x8_magic_1/RBL1_2
rlabel locali 1696 -2108 1711 -2066 1 10T_8x8_magic_1/RBL0_2
rlabel locali 1739 -2108 1754 -2066 1 10T_8x8_magic_1/RBL1_3
rlabel locali 2276 -2108 2291 -2066 1 10T_8x8_magic_1/RBL0_3
rlabel locali 2319 -2108 2334 -2066 1 10T_8x8_magic_1/RBL1_4
rlabel locali 2856 -2108 2871 -2066 1 10T_8x8_magic_1/RBL0_4
rlabel locali 2899 -2108 2914 -2066 1 10T_8x8_magic_1/RBL1_5
rlabel locali 3436 -2108 3451 -2066 1 10T_8x8_magic_1/RBL0_5
rlabel locali 3479 -2108 3494 -2066 1 10T_8x8_magic_1/RBL1_6
rlabel locali 4016 -2108 4031 -2066 1 10T_8x8_magic_1/RBL0_6
rlabel locali 4059 -2108 4074 -2066 1 10T_8x8_magic_1/RBL1_7
rlabel locali 4596 -2108 4611 -2066 1 10T_8x8_magic_1/RBL0_7
rlabel locali 463 -1962 478 -1933 1 10T_8x8_magic_1/WBL_0
rlabel locali 73 -1962 88 -1934 1 10T_8x8_magic_1/WBLb_0
rlabel locali 1043 -1962 1058 -1933 1 10T_8x8_magic_1/WBL_1
rlabel locali 653 -1962 668 -1934 1 10T_8x8_magic_1/WBLb_1
rlabel locali 1623 -1962 1638 -1933 1 10T_8x8_magic_1/WBL_2
rlabel locali 1233 -1962 1248 -1934 1 10T_8x8_magic_1/WBLb_2
rlabel locali 2203 -1962 2218 -1933 1 10T_8x8_magic_1/WBL_3
rlabel locali 1813 -1962 1828 -1934 1 10T_8x8_magic_1/WBLb_3
rlabel locali 2783 -1962 2798 -1933 1 10T_8x8_magic_1/WBL_4
rlabel locali 2393 -1962 2408 -1934 1 10T_8x8_magic_1/WBLb_4
rlabel locali 3363 -1962 3378 -1933 1 10T_8x8_magic_1/WBL_5
rlabel locali 2973 -1962 2988 -1934 1 10T_8x8_magic_1/WBLb_5
rlabel locali 3943 -1962 3958 -1933 1 10T_8x8_magic_1/WBL_6
rlabel locali 3553 -1962 3568 -1934 1 10T_8x8_magic_1/WBLb_6
rlabel locali 4523 -1962 4538 -1933 1 10T_8x8_magic_1/WBL_7
rlabel locali 4133 -1962 4148 -1934 1 10T_8x8_magic_1/WBLb_7
rlabel poly -1 -16 29 14 1 10T_8x8_magic_1/WWL_0
rlabel metal1 -1 -154 14 -120 1 10T_8x8_magic_1/RWL_0
rlabel poly -1 -286 29 -256 1 10T_8x8_magic_1/WWL_1
rlabel metal1 -1 -424 14 -390 1 10T_8x8_magic_1/RWL_1
rlabel poly -1 -556 29 -526 1 10T_8x8_magic_1/WWL_2
rlabel metal1 -1 -694 14 -660 1 10T_8x8_magic_1/RWL_2
rlabel poly -1 -826 29 -796 1 10T_8x8_magic_1/WWL_3
rlabel metal1 -1 -964 14 -930 1 10T_8x8_magic_1/RWL_3
rlabel poly -1 -1096 29 -1066 1 10T_8x8_magic_1/WWL_4
rlabel metal1 -1 -1234 14 -1200 1 10T_8x8_magic_1/RWL_4
rlabel poly -1 -1366 29 -1336 1 10T_8x8_magic_1/WWL_5
rlabel metal1 -1 -1504 14 -1470 1 10T_8x8_magic_1/RWL_5
rlabel poly -1 -1636 29 -1606 1 10T_8x8_magic_1/WWL_6
rlabel metal1 -1 -1774 14 -1740 1 10T_8x8_magic_1/RWL_6
rlabel poly -1 -1906 29 -1876 1 10T_8x8_magic_1/WWL_7
rlabel metal1 -1 -2044 14 -2010 1 10T_8x8_magic_1/RWL_7
rlabel metal1 -1 -30 14 -16 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -256 14 -242 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -570 14 -556 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -840 14 -826 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -300 14 -286 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -1110 14 -1096 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -1650 14 -1636 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -1920 14 -1906 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -1380 14 -1366 1 10T_8x8_magic_1/VDD
rlabel metal1 -1 -1066 14 -1052 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -796 14 -782 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -526 14 -512 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -1336 14 -1322 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -2146 14 -2132 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -1876 14 -1862 1 10T_8x8_magic_1/GND
rlabel metal1 -1 -1606 14 -1592 1 10T_8x8_magic_1/GND
rlabel poly -1 -1366 29 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/WWL
rlabel metal1 -1 -1504 14 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/RWL
rlabel corelocali 73 -1422 88 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_0
rlabel corelocali 463 -1422 478 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_0
rlabel corelocali -1 -1568 14 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_0
rlabel corelocali 536 -1568 551 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_0
rlabel corelocali 653 -1422 668 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_1
rlabel corelocali 1043 -1422 1058 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_1
rlabel corelocali 579 -1568 594 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_1
rlabel corelocali 1116 -1568 1131 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_1
rlabel corelocali 1233 -1422 1248 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_2
rlabel corelocali 1623 -1422 1638 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_2
rlabel corelocali 1159 -1568 1174 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_2
rlabel corelocali 1696 -1568 1711 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_2
rlabel corelocali 1813 -1422 1828 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_3
rlabel corelocali 2203 -1422 2218 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_3
rlabel corelocali 1739 -1568 1754 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_3
rlabel corelocali 2276 -1568 2291 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_3
rlabel corelocali 2393 -1422 2408 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_4
rlabel corelocali 2783 -1422 2798 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_4
rlabel corelocali 2319 -1568 2334 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_4
rlabel corelocali 2856 -1568 2871 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_4
rlabel corelocali 2973 -1422 2988 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_5
rlabel corelocali 3363 -1422 3378 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_5
rlabel corelocali 2899 -1568 2914 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_5
rlabel corelocali 3436 -1568 3451 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_5
rlabel corelocali 3553 -1422 3568 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_6
rlabel corelocali 3943 -1422 3958 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_6
rlabel corelocali 3479 -1568 3494 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_6
rlabel corelocali 4016 -1568 4031 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_6
rlabel corelocali 4133 -1422 4148 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/WBLb_7
rlabel corelocali 4523 -1422 4538 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/WBL_7
rlabel corelocali 4059 -1568 4074 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL1_7
rlabel corelocali 4596 -1568 4611 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/RBL0_7
rlabel metal1 -1 -1380 14 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/VDD
rlabel metal1 -1 -1606 14 -1592 1 10T_8x8_magic_1/10T_1x8_magic_7/GND
rlabel poly -1 -1366 551 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/WWL
rlabel locali 478 -1504 508 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/RWL
rlabel locali 42 -1504 72 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/RWL
rlabel locali 463 -1422 478 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/WBL
rlabel locali 73 -1422 88 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/WBLb
rlabel locali 536 -1568 551 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/RBL0
rlabel locali -1 -1568 14 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/RBL1
rlabel metal1 259 -1380 291 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/VDD
rlabel metal1 259 -1606 291 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/GND
rlabel polycont 221 -1499 251 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/junc0
rlabel polycont 299 -1499 329 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/junc1
rlabel ndiff 72 -1568 128 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -1568 478 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -1366 1131 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/WWL
rlabel locali 1058 -1504 1088 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/RWL
rlabel locali 622 -1504 652 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/RWL
rlabel locali 1043 -1422 1058 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/WBL
rlabel locali 653 -1422 668 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/WBLb
rlabel locali 1116 -1568 1131 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/RBL0
rlabel locali 579 -1568 594 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/RBL1
rlabel metal1 839 -1380 871 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/VDD
rlabel metal1 839 -1606 871 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/GND
rlabel polycont 801 -1499 831 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/junc0
rlabel polycont 879 -1499 909 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/junc1
rlabel ndiff 652 -1568 708 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -1568 1058 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -1366 1711 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/WWL
rlabel locali 1638 -1504 1668 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/RWL
rlabel locali 1202 -1504 1232 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/RWL
rlabel locali 1623 -1422 1638 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/WBL
rlabel locali 1233 -1422 1248 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/WBLb
rlabel locali 1696 -1568 1711 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/RBL0
rlabel locali 1159 -1568 1174 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/RBL1
rlabel metal1 1419 -1380 1451 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/VDD
rlabel metal1 1419 -1606 1451 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/GND
rlabel polycont 1381 -1499 1411 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/junc0
rlabel polycont 1459 -1499 1489 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/junc1
rlabel ndiff 1232 -1568 1288 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -1568 1638 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -1366 2291 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/WWL
rlabel locali 2218 -1504 2248 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/RWL
rlabel locali 1782 -1504 1812 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/RWL
rlabel locali 2203 -1422 2218 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/WBL
rlabel locali 1813 -1422 1828 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/WBLb
rlabel locali 2276 -1568 2291 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/RBL0
rlabel locali 1739 -1568 1754 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/RBL1
rlabel metal1 1999 -1380 2031 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/VDD
rlabel metal1 1999 -1606 2031 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/GND
rlabel polycont 1961 -1499 1991 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/junc0
rlabel polycont 2039 -1499 2069 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/junc1
rlabel ndiff 1812 -1568 1868 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -1568 2218 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -1366 2871 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/WWL
rlabel locali 2798 -1504 2828 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/RWL
rlabel locali 2362 -1504 2392 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/RWL
rlabel locali 2783 -1422 2798 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/WBL
rlabel locali 2393 -1422 2408 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/WBLb
rlabel locali 2856 -1568 2871 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/RBL0
rlabel locali 2319 -1568 2334 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/RBL1
rlabel metal1 2579 -1380 2611 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/VDD
rlabel metal1 2579 -1606 2611 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/GND
rlabel polycont 2541 -1499 2571 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/junc0
rlabel polycont 2619 -1499 2649 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/junc1
rlabel ndiff 2392 -1568 2448 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -1568 2798 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -1366 3451 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/WWL
rlabel locali 3378 -1504 3408 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/RWL
rlabel locali 2942 -1504 2972 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/RWL
rlabel locali 3363 -1422 3378 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/WBL
rlabel locali 2973 -1422 2988 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/WBLb
rlabel locali 3436 -1568 3451 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/RBL0
rlabel locali 2899 -1568 2914 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/RBL1
rlabel metal1 3159 -1380 3191 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/VDD
rlabel metal1 3159 -1606 3191 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/GND
rlabel polycont 3121 -1499 3151 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/junc0
rlabel polycont 3199 -1499 3229 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/junc1
rlabel ndiff 2972 -1568 3028 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -1568 3378 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -1366 4611 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/WWL
rlabel locali 4538 -1504 4568 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/RWL
rlabel locali 4102 -1504 4132 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/RWL
rlabel locali 4523 -1422 4538 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/WBL
rlabel locali 4133 -1422 4148 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/WBLb
rlabel locali 4596 -1568 4611 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/RBL0
rlabel locali 4059 -1568 4074 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/RBL1
rlabel metal1 4319 -1380 4351 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/VDD
rlabel metal1 4319 -1606 4351 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/GND
rlabel polycont 4281 -1499 4311 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/junc0
rlabel polycont 4359 -1499 4389 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/junc1
rlabel ndiff 4132 -1568 4188 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -1568 4538 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -1366 4031 -1336 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/WWL
rlabel locali 3958 -1504 3988 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/RWL
rlabel locali 3522 -1504 3552 -1470 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/RWL
rlabel locali 3943 -1422 3958 -1393 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/WBL
rlabel locali 3553 -1422 3568 -1394 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/WBLb
rlabel locali 4016 -1568 4031 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/RBL0
rlabel locali 3479 -1568 3494 -1526 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/RBL1
rlabel metal1 3739 -1380 3771 -1366 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/VDD
rlabel metal1 3739 -1606 3771 -1592 7 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/GND
rlabel polycont 3701 -1499 3731 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/junc0
rlabel polycont 3779 -1499 3809 -1465 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/junc1
rlabel ndiff 3552 -1568 3608 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -1568 3958 -1540 1 10T_8x8_magic_1/10T_1x8_magic_7/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -1096 29 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/WWL
rlabel metal1 -1 -1234 14 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/RWL
rlabel corelocali 73 -1152 88 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_0
rlabel corelocali 463 -1152 478 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_0
rlabel corelocali -1 -1298 14 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_0
rlabel corelocali 536 -1298 551 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_0
rlabel corelocali 653 -1152 668 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_1
rlabel corelocali 1043 -1152 1058 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_1
rlabel corelocali 579 -1298 594 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_1
rlabel corelocali 1116 -1298 1131 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_1
rlabel corelocali 1233 -1152 1248 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_2
rlabel corelocali 1623 -1152 1638 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_2
rlabel corelocali 1159 -1298 1174 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_2
rlabel corelocali 1696 -1298 1711 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_2
rlabel corelocali 1813 -1152 1828 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_3
rlabel corelocali 2203 -1152 2218 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_3
rlabel corelocali 1739 -1298 1754 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_3
rlabel corelocali 2276 -1298 2291 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_3
rlabel corelocali 2393 -1152 2408 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_4
rlabel corelocali 2783 -1152 2798 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_4
rlabel corelocali 2319 -1298 2334 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_4
rlabel corelocali 2856 -1298 2871 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_4
rlabel corelocali 2973 -1152 2988 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_5
rlabel corelocali 3363 -1152 3378 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_5
rlabel corelocali 2899 -1298 2914 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_5
rlabel corelocali 3436 -1298 3451 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_5
rlabel corelocali 3553 -1152 3568 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_6
rlabel corelocali 3943 -1152 3958 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_6
rlabel corelocali 3479 -1298 3494 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_6
rlabel corelocali 4016 -1298 4031 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_6
rlabel corelocali 4133 -1152 4148 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/WBLb_7
rlabel corelocali 4523 -1152 4538 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/WBL_7
rlabel corelocali 4059 -1298 4074 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL1_7
rlabel corelocali 4596 -1298 4611 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/RBL0_7
rlabel metal1 -1 -1110 14 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/VDD
rlabel metal1 -1 -1336 14 -1322 1 10T_8x8_magic_1/10T_1x8_magic_6/GND
rlabel poly -1 -1096 551 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/WWL
rlabel locali 478 -1234 508 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/RWL
rlabel locali 42 -1234 72 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/RWL
rlabel locali 463 -1152 478 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/WBL
rlabel locali 73 -1152 88 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/WBLb
rlabel locali 536 -1298 551 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/RBL0
rlabel locali -1 -1298 14 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/RBL1
rlabel metal1 259 -1110 291 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/VDD
rlabel metal1 259 -1336 291 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/GND
rlabel polycont 221 -1229 251 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/junc0
rlabel polycont 299 -1229 329 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/junc1
rlabel ndiff 72 -1298 128 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -1298 478 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -1096 1131 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/WWL
rlabel locali 1058 -1234 1088 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/RWL
rlabel locali 622 -1234 652 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/RWL
rlabel locali 1043 -1152 1058 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/WBL
rlabel locali 653 -1152 668 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/WBLb
rlabel locali 1116 -1298 1131 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/RBL0
rlabel locali 579 -1298 594 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/RBL1
rlabel metal1 839 -1110 871 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/VDD
rlabel metal1 839 -1336 871 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/GND
rlabel polycont 801 -1229 831 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/junc0
rlabel polycont 879 -1229 909 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/junc1
rlabel ndiff 652 -1298 708 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -1298 1058 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -1096 1711 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/WWL
rlabel locali 1638 -1234 1668 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/RWL
rlabel locali 1202 -1234 1232 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/RWL
rlabel locali 1623 -1152 1638 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/WBL
rlabel locali 1233 -1152 1248 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/WBLb
rlabel locali 1696 -1298 1711 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/RBL0
rlabel locali 1159 -1298 1174 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/RBL1
rlabel metal1 1419 -1110 1451 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/VDD
rlabel metal1 1419 -1336 1451 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/GND
rlabel polycont 1381 -1229 1411 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/junc0
rlabel polycont 1459 -1229 1489 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/junc1
rlabel ndiff 1232 -1298 1288 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -1298 1638 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -1096 2291 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/WWL
rlabel locali 2218 -1234 2248 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/RWL
rlabel locali 1782 -1234 1812 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/RWL
rlabel locali 2203 -1152 2218 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/WBL
rlabel locali 1813 -1152 1828 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/WBLb
rlabel locali 2276 -1298 2291 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/RBL0
rlabel locali 1739 -1298 1754 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/RBL1
rlabel metal1 1999 -1110 2031 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/VDD
rlabel metal1 1999 -1336 2031 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/GND
rlabel polycont 1961 -1229 1991 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/junc0
rlabel polycont 2039 -1229 2069 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/junc1
rlabel ndiff 1812 -1298 1868 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -1298 2218 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -1096 2871 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/WWL
rlabel locali 2798 -1234 2828 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/RWL
rlabel locali 2362 -1234 2392 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/RWL
rlabel locali 2783 -1152 2798 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/WBL
rlabel locali 2393 -1152 2408 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/WBLb
rlabel locali 2856 -1298 2871 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/RBL0
rlabel locali 2319 -1298 2334 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/RBL1
rlabel metal1 2579 -1110 2611 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/VDD
rlabel metal1 2579 -1336 2611 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/GND
rlabel polycont 2541 -1229 2571 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/junc0
rlabel polycont 2619 -1229 2649 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/junc1
rlabel ndiff 2392 -1298 2448 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -1298 2798 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -1096 3451 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/WWL
rlabel locali 3378 -1234 3408 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/RWL
rlabel locali 2942 -1234 2972 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/RWL
rlabel locali 3363 -1152 3378 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/WBL
rlabel locali 2973 -1152 2988 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/WBLb
rlabel locali 3436 -1298 3451 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/RBL0
rlabel locali 2899 -1298 2914 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/RBL1
rlabel metal1 3159 -1110 3191 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/VDD
rlabel metal1 3159 -1336 3191 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/GND
rlabel polycont 3121 -1229 3151 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/junc0
rlabel polycont 3199 -1229 3229 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/junc1
rlabel ndiff 2972 -1298 3028 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -1298 3378 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -1096 4611 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/WWL
rlabel locali 4538 -1234 4568 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/RWL
rlabel locali 4102 -1234 4132 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/RWL
rlabel locali 4523 -1152 4538 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/WBL
rlabel locali 4133 -1152 4148 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/WBLb
rlabel locali 4596 -1298 4611 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/RBL0
rlabel locali 4059 -1298 4074 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/RBL1
rlabel metal1 4319 -1110 4351 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/VDD
rlabel metal1 4319 -1336 4351 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/GND
rlabel polycont 4281 -1229 4311 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/junc0
rlabel polycont 4359 -1229 4389 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/junc1
rlabel ndiff 4132 -1298 4188 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -1298 4538 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -1096 4031 -1066 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/WWL
rlabel locali 3958 -1234 3988 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/RWL
rlabel locali 3522 -1234 3552 -1200 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/RWL
rlabel locali 3943 -1152 3958 -1123 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/WBL
rlabel locali 3553 -1152 3568 -1124 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/WBLb
rlabel locali 4016 -1298 4031 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/RBL0
rlabel locali 3479 -1298 3494 -1256 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/RBL1
rlabel metal1 3739 -1110 3771 -1096 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/VDD
rlabel metal1 3739 -1336 3771 -1322 7 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/GND
rlabel polycont 3701 -1229 3731 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/junc0
rlabel polycont 3779 -1229 3809 -1195 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/junc1
rlabel ndiff 3552 -1298 3608 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -1298 3958 -1270 1 10T_8x8_magic_1/10T_1x8_magic_6/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -1636 29 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/WWL
rlabel metal1 -1 -1774 14 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/RWL
rlabel corelocali 73 -1692 88 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_0
rlabel corelocali 463 -1692 478 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_0
rlabel corelocali -1 -1838 14 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_0
rlabel corelocali 536 -1838 551 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_0
rlabel corelocali 653 -1692 668 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_1
rlabel corelocali 1043 -1692 1058 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_1
rlabel corelocali 579 -1838 594 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_1
rlabel corelocali 1116 -1838 1131 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_1
rlabel corelocali 1233 -1692 1248 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_2
rlabel corelocali 1623 -1692 1638 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_2
rlabel corelocali 1159 -1838 1174 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_2
rlabel corelocali 1696 -1838 1711 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_2
rlabel corelocali 1813 -1692 1828 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_3
rlabel corelocali 2203 -1692 2218 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_3
rlabel corelocali 1739 -1838 1754 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_3
rlabel corelocali 2276 -1838 2291 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_3
rlabel corelocali 2393 -1692 2408 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_4
rlabel corelocali 2783 -1692 2798 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_4
rlabel corelocali 2319 -1838 2334 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_4
rlabel corelocali 2856 -1838 2871 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_4
rlabel corelocali 2973 -1692 2988 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_5
rlabel corelocali 3363 -1692 3378 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_5
rlabel corelocali 2899 -1838 2914 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_5
rlabel corelocali 3436 -1838 3451 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_5
rlabel corelocali 3553 -1692 3568 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_6
rlabel corelocali 3943 -1692 3958 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_6
rlabel corelocali 3479 -1838 3494 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_6
rlabel corelocali 4016 -1838 4031 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_6
rlabel corelocali 4133 -1692 4148 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/WBLb_7
rlabel corelocali 4523 -1692 4538 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/WBL_7
rlabel corelocali 4059 -1838 4074 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL1_7
rlabel corelocali 4596 -1838 4611 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/RBL0_7
rlabel metal1 -1 -1650 14 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/VDD
rlabel metal1 -1 -1876 14 -1862 1 10T_8x8_magic_1/10T_1x8_magic_5/GND
rlabel poly -1 -1636 551 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/WWL
rlabel locali 478 -1774 508 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/RWL
rlabel locali 42 -1774 72 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/RWL
rlabel locali 463 -1692 478 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/WBL
rlabel locali 73 -1692 88 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/WBLb
rlabel locali 536 -1838 551 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/RBL0
rlabel locali -1 -1838 14 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/RBL1
rlabel metal1 259 -1650 291 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/VDD
rlabel metal1 259 -1876 291 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/GND
rlabel polycont 221 -1769 251 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/junc0
rlabel polycont 299 -1769 329 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/junc1
rlabel ndiff 72 -1838 128 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -1838 478 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -1636 1131 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/WWL
rlabel locali 1058 -1774 1088 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/RWL
rlabel locali 622 -1774 652 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/RWL
rlabel locali 1043 -1692 1058 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/WBL
rlabel locali 653 -1692 668 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/WBLb
rlabel locali 1116 -1838 1131 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/RBL0
rlabel locali 579 -1838 594 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/RBL1
rlabel metal1 839 -1650 871 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/VDD
rlabel metal1 839 -1876 871 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/GND
rlabel polycont 801 -1769 831 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/junc0
rlabel polycont 879 -1769 909 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/junc1
rlabel ndiff 652 -1838 708 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -1838 1058 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -1636 1711 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/WWL
rlabel locali 1638 -1774 1668 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/RWL
rlabel locali 1202 -1774 1232 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/RWL
rlabel locali 1623 -1692 1638 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/WBL
rlabel locali 1233 -1692 1248 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/WBLb
rlabel locali 1696 -1838 1711 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/RBL0
rlabel locali 1159 -1838 1174 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/RBL1
rlabel metal1 1419 -1650 1451 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/VDD
rlabel metal1 1419 -1876 1451 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/GND
rlabel polycont 1381 -1769 1411 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/junc0
rlabel polycont 1459 -1769 1489 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/junc1
rlabel ndiff 1232 -1838 1288 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -1838 1638 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -1636 2291 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/WWL
rlabel locali 2218 -1774 2248 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/RWL
rlabel locali 1782 -1774 1812 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/RWL
rlabel locali 2203 -1692 2218 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/WBL
rlabel locali 1813 -1692 1828 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/WBLb
rlabel locali 2276 -1838 2291 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/RBL0
rlabel locali 1739 -1838 1754 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/RBL1
rlabel metal1 1999 -1650 2031 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/VDD
rlabel metal1 1999 -1876 2031 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/GND
rlabel polycont 1961 -1769 1991 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/junc0
rlabel polycont 2039 -1769 2069 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/junc1
rlabel ndiff 1812 -1838 1868 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -1838 2218 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -1636 2871 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/WWL
rlabel locali 2798 -1774 2828 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/RWL
rlabel locali 2362 -1774 2392 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/RWL
rlabel locali 2783 -1692 2798 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/WBL
rlabel locali 2393 -1692 2408 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/WBLb
rlabel locali 2856 -1838 2871 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/RBL0
rlabel locali 2319 -1838 2334 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/RBL1
rlabel metal1 2579 -1650 2611 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/VDD
rlabel metal1 2579 -1876 2611 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/GND
rlabel polycont 2541 -1769 2571 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/junc0
rlabel polycont 2619 -1769 2649 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/junc1
rlabel ndiff 2392 -1838 2448 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -1838 2798 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -1636 3451 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/WWL
rlabel locali 3378 -1774 3408 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/RWL
rlabel locali 2942 -1774 2972 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/RWL
rlabel locali 3363 -1692 3378 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/WBL
rlabel locali 2973 -1692 2988 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/WBLb
rlabel locali 3436 -1838 3451 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/RBL0
rlabel locali 2899 -1838 2914 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/RBL1
rlabel metal1 3159 -1650 3191 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/VDD
rlabel metal1 3159 -1876 3191 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/GND
rlabel polycont 3121 -1769 3151 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/junc0
rlabel polycont 3199 -1769 3229 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/junc1
rlabel ndiff 2972 -1838 3028 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -1838 3378 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -1636 4611 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/WWL
rlabel locali 4538 -1774 4568 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/RWL
rlabel locali 4102 -1774 4132 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/RWL
rlabel locali 4523 -1692 4538 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/WBL
rlabel locali 4133 -1692 4148 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/WBLb
rlabel locali 4596 -1838 4611 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/RBL0
rlabel locali 4059 -1838 4074 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/RBL1
rlabel metal1 4319 -1650 4351 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/VDD
rlabel metal1 4319 -1876 4351 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/GND
rlabel polycont 4281 -1769 4311 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/junc0
rlabel polycont 4359 -1769 4389 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/junc1
rlabel ndiff 4132 -1838 4188 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -1838 4538 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -1636 4031 -1606 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/WWL
rlabel locali 3958 -1774 3988 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/RWL
rlabel locali 3522 -1774 3552 -1740 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/RWL
rlabel locali 3943 -1692 3958 -1663 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/WBL
rlabel locali 3553 -1692 3568 -1664 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/WBLb
rlabel locali 4016 -1838 4031 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/RBL0
rlabel locali 3479 -1838 3494 -1796 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/RBL1
rlabel metal1 3739 -1650 3771 -1636 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/VDD
rlabel metal1 3739 -1876 3771 -1862 7 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/GND
rlabel polycont 3701 -1769 3731 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/junc0
rlabel polycont 3779 -1769 3809 -1735 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/junc1
rlabel ndiff 3552 -1838 3608 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -1838 3958 -1810 1 10T_8x8_magic_1/10T_1x8_magic_5/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -1906 29 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/WWL
rlabel metal1 -1 -2044 14 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/RWL
rlabel corelocali 73 -1962 88 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_0
rlabel corelocali 463 -1962 478 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_0
rlabel corelocali -1 -2108 14 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_0
rlabel corelocali 536 -2108 551 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_0
rlabel corelocali 653 -1962 668 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_1
rlabel corelocali 1043 -1962 1058 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_1
rlabel corelocali 579 -2108 594 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_1
rlabel corelocali 1116 -2108 1131 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_1
rlabel corelocali 1233 -1962 1248 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_2
rlabel corelocali 1623 -1962 1638 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_2
rlabel corelocali 1159 -2108 1174 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_2
rlabel corelocali 1696 -2108 1711 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_2
rlabel corelocali 1813 -1962 1828 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_3
rlabel corelocali 2203 -1962 2218 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_3
rlabel corelocali 1739 -2108 1754 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_3
rlabel corelocali 2276 -2108 2291 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_3
rlabel corelocali 2393 -1962 2408 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_4
rlabel corelocali 2783 -1962 2798 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_4
rlabel corelocali 2319 -2108 2334 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_4
rlabel corelocali 2856 -2108 2871 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_4
rlabel corelocali 2973 -1962 2988 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_5
rlabel corelocali 3363 -1962 3378 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_5
rlabel corelocali 2899 -2108 2914 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_5
rlabel corelocali 3436 -2108 3451 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_5
rlabel corelocali 3553 -1962 3568 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_6
rlabel corelocali 3943 -1962 3958 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_6
rlabel corelocali 3479 -2108 3494 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_6
rlabel corelocali 4016 -2108 4031 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_6
rlabel corelocali 4133 -1962 4148 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/WBLb_7
rlabel corelocali 4523 -1962 4538 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/WBL_7
rlabel corelocali 4059 -2108 4074 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL1_7
rlabel corelocali 4596 -2108 4611 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/RBL0_7
rlabel metal1 -1 -1920 14 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/VDD
rlabel metal1 -1 -2146 14 -2132 1 10T_8x8_magic_1/10T_1x8_magic_4/GND
rlabel poly -1 -1906 551 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/WWL
rlabel locali 478 -2044 508 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/RWL
rlabel locali 42 -2044 72 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/RWL
rlabel locali 463 -1962 478 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/WBL
rlabel locali 73 -1962 88 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/WBLb
rlabel locali 536 -2108 551 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/RBL0
rlabel locali -1 -2108 14 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/RBL1
rlabel metal1 259 -1920 291 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/VDD
rlabel metal1 259 -2146 291 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/GND
rlabel polycont 221 -2039 251 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/junc0
rlabel polycont 299 -2039 329 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/junc1
rlabel ndiff 72 -2108 128 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -2108 478 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -1906 1131 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/WWL
rlabel locali 1058 -2044 1088 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/RWL
rlabel locali 622 -2044 652 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/RWL
rlabel locali 1043 -1962 1058 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/WBL
rlabel locali 653 -1962 668 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/WBLb
rlabel locali 1116 -2108 1131 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/RBL0
rlabel locali 579 -2108 594 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/RBL1
rlabel metal1 839 -1920 871 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/VDD
rlabel metal1 839 -2146 871 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/GND
rlabel polycont 801 -2039 831 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/junc0
rlabel polycont 879 -2039 909 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/junc1
rlabel ndiff 652 -2108 708 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -2108 1058 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -1906 1711 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/WWL
rlabel locali 1638 -2044 1668 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/RWL
rlabel locali 1202 -2044 1232 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/RWL
rlabel locali 1623 -1962 1638 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/WBL
rlabel locali 1233 -1962 1248 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/WBLb
rlabel locali 1696 -2108 1711 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/RBL0
rlabel locali 1159 -2108 1174 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/RBL1
rlabel metal1 1419 -1920 1451 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/VDD
rlabel metal1 1419 -2146 1451 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/GND
rlabel polycont 1381 -2039 1411 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/junc0
rlabel polycont 1459 -2039 1489 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/junc1
rlabel ndiff 1232 -2108 1288 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -2108 1638 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -1906 2291 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/WWL
rlabel locali 2218 -2044 2248 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/RWL
rlabel locali 1782 -2044 1812 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/RWL
rlabel locali 2203 -1962 2218 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/WBL
rlabel locali 1813 -1962 1828 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/WBLb
rlabel locali 2276 -2108 2291 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/RBL0
rlabel locali 1739 -2108 1754 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/RBL1
rlabel metal1 1999 -1920 2031 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/VDD
rlabel metal1 1999 -2146 2031 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/GND
rlabel polycont 1961 -2039 1991 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/junc0
rlabel polycont 2039 -2039 2069 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/junc1
rlabel ndiff 1812 -2108 1868 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -2108 2218 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -1906 2871 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/WWL
rlabel locali 2798 -2044 2828 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/RWL
rlabel locali 2362 -2044 2392 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/RWL
rlabel locali 2783 -1962 2798 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/WBL
rlabel locali 2393 -1962 2408 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/WBLb
rlabel locali 2856 -2108 2871 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/RBL0
rlabel locali 2319 -2108 2334 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/RBL1
rlabel metal1 2579 -1920 2611 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/VDD
rlabel metal1 2579 -2146 2611 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/GND
rlabel polycont 2541 -2039 2571 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/junc0
rlabel polycont 2619 -2039 2649 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/junc1
rlabel ndiff 2392 -2108 2448 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -2108 2798 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -1906 3451 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/WWL
rlabel locali 3378 -2044 3408 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/RWL
rlabel locali 2942 -2044 2972 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/RWL
rlabel locali 3363 -1962 3378 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/WBL
rlabel locali 2973 -1962 2988 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/WBLb
rlabel locali 3436 -2108 3451 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/RBL0
rlabel locali 2899 -2108 2914 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/RBL1
rlabel metal1 3159 -1920 3191 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/VDD
rlabel metal1 3159 -2146 3191 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/GND
rlabel polycont 3121 -2039 3151 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/junc0
rlabel polycont 3199 -2039 3229 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/junc1
rlabel ndiff 2972 -2108 3028 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -2108 3378 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -1906 4611 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/WWL
rlabel locali 4538 -2044 4568 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/RWL
rlabel locali 4102 -2044 4132 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/RWL
rlabel locali 4523 -1962 4538 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/WBL
rlabel locali 4133 -1962 4148 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/WBLb
rlabel locali 4596 -2108 4611 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/RBL0
rlabel locali 4059 -2108 4074 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/RBL1
rlabel metal1 4319 -1920 4351 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/VDD
rlabel metal1 4319 -2146 4351 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/GND
rlabel polycont 4281 -2039 4311 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/junc0
rlabel polycont 4359 -2039 4389 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/junc1
rlabel ndiff 4132 -2108 4188 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -2108 4538 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -1906 4031 -1876 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/WWL
rlabel locali 3958 -2044 3988 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/RWL
rlabel locali 3522 -2044 3552 -2010 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/RWL
rlabel locali 3943 -1962 3958 -1933 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/WBL
rlabel locali 3553 -1962 3568 -1934 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/WBLb
rlabel locali 4016 -2108 4031 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/RBL0
rlabel locali 3479 -2108 3494 -2066 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/RBL1
rlabel metal1 3739 -1920 3771 -1906 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/VDD
rlabel metal1 3739 -2146 3771 -2132 7 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/GND
rlabel polycont 3701 -2039 3731 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/junc0
rlabel polycont 3779 -2039 3809 -2005 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/junc1
rlabel ndiff 3552 -2108 3608 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -2108 3958 -2080 1 10T_8x8_magic_1/10T_1x8_magic_4/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -286 29 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/WWL
rlabel metal1 -1 -424 14 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/RWL
rlabel corelocali 73 -342 88 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_0
rlabel corelocali 463 -342 478 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_0
rlabel corelocali -1 -488 14 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_0
rlabel corelocali 536 -488 551 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_0
rlabel corelocali 653 -342 668 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_1
rlabel corelocali 1043 -342 1058 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_1
rlabel corelocali 579 -488 594 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_1
rlabel corelocali 1116 -488 1131 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_1
rlabel corelocali 1233 -342 1248 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_2
rlabel corelocali 1623 -342 1638 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_2
rlabel corelocali 1159 -488 1174 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_2
rlabel corelocali 1696 -488 1711 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_2
rlabel corelocali 1813 -342 1828 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_3
rlabel corelocali 2203 -342 2218 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_3
rlabel corelocali 1739 -488 1754 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_3
rlabel corelocali 2276 -488 2291 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_3
rlabel corelocali 2393 -342 2408 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_4
rlabel corelocali 2783 -342 2798 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_4
rlabel corelocali 2319 -488 2334 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_4
rlabel corelocali 2856 -488 2871 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_4
rlabel corelocali 2973 -342 2988 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_5
rlabel corelocali 3363 -342 3378 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_5
rlabel corelocali 2899 -488 2914 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_5
rlabel corelocali 3436 -488 3451 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_5
rlabel corelocali 3553 -342 3568 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_6
rlabel corelocali 3943 -342 3958 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_6
rlabel corelocali 3479 -488 3494 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_6
rlabel corelocali 4016 -488 4031 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_6
rlabel corelocali 4133 -342 4148 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/WBLb_7
rlabel corelocali 4523 -342 4538 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/WBL_7
rlabel corelocali 4059 -488 4074 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL1_7
rlabel corelocali 4596 -488 4611 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/RBL0_7
rlabel metal1 -1 -300 14 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/VDD
rlabel metal1 -1 -526 14 -512 1 10T_8x8_magic_1/10T_1x8_magic_3/GND
rlabel poly -1 -286 551 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/WWL
rlabel locali 478 -424 508 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/RWL
rlabel locali 42 -424 72 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/RWL
rlabel locali 463 -342 478 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/WBL
rlabel locali 73 -342 88 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/WBLb
rlabel locali 536 -488 551 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/RBL0
rlabel locali -1 -488 14 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/RBL1
rlabel metal1 259 -300 291 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/VDD
rlabel metal1 259 -526 291 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/GND
rlabel polycont 221 -419 251 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/junc0
rlabel polycont 299 -419 329 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/junc1
rlabel ndiff 72 -488 128 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -488 478 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -286 1131 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/WWL
rlabel locali 1058 -424 1088 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/RWL
rlabel locali 622 -424 652 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/RWL
rlabel locali 1043 -342 1058 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/WBL
rlabel locali 653 -342 668 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/WBLb
rlabel locali 1116 -488 1131 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/RBL0
rlabel locali 579 -488 594 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/RBL1
rlabel metal1 839 -300 871 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/VDD
rlabel metal1 839 -526 871 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/GND
rlabel polycont 801 -419 831 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/junc0
rlabel polycont 879 -419 909 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/junc1
rlabel ndiff 652 -488 708 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -488 1058 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -286 1711 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/WWL
rlabel locali 1638 -424 1668 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/RWL
rlabel locali 1202 -424 1232 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/RWL
rlabel locali 1623 -342 1638 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/WBL
rlabel locali 1233 -342 1248 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/WBLb
rlabel locali 1696 -488 1711 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/RBL0
rlabel locali 1159 -488 1174 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/RBL1
rlabel metal1 1419 -300 1451 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/VDD
rlabel metal1 1419 -526 1451 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/GND
rlabel polycont 1381 -419 1411 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/junc0
rlabel polycont 1459 -419 1489 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/junc1
rlabel ndiff 1232 -488 1288 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -488 1638 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -286 2291 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/WWL
rlabel locali 2218 -424 2248 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/RWL
rlabel locali 1782 -424 1812 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/RWL
rlabel locali 2203 -342 2218 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/WBL
rlabel locali 1813 -342 1828 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/WBLb
rlabel locali 2276 -488 2291 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/RBL0
rlabel locali 1739 -488 1754 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/RBL1
rlabel metal1 1999 -300 2031 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/VDD
rlabel metal1 1999 -526 2031 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/GND
rlabel polycont 1961 -419 1991 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/junc0
rlabel polycont 2039 -419 2069 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/junc1
rlabel ndiff 1812 -488 1868 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -488 2218 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -286 2871 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/WWL
rlabel locali 2798 -424 2828 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/RWL
rlabel locali 2362 -424 2392 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/RWL
rlabel locali 2783 -342 2798 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/WBL
rlabel locali 2393 -342 2408 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/WBLb
rlabel locali 2856 -488 2871 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/RBL0
rlabel locali 2319 -488 2334 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/RBL1
rlabel metal1 2579 -300 2611 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/VDD
rlabel metal1 2579 -526 2611 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/GND
rlabel polycont 2541 -419 2571 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/junc0
rlabel polycont 2619 -419 2649 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/junc1
rlabel ndiff 2392 -488 2448 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -488 2798 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -286 3451 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/WWL
rlabel locali 3378 -424 3408 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/RWL
rlabel locali 2942 -424 2972 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/RWL
rlabel locali 3363 -342 3378 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/WBL
rlabel locali 2973 -342 2988 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/WBLb
rlabel locali 3436 -488 3451 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/RBL0
rlabel locali 2899 -488 2914 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/RBL1
rlabel metal1 3159 -300 3191 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/VDD
rlabel metal1 3159 -526 3191 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/GND
rlabel polycont 3121 -419 3151 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/junc0
rlabel polycont 3199 -419 3229 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/junc1
rlabel ndiff 2972 -488 3028 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -488 3378 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -286 4611 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/WWL
rlabel locali 4538 -424 4568 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/RWL
rlabel locali 4102 -424 4132 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/RWL
rlabel locali 4523 -342 4538 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/WBL
rlabel locali 4133 -342 4148 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/WBLb
rlabel locali 4596 -488 4611 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/RBL0
rlabel locali 4059 -488 4074 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/RBL1
rlabel metal1 4319 -300 4351 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/VDD
rlabel metal1 4319 -526 4351 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/GND
rlabel polycont 4281 -419 4311 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/junc0
rlabel polycont 4359 -419 4389 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/junc1
rlabel ndiff 4132 -488 4188 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -488 4538 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -286 4031 -256 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/WWL
rlabel locali 3958 -424 3988 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/RWL
rlabel locali 3522 -424 3552 -390 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/RWL
rlabel locali 3943 -342 3958 -313 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/WBL
rlabel locali 3553 -342 3568 -314 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/WBLb
rlabel locali 4016 -488 4031 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/RBL0
rlabel locali 3479 -488 3494 -446 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/RBL1
rlabel metal1 3739 -300 3771 -286 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/VDD
rlabel metal1 3739 -526 3771 -512 7 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/GND
rlabel polycont 3701 -419 3731 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/junc0
rlabel polycont 3779 -419 3809 -385 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/junc1
rlabel ndiff 3552 -488 3608 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -488 3958 -460 1 10T_8x8_magic_1/10T_1x8_magic_3/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -16 29 14 1 10T_8x8_magic_1/10T_1x8_magic_2/WWL
rlabel metal1 -1 -154 14 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/RWL
rlabel corelocali 73 -72 88 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_0
rlabel corelocali 463 -72 478 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_0
rlabel corelocali -1 -218 14 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_0
rlabel corelocali 536 -218 551 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_0
rlabel corelocali 653 -72 668 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_1
rlabel corelocali 1043 -72 1058 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_1
rlabel corelocali 579 -218 594 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_1
rlabel corelocali 1116 -218 1131 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_1
rlabel corelocali 1233 -72 1248 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_2
rlabel corelocali 1623 -72 1638 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_2
rlabel corelocali 1159 -218 1174 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_2
rlabel corelocali 1696 -218 1711 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_2
rlabel corelocali 1813 -72 1828 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_3
rlabel corelocali 2203 -72 2218 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_3
rlabel corelocali 1739 -218 1754 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_3
rlabel corelocali 2276 -218 2291 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_3
rlabel corelocali 2393 -72 2408 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_4
rlabel corelocali 2783 -72 2798 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_4
rlabel corelocali 2319 -218 2334 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_4
rlabel corelocali 2856 -218 2871 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_4
rlabel corelocali 2973 -72 2988 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_5
rlabel corelocali 3363 -72 3378 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_5
rlabel corelocali 2899 -218 2914 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_5
rlabel corelocali 3436 -218 3451 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_5
rlabel corelocali 3553 -72 3568 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_6
rlabel corelocali 3943 -72 3958 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_6
rlabel corelocali 3479 -218 3494 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_6
rlabel corelocali 4016 -218 4031 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_6
rlabel corelocali 4133 -72 4148 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/WBLb_7
rlabel corelocali 4523 -72 4538 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/WBL_7
rlabel corelocali 4059 -218 4074 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL1_7
rlabel corelocali 4596 -218 4611 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/RBL0_7
rlabel metal1 -1 -30 14 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/VDD
rlabel metal1 -1 -256 14 -242 1 10T_8x8_magic_1/10T_1x8_magic_2/GND
rlabel poly -1 -16 551 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/WWL
rlabel locali 478 -154 508 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/RWL
rlabel locali 42 -154 72 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/RWL
rlabel locali 463 -72 478 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/WBL
rlabel locali 73 -72 88 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/WBLb
rlabel locali 536 -218 551 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/RBL0
rlabel locali -1 -218 14 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/RBL1
rlabel metal1 259 -30 291 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/VDD
rlabel metal1 259 -256 291 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/GND
rlabel polycont 221 -149 251 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/junc0
rlabel polycont 299 -149 329 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/junc1
rlabel ndiff 72 -218 128 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -218 478 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -16 1131 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/WWL
rlabel locali 1058 -154 1088 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/RWL
rlabel locali 622 -154 652 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/RWL
rlabel locali 1043 -72 1058 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/WBL
rlabel locali 653 -72 668 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/WBLb
rlabel locali 1116 -218 1131 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/RBL0
rlabel locali 579 -218 594 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/RBL1
rlabel metal1 839 -30 871 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/VDD
rlabel metal1 839 -256 871 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/GND
rlabel polycont 801 -149 831 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/junc0
rlabel polycont 879 -149 909 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/junc1
rlabel ndiff 652 -218 708 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -218 1058 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -16 1711 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/WWL
rlabel locali 1638 -154 1668 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/RWL
rlabel locali 1202 -154 1232 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/RWL
rlabel locali 1623 -72 1638 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/WBL
rlabel locali 1233 -72 1248 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/WBLb
rlabel locali 1696 -218 1711 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/RBL0
rlabel locali 1159 -218 1174 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/RBL1
rlabel metal1 1419 -30 1451 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/VDD
rlabel metal1 1419 -256 1451 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/GND
rlabel polycont 1381 -149 1411 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/junc0
rlabel polycont 1459 -149 1489 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/junc1
rlabel ndiff 1232 -218 1288 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -218 1638 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -16 2291 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/WWL
rlabel locali 2218 -154 2248 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/RWL
rlabel locali 1782 -154 1812 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/RWL
rlabel locali 2203 -72 2218 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/WBL
rlabel locali 1813 -72 1828 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/WBLb
rlabel locali 2276 -218 2291 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/RBL0
rlabel locali 1739 -218 1754 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/RBL1
rlabel metal1 1999 -30 2031 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/VDD
rlabel metal1 1999 -256 2031 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/GND
rlabel polycont 1961 -149 1991 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/junc0
rlabel polycont 2039 -149 2069 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/junc1
rlabel ndiff 1812 -218 1868 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -218 2218 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -16 2871 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/WWL
rlabel locali 2798 -154 2828 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/RWL
rlabel locali 2362 -154 2392 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/RWL
rlabel locali 2783 -72 2798 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/WBL
rlabel locali 2393 -72 2408 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/WBLb
rlabel locali 2856 -218 2871 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/RBL0
rlabel locali 2319 -218 2334 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/RBL1
rlabel metal1 2579 -30 2611 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/VDD
rlabel metal1 2579 -256 2611 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/GND
rlabel polycont 2541 -149 2571 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/junc0
rlabel polycont 2619 -149 2649 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/junc1
rlabel ndiff 2392 -218 2448 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -218 2798 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -16 3451 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/WWL
rlabel locali 3378 -154 3408 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/RWL
rlabel locali 2942 -154 2972 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/RWL
rlabel locali 3363 -72 3378 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/WBL
rlabel locali 2973 -72 2988 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/WBLb
rlabel locali 3436 -218 3451 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/RBL0
rlabel locali 2899 -218 2914 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/RBL1
rlabel metal1 3159 -30 3191 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/VDD
rlabel metal1 3159 -256 3191 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/GND
rlabel polycont 3121 -149 3151 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/junc0
rlabel polycont 3199 -149 3229 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/junc1
rlabel ndiff 2972 -218 3028 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -218 3378 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -16 4611 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/WWL
rlabel locali 4538 -154 4568 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/RWL
rlabel locali 4102 -154 4132 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/RWL
rlabel locali 4523 -72 4538 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/WBL
rlabel locali 4133 -72 4148 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/WBLb
rlabel locali 4596 -218 4611 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/RBL0
rlabel locali 4059 -218 4074 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/RBL1
rlabel metal1 4319 -30 4351 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/VDD
rlabel metal1 4319 -256 4351 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/GND
rlabel polycont 4281 -149 4311 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/junc0
rlabel polycont 4359 -149 4389 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/junc1
rlabel ndiff 4132 -218 4188 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -218 4538 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -16 4031 14 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/WWL
rlabel locali 3958 -154 3988 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/RWL
rlabel locali 3522 -154 3552 -120 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/RWL
rlabel locali 3943 -72 3958 -43 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/WBL
rlabel locali 3553 -72 3568 -44 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/WBLb
rlabel locali 4016 -218 4031 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/RBL0
rlabel locali 3479 -218 3494 -176 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/RBL1
rlabel metal1 3739 -30 3771 -16 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/VDD
rlabel metal1 3739 -256 3771 -242 7 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/GND
rlabel polycont 3701 -149 3731 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/junc0
rlabel polycont 3779 -149 3809 -115 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/junc1
rlabel ndiff 3552 -218 3608 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -218 3958 -190 1 10T_8x8_magic_1/10T_1x8_magic_2/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -826 29 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/WWL
rlabel metal1 -1 -964 14 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/RWL
rlabel corelocali 73 -882 88 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_0
rlabel corelocali 463 -882 478 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_0
rlabel corelocali -1 -1028 14 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_0
rlabel corelocali 536 -1028 551 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_0
rlabel corelocali 653 -882 668 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_1
rlabel corelocali 1043 -882 1058 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_1
rlabel corelocali 579 -1028 594 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_1
rlabel corelocali 1116 -1028 1131 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_1
rlabel corelocali 1233 -882 1248 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_2
rlabel corelocali 1623 -882 1638 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_2
rlabel corelocali 1159 -1028 1174 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_2
rlabel corelocali 1696 -1028 1711 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_2
rlabel corelocali 1813 -882 1828 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_3
rlabel corelocali 2203 -882 2218 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_3
rlabel corelocali 1739 -1028 1754 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_3
rlabel corelocali 2276 -1028 2291 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_3
rlabel corelocali 2393 -882 2408 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_4
rlabel corelocali 2783 -882 2798 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_4
rlabel corelocali 2319 -1028 2334 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_4
rlabel corelocali 2856 -1028 2871 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_4
rlabel corelocali 2973 -882 2988 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_5
rlabel corelocali 3363 -882 3378 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_5
rlabel corelocali 2899 -1028 2914 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_5
rlabel corelocali 3436 -1028 3451 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_5
rlabel corelocali 3553 -882 3568 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_6
rlabel corelocali 3943 -882 3958 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_6
rlabel corelocali 3479 -1028 3494 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_6
rlabel corelocali 4016 -1028 4031 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_6
rlabel corelocali 4133 -882 4148 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/WBLb_7
rlabel corelocali 4523 -882 4538 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/WBL_7
rlabel corelocali 4059 -1028 4074 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL1_7
rlabel corelocali 4596 -1028 4611 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/RBL0_7
rlabel metal1 -1 -840 14 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/VDD
rlabel metal1 -1 -1066 14 -1052 1 10T_8x8_magic_1/10T_1x8_magic_1/GND
rlabel poly -1 -826 551 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/WWL
rlabel locali 478 -964 508 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/RWL
rlabel locali 42 -964 72 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/RWL
rlabel locali 463 -882 478 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/WBL
rlabel locali 73 -882 88 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/WBLb
rlabel locali 536 -1028 551 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/RBL0
rlabel locali -1 -1028 14 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/RBL1
rlabel metal1 259 -840 291 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/VDD
rlabel metal1 259 -1066 291 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/GND
rlabel polycont 221 -959 251 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/junc0
rlabel polycont 299 -959 329 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/junc1
rlabel ndiff 72 -1028 128 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -1028 478 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -826 1131 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/WWL
rlabel locali 1058 -964 1088 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/RWL
rlabel locali 622 -964 652 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/RWL
rlabel locali 1043 -882 1058 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/WBL
rlabel locali 653 -882 668 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/WBLb
rlabel locali 1116 -1028 1131 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/RBL0
rlabel locali 579 -1028 594 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/RBL1
rlabel metal1 839 -840 871 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/VDD
rlabel metal1 839 -1066 871 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/GND
rlabel polycont 801 -959 831 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/junc0
rlabel polycont 879 -959 909 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/junc1
rlabel ndiff 652 -1028 708 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -1028 1058 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -826 1711 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/WWL
rlabel locali 1638 -964 1668 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/RWL
rlabel locali 1202 -964 1232 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/RWL
rlabel locali 1623 -882 1638 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/WBL
rlabel locali 1233 -882 1248 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/WBLb
rlabel locali 1696 -1028 1711 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/RBL0
rlabel locali 1159 -1028 1174 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/RBL1
rlabel metal1 1419 -840 1451 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/VDD
rlabel metal1 1419 -1066 1451 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/GND
rlabel polycont 1381 -959 1411 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/junc0
rlabel polycont 1459 -959 1489 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/junc1
rlabel ndiff 1232 -1028 1288 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -1028 1638 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -826 2291 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/WWL
rlabel locali 2218 -964 2248 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/RWL
rlabel locali 1782 -964 1812 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/RWL
rlabel locali 2203 -882 2218 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/WBL
rlabel locali 1813 -882 1828 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/WBLb
rlabel locali 2276 -1028 2291 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/RBL0
rlabel locali 1739 -1028 1754 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/RBL1
rlabel metal1 1999 -840 2031 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/VDD
rlabel metal1 1999 -1066 2031 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/GND
rlabel polycont 1961 -959 1991 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/junc0
rlabel polycont 2039 -959 2069 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/junc1
rlabel ndiff 1812 -1028 1868 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -1028 2218 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -826 2871 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/WWL
rlabel locali 2798 -964 2828 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/RWL
rlabel locali 2362 -964 2392 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/RWL
rlabel locali 2783 -882 2798 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/WBL
rlabel locali 2393 -882 2408 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/WBLb
rlabel locali 2856 -1028 2871 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/RBL0
rlabel locali 2319 -1028 2334 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/RBL1
rlabel metal1 2579 -840 2611 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/VDD
rlabel metal1 2579 -1066 2611 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/GND
rlabel polycont 2541 -959 2571 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/junc0
rlabel polycont 2619 -959 2649 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/junc1
rlabel ndiff 2392 -1028 2448 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -1028 2798 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -826 3451 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/WWL
rlabel locali 3378 -964 3408 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/RWL
rlabel locali 2942 -964 2972 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/RWL
rlabel locali 3363 -882 3378 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/WBL
rlabel locali 2973 -882 2988 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/WBLb
rlabel locali 3436 -1028 3451 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/RBL0
rlabel locali 2899 -1028 2914 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/RBL1
rlabel metal1 3159 -840 3191 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/VDD
rlabel metal1 3159 -1066 3191 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/GND
rlabel polycont 3121 -959 3151 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/junc0
rlabel polycont 3199 -959 3229 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/junc1
rlabel ndiff 2972 -1028 3028 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -1028 3378 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -826 4611 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/WWL
rlabel locali 4538 -964 4568 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/RWL
rlabel locali 4102 -964 4132 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/RWL
rlabel locali 4523 -882 4538 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/WBL
rlabel locali 4133 -882 4148 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/WBLb
rlabel locali 4596 -1028 4611 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/RBL0
rlabel locali 4059 -1028 4074 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/RBL1
rlabel metal1 4319 -840 4351 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/VDD
rlabel metal1 4319 -1066 4351 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/GND
rlabel polycont 4281 -959 4311 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/junc0
rlabel polycont 4359 -959 4389 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/junc1
rlabel ndiff 4132 -1028 4188 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -1028 4538 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -826 4031 -796 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/WWL
rlabel locali 3958 -964 3988 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/RWL
rlabel locali 3522 -964 3552 -930 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/RWL
rlabel locali 3943 -882 3958 -853 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/WBL
rlabel locali 3553 -882 3568 -854 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/WBLb
rlabel locali 4016 -1028 4031 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/RBL0
rlabel locali 3479 -1028 3494 -986 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/RBL1
rlabel metal1 3739 -840 3771 -826 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/VDD
rlabel metal1 3739 -1066 3771 -1052 7 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/GND
rlabel polycont 3701 -959 3731 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/junc0
rlabel polycont 3779 -959 3809 -925 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/junc1
rlabel ndiff 3552 -1028 3608 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -1028 3958 -1000 1 10T_8x8_magic_1/10T_1x8_magic_1/10T_toy_magic_0/RWL0_junc
rlabel poly -1 -556 29 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/WWL
rlabel metal1 -1 -694 14 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/RWL
rlabel corelocali 73 -612 88 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_0
rlabel corelocali 463 -612 478 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_0
rlabel corelocali -1 -758 14 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_0
rlabel corelocali 536 -758 551 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_0
rlabel corelocali 653 -612 668 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_1
rlabel corelocali 1043 -612 1058 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_1
rlabel corelocali 579 -758 594 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_1
rlabel corelocali 1116 -758 1131 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_1
rlabel corelocali 1233 -612 1248 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_2
rlabel corelocali 1623 -612 1638 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_2
rlabel corelocali 1159 -758 1174 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_2
rlabel corelocali 1696 -758 1711 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_2
rlabel corelocali 1813 -612 1828 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_3
rlabel corelocali 2203 -612 2218 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_3
rlabel corelocali 1739 -758 1754 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_3
rlabel corelocali 2276 -758 2291 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_3
rlabel corelocali 2393 -612 2408 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_4
rlabel corelocali 2783 -612 2798 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_4
rlabel corelocali 2319 -758 2334 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_4
rlabel corelocali 2856 -758 2871 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_4
rlabel corelocali 2973 -612 2988 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_5
rlabel corelocali 3363 -612 3378 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_5
rlabel corelocali 2899 -758 2914 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_5
rlabel corelocali 3436 -758 3451 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_5
rlabel corelocali 3553 -612 3568 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_6
rlabel corelocali 3943 -612 3958 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_6
rlabel corelocali 3479 -758 3494 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_6
rlabel corelocali 4016 -758 4031 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_6
rlabel corelocali 4133 -612 4148 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/WBLb_7
rlabel corelocali 4523 -612 4538 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/WBL_7
rlabel corelocali 4059 -758 4074 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL1_7
rlabel corelocali 4596 -758 4611 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/RBL0_7
rlabel metal1 -1 -570 14 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/VDD
rlabel metal1 -1 -796 14 -782 1 10T_8x8_magic_1/10T_1x8_magic_0/GND
rlabel poly -1 -556 551 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/WWL
rlabel locali 478 -694 508 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/RWL
rlabel locali 42 -694 72 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/RWL
rlabel locali 463 -612 478 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/WBL
rlabel locali 73 -612 88 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/WBLb
rlabel locali 536 -758 551 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/RBL0
rlabel locali -1 -758 14 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/RBL1
rlabel metal1 259 -570 291 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/VDD
rlabel metal1 259 -796 291 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/GND
rlabel polycont 221 -689 251 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/junc0
rlabel polycont 299 -689 329 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/junc1
rlabel ndiff 72 -758 128 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/RWL1_junc
rlabel ndiff 422 -758 478 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_7/RWL0_junc
rlabel poly 579 -556 1131 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/WWL
rlabel locali 1058 -694 1088 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/RWL
rlabel locali 622 -694 652 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/RWL
rlabel locali 1043 -612 1058 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/WBL
rlabel locali 653 -612 668 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/WBLb
rlabel locali 1116 -758 1131 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/RBL0
rlabel locali 579 -758 594 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/RBL1
rlabel metal1 839 -570 871 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/VDD
rlabel metal1 839 -796 871 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/GND
rlabel polycont 801 -689 831 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/junc0
rlabel polycont 879 -689 909 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/junc1
rlabel ndiff 652 -758 708 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/RWL1_junc
rlabel ndiff 1002 -758 1058 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_6/RWL0_junc
rlabel poly 1159 -556 1711 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/WWL
rlabel locali 1638 -694 1668 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/RWL
rlabel locali 1202 -694 1232 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/RWL
rlabel locali 1623 -612 1638 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/WBL
rlabel locali 1233 -612 1248 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/WBLb
rlabel locali 1696 -758 1711 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/RBL0
rlabel locali 1159 -758 1174 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/RBL1
rlabel metal1 1419 -570 1451 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/VDD
rlabel metal1 1419 -796 1451 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/GND
rlabel polycont 1381 -689 1411 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/junc0
rlabel polycont 1459 -689 1489 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/junc1
rlabel ndiff 1232 -758 1288 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/RWL1_junc
rlabel ndiff 1582 -758 1638 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_5/RWL0_junc
rlabel poly 1739 -556 2291 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/WWL
rlabel locali 2218 -694 2248 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/RWL
rlabel locali 1782 -694 1812 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/RWL
rlabel locali 2203 -612 2218 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/WBL
rlabel locali 1813 -612 1828 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/WBLb
rlabel locali 2276 -758 2291 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/RBL0
rlabel locali 1739 -758 1754 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/RBL1
rlabel metal1 1999 -570 2031 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/VDD
rlabel metal1 1999 -796 2031 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/GND
rlabel polycont 1961 -689 1991 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/junc0
rlabel polycont 2039 -689 2069 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/junc1
rlabel ndiff 1812 -758 1868 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/RWL1_junc
rlabel ndiff 2162 -758 2218 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_4/RWL0_junc
rlabel poly 2319 -556 2871 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/WWL
rlabel locali 2798 -694 2828 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/RWL
rlabel locali 2362 -694 2392 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/RWL
rlabel locali 2783 -612 2798 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/WBL
rlabel locali 2393 -612 2408 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/WBLb
rlabel locali 2856 -758 2871 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/RBL0
rlabel locali 2319 -758 2334 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/RBL1
rlabel metal1 2579 -570 2611 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/VDD
rlabel metal1 2579 -796 2611 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/GND
rlabel polycont 2541 -689 2571 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/junc0
rlabel polycont 2619 -689 2649 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/junc1
rlabel ndiff 2392 -758 2448 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/RWL1_junc
rlabel ndiff 2742 -758 2798 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_3/RWL0_junc
rlabel poly 2899 -556 3451 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/WWL
rlabel locali 3378 -694 3408 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/RWL
rlabel locali 2942 -694 2972 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/RWL
rlabel locali 3363 -612 3378 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/WBL
rlabel locali 2973 -612 2988 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/WBLb
rlabel locali 3436 -758 3451 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/RBL0
rlabel locali 2899 -758 2914 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/RBL1
rlabel metal1 3159 -570 3191 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/VDD
rlabel metal1 3159 -796 3191 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/GND
rlabel polycont 3121 -689 3151 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/junc0
rlabel polycont 3199 -689 3229 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/junc1
rlabel ndiff 2972 -758 3028 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/RWL1_junc
rlabel ndiff 3322 -758 3378 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_2/RWL0_junc
rlabel poly 4059 -556 4611 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/WWL
rlabel locali 4538 -694 4568 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/RWL
rlabel locali 4102 -694 4132 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/RWL
rlabel locali 4523 -612 4538 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/WBL
rlabel locali 4133 -612 4148 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/WBLb
rlabel locali 4596 -758 4611 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/RBL0
rlabel locali 4059 -758 4074 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/RBL1
rlabel metal1 4319 -570 4351 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/VDD
rlabel metal1 4319 -796 4351 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/GND
rlabel polycont 4281 -689 4311 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/junc0
rlabel polycont 4359 -689 4389 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/junc1
rlabel ndiff 4132 -758 4188 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/RWL1_junc
rlabel ndiff 4482 -758 4538 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_1/RWL0_junc
rlabel poly 3479 -556 4031 -526 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/WWL
rlabel locali 3958 -694 3988 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/RWL
rlabel locali 3522 -694 3552 -660 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/RWL
rlabel locali 3943 -612 3958 -583 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/WBL
rlabel locali 3553 -612 3568 -584 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/WBLb
rlabel locali 4016 -758 4031 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/RBL0
rlabel locali 3479 -758 3494 -716 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/RBL1
rlabel metal1 3739 -570 3771 -556 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/VDD
rlabel metal1 3739 -796 3771 -782 7 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/GND
rlabel polycont 3701 -689 3731 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/junc0
rlabel polycont 3779 -689 3809 -655 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/junc1
rlabel ndiff 3552 -758 3608 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/RWL1_junc
rlabel ndiff 3902 -758 3958 -730 1 10T_8x8_magic_1/10T_1x8_magic_0/10T_toy_magic_0/RWL0_junc
rlabel poly 4591 1063 4621 1093 1 10T_4x4_magic_0/WWL_0
rlabel poly 4591 793 4621 823 1 10T_4x4_magic_0/WWL_1
rlabel metal1 4591 1049 4621 1063 1 10T_4x4_magic_0/VDD
rlabel metal1 4591 779 4621 793 1 10T_4x4_magic_0/VDD
rlabel metal1 4591 823 4621 837 1 10T_4x4_magic_0/GND
rlabel metal1 4591 553 4621 567 1 10T_4x4_magic_0/GND
rlabel corelocali 4639 505 4654 535 1 10T_4x4_magic_0/RBL1_0
rlabel corelocali 5176 505 5191 535 1 10T_4x4_magic_0/RBL0_0
rlabel corelocali 5219 505 5234 535 1 10T_4x4_magic_0/RBL1_1
rlabel corelocali 5756 505 5771 535 1 10T_4x4_magic_0/RBL0_1
rlabel metal1 4591 655 4621 689 1 10T_4x4_magic_0/RWL_1
rlabel metal1 4591 925 4621 959 1 10T_4x4_magic_0/RWL_0
rlabel poly 5219 793 5771 823 1 10T_4x4_magic_0/10T_toy_magic_3/WWL
rlabel locali 5698 655 5728 689 1 10T_4x4_magic_0/10T_toy_magic_3/RWL
rlabel locali 5262 655 5292 689 1 10T_4x4_magic_0/10T_toy_magic_3/RWL
rlabel locali 5683 737 5698 766 1 10T_4x4_magic_0/10T_toy_magic_3/WBL
rlabel locali 5293 737 5308 765 1 10T_4x4_magic_0/10T_toy_magic_3/WBLb
rlabel locali 5756 591 5771 633 1 10T_4x4_magic_0/10T_toy_magic_3/RBL0
rlabel locali 5219 591 5234 633 1 10T_4x4_magic_0/10T_toy_magic_3/RBL1
rlabel metal1 5479 779 5511 793 1 10T_4x4_magic_0/10T_toy_magic_3/VDD
rlabel metal1 5479 553 5511 567 7 10T_4x4_magic_0/10T_toy_magic_3/GND
rlabel polycont 5441 660 5471 694 1 10T_4x4_magic_0/10T_toy_magic_3/junc0
rlabel polycont 5519 660 5549 694 1 10T_4x4_magic_0/10T_toy_magic_3/junc1
rlabel ndiff 5292 591 5348 619 1 10T_4x4_magic_0/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 591 5698 619 1 10T_4x4_magic_0/10T_toy_magic_3/RWL0_junc
rlabel poly 4639 793 5191 823 1 10T_4x4_magic_0/10T_toy_magic_2/WWL
rlabel locali 5118 655 5148 689 1 10T_4x4_magic_0/10T_toy_magic_2/RWL
rlabel locali 4682 655 4712 689 1 10T_4x4_magic_0/10T_toy_magic_2/RWL
rlabel locali 5103 737 5118 766 1 10T_4x4_magic_0/10T_toy_magic_2/WBL
rlabel locali 4713 737 4728 765 1 10T_4x4_magic_0/10T_toy_magic_2/WBLb
rlabel locali 5176 591 5191 633 1 10T_4x4_magic_0/10T_toy_magic_2/RBL0
rlabel locali 4639 591 4654 633 1 10T_4x4_magic_0/10T_toy_magic_2/RBL1
rlabel metal1 4899 779 4931 793 1 10T_4x4_magic_0/10T_toy_magic_2/VDD
rlabel metal1 4899 553 4931 567 7 10T_4x4_magic_0/10T_toy_magic_2/GND
rlabel polycont 4861 660 4891 694 1 10T_4x4_magic_0/10T_toy_magic_2/junc0
rlabel polycont 4939 660 4969 694 1 10T_4x4_magic_0/10T_toy_magic_2/junc1
rlabel ndiff 4712 591 4768 619 1 10T_4x4_magic_0/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 591 5118 619 1 10T_4x4_magic_0/10T_toy_magic_2/RWL0_junc
rlabel poly 5219 1063 5771 1093 1 10T_4x4_magic_0/10T_toy_magic_1/WWL
rlabel locali 5698 925 5728 959 1 10T_4x4_magic_0/10T_toy_magic_1/RWL
rlabel locali 5262 925 5292 959 1 10T_4x4_magic_0/10T_toy_magic_1/RWL
rlabel locali 5683 1007 5698 1036 1 10T_4x4_magic_0/10T_toy_magic_1/WBL
rlabel locali 5293 1007 5308 1035 1 10T_4x4_magic_0/10T_toy_magic_1/WBLb
rlabel locali 5756 861 5771 903 1 10T_4x4_magic_0/10T_toy_magic_1/RBL0
rlabel locali 5219 861 5234 903 1 10T_4x4_magic_0/10T_toy_magic_1/RBL1
rlabel metal1 5479 1049 5511 1063 1 10T_4x4_magic_0/10T_toy_magic_1/VDD
rlabel metal1 5479 823 5511 837 7 10T_4x4_magic_0/10T_toy_magic_1/GND
rlabel polycont 5441 930 5471 964 1 10T_4x4_magic_0/10T_toy_magic_1/junc0
rlabel polycont 5519 930 5549 964 1 10T_4x4_magic_0/10T_toy_magic_1/junc1
rlabel ndiff 5292 861 5348 889 1 10T_4x4_magic_0/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 861 5698 889 1 10T_4x4_magic_0/10T_toy_magic_1/RWL0_junc
rlabel poly 4639 1063 5191 1093 1 10T_4x4_magic_0/10T_toy_magic_0/WWL
rlabel locali 5118 925 5148 959 1 10T_4x4_magic_0/10T_toy_magic_0/RWL
rlabel locali 4682 925 4712 959 1 10T_4x4_magic_0/10T_toy_magic_0/RWL
rlabel locali 5103 1007 5118 1036 1 10T_4x4_magic_0/10T_toy_magic_0/WBL
rlabel locali 4713 1007 4728 1035 1 10T_4x4_magic_0/10T_toy_magic_0/WBLb
rlabel locali 5176 861 5191 903 1 10T_4x4_magic_0/10T_toy_magic_0/RBL0
rlabel locali 4639 861 4654 903 1 10T_4x4_magic_0/10T_toy_magic_0/RBL1
rlabel metal1 4899 1049 4931 1063 1 10T_4x4_magic_0/10T_toy_magic_0/VDD
rlabel metal1 4899 823 4931 837 7 10T_4x4_magic_0/10T_toy_magic_0/GND
rlabel polycont 4861 930 4891 964 1 10T_4x4_magic_0/10T_toy_magic_0/junc0
rlabel polycont 4939 930 4969 964 1 10T_4x4_magic_0/10T_toy_magic_0/junc1
rlabel ndiff 4712 861 4768 889 1 10T_4x4_magic_0/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 861 5118 889 1 10T_4x4_magic_0/10T_toy_magic_0/RWL0_junc
rlabel metal1 4591 2130 4621 2144 1 10T_4x4_magic_1/VDD
rlabel metal1 4591 1860 4621 1874 1 10T_4x4_magic_1/VDD
rlabel metal1 4591 1904 4621 1918 1 10T_4x4_magic_1/GND
rlabel metal1 4591 1634 4621 1648 1 10T_4x4_magic_1/GND
rlabel corelocali 4639 1586 4654 1616 1 10T_4x4_magic_1/RBL1_0
rlabel corelocali 5176 1586 5191 1616 1 10T_4x4_magic_1/RBL0_0
rlabel corelocali 5219 1586 5234 1616 1 10T_4x4_magic_1/RBL1_1
rlabel corelocali 5756 1586 5771 1616 1 10T_4x4_magic_1/RBL0_1
rlabel metal1 4591 1736 4621 1770 1 10T_4x4_magic_1/RWL_1
rlabel metal1 4591 2006 4621 2040 1 10T_4x4_magic_1/RWL_0
rlabel locali 5698 1736 5728 1770 1 10T_4x4_magic_1/10T_toy_magic_3/RWL
rlabel locali 5262 1736 5292 1770 1 10T_4x4_magic_1/10T_toy_magic_3/RWL
rlabel locali 5683 1818 5698 1847 1 10T_4x4_magic_1/10T_toy_magic_3/WBL
rlabel locali 5293 1818 5308 1846 1 10T_4x4_magic_1/10T_toy_magic_3/WBLb
rlabel locali 5756 1672 5771 1714 1 10T_4x4_magic_1/10T_toy_magic_3/RBL0
rlabel locali 5219 1672 5234 1714 1 10T_4x4_magic_1/10T_toy_magic_3/RBL1
rlabel metal1 5479 1860 5511 1874 1 10T_4x4_magic_1/10T_toy_magic_3/VDD
rlabel metal1 5479 1634 5511 1648 7 10T_4x4_magic_1/10T_toy_magic_3/GND
rlabel polycont 5441 1741 5471 1775 1 10T_4x4_magic_1/10T_toy_magic_3/junc0
rlabel polycont 5519 1741 5549 1775 1 10T_4x4_magic_1/10T_toy_magic_3/junc1
rlabel ndiff 5292 1672 5348 1700 1 10T_4x4_magic_1/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 1672 5698 1700 1 10T_4x4_magic_1/10T_toy_magic_3/RWL0_junc
rlabel locali 5118 1736 5148 1770 1 10T_4x4_magic_1/10T_toy_magic_2/RWL
rlabel locali 4682 1736 4712 1770 1 10T_4x4_magic_1/10T_toy_magic_2/RWL
rlabel locali 5103 1818 5118 1847 1 10T_4x4_magic_1/10T_toy_magic_2/WBL
rlabel locali 4713 1818 4728 1846 1 10T_4x4_magic_1/10T_toy_magic_2/WBLb
rlabel locali 5176 1672 5191 1714 1 10T_4x4_magic_1/10T_toy_magic_2/RBL0
rlabel locali 4639 1672 4654 1714 1 10T_4x4_magic_1/10T_toy_magic_2/RBL1
rlabel metal1 4899 1860 4931 1874 1 10T_4x4_magic_1/10T_toy_magic_2/VDD
rlabel metal1 4899 1634 4931 1648 7 10T_4x4_magic_1/10T_toy_magic_2/GND
rlabel polycont 4861 1741 4891 1775 1 10T_4x4_magic_1/10T_toy_magic_2/junc0
rlabel polycont 4939 1741 4969 1775 1 10T_4x4_magic_1/10T_toy_magic_2/junc1
rlabel ndiff 4712 1672 4768 1700 1 10T_4x4_magic_1/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 1672 5118 1700 1 10T_4x4_magic_1/10T_toy_magic_2/RWL0_junc
rlabel locali 5698 2006 5728 2040 1 10T_4x4_magic_1/10T_toy_magic_1/RWL
rlabel locali 5262 2006 5292 2040 1 10T_4x4_magic_1/10T_toy_magic_1/RWL
rlabel locali 5683 2088 5698 2117 1 10T_4x4_magic_1/10T_toy_magic_1/WBL
rlabel locali 5293 2088 5308 2116 1 10T_4x4_magic_1/10T_toy_magic_1/WBLb
rlabel locali 5756 1942 5771 1984 1 10T_4x4_magic_1/10T_toy_magic_1/RBL0
rlabel locali 5219 1942 5234 1984 1 10T_4x4_magic_1/10T_toy_magic_1/RBL1
rlabel metal1 5479 2130 5511 2144 1 10T_4x4_magic_1/10T_toy_magic_1/VDD
rlabel metal1 5479 1904 5511 1918 7 10T_4x4_magic_1/10T_toy_magic_1/GND
rlabel polycont 5441 2011 5471 2045 1 10T_4x4_magic_1/10T_toy_magic_1/junc0
rlabel polycont 5519 2011 5549 2045 1 10T_4x4_magic_1/10T_toy_magic_1/junc1
rlabel ndiff 5292 1942 5348 1970 1 10T_4x4_magic_1/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 1942 5698 1970 1 10T_4x4_magic_1/10T_toy_magic_1/RWL0_junc
rlabel locali 5118 2006 5148 2040 1 10T_4x4_magic_1/10T_toy_magic_0/RWL
rlabel locali 4682 2006 4712 2040 1 10T_4x4_magic_1/10T_toy_magic_0/RWL
rlabel locali 5103 2088 5118 2117 1 10T_4x4_magic_1/10T_toy_magic_0/WBL
rlabel locali 4713 2088 4728 2116 1 10T_4x4_magic_1/10T_toy_magic_0/WBLb
rlabel locali 5176 1942 5191 1984 1 10T_4x4_magic_1/10T_toy_magic_0/RBL0
rlabel locali 4639 1942 4654 1984 1 10T_4x4_magic_1/10T_toy_magic_0/RBL1
rlabel metal1 4899 2130 4931 2144 1 10T_4x4_magic_1/10T_toy_magic_0/VDD
rlabel metal1 4899 1904 4931 1918 7 10T_4x4_magic_1/10T_toy_magic_0/GND
rlabel polycont 4861 2011 4891 2045 1 10T_4x4_magic_1/10T_toy_magic_0/junc0
rlabel polycont 4939 2011 4969 2045 1 10T_4x4_magic_1/10T_toy_magic_0/junc1
rlabel ndiff 4712 1942 4768 1970 1 10T_4x4_magic_1/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 1942 5118 1970 1 10T_4x4_magic_1/10T_toy_magic_0/RWL0_junc
rlabel metal1 4591 1590 4621 1604 1 10T_4x4_magic_2/VDD
rlabel metal1 4591 1320 4621 1334 1 10T_4x4_magic_2/VDD
rlabel metal1 4591 1364 4621 1378 1 10T_4x4_magic_2/GND
rlabel metal1 4591 1094 4621 1108 1 10T_4x4_magic_2/GND
rlabel corelocali 4639 1046 4654 1076 1 10T_4x4_magic_2/RBL1_0
rlabel corelocali 5176 1046 5191 1076 1 10T_4x4_magic_2/RBL0_0
rlabel corelocali 5219 1046 5234 1076 1 10T_4x4_magic_2/RBL1_1
rlabel corelocali 5756 1046 5771 1076 1 10T_4x4_magic_2/RBL0_1
rlabel metal1 4591 1196 4621 1230 1 10T_4x4_magic_2/RWL_1
rlabel metal1 4591 1466 4621 1500 1 10T_4x4_magic_2/RWL_0
rlabel locali 5698 1196 5728 1230 1 10T_4x4_magic_2/10T_toy_magic_3/RWL
rlabel locali 5262 1196 5292 1230 1 10T_4x4_magic_2/10T_toy_magic_3/RWL
rlabel locali 5683 1278 5698 1307 1 10T_4x4_magic_2/10T_toy_magic_3/WBL
rlabel locali 5293 1278 5308 1306 1 10T_4x4_magic_2/10T_toy_magic_3/WBLb
rlabel locali 5756 1132 5771 1174 1 10T_4x4_magic_2/10T_toy_magic_3/RBL0
rlabel locali 5219 1132 5234 1174 1 10T_4x4_magic_2/10T_toy_magic_3/RBL1
rlabel metal1 5479 1320 5511 1334 1 10T_4x4_magic_2/10T_toy_magic_3/VDD
rlabel metal1 5479 1094 5511 1108 7 10T_4x4_magic_2/10T_toy_magic_3/GND
rlabel polycont 5441 1201 5471 1235 1 10T_4x4_magic_2/10T_toy_magic_3/junc0
rlabel polycont 5519 1201 5549 1235 1 10T_4x4_magic_2/10T_toy_magic_3/junc1
rlabel ndiff 5292 1132 5348 1160 1 10T_4x4_magic_2/10T_toy_magic_3/RWL1_junc
rlabel ndiff 5642 1132 5698 1160 1 10T_4x4_magic_2/10T_toy_magic_3/RWL0_junc
rlabel locali 5118 1196 5148 1230 1 10T_4x4_magic_2/10T_toy_magic_2/RWL
rlabel locali 4682 1196 4712 1230 1 10T_4x4_magic_2/10T_toy_magic_2/RWL
rlabel locali 5103 1278 5118 1307 1 10T_4x4_magic_2/10T_toy_magic_2/WBL
rlabel locali 4713 1278 4728 1306 1 10T_4x4_magic_2/10T_toy_magic_2/WBLb
rlabel locali 5176 1132 5191 1174 1 10T_4x4_magic_2/10T_toy_magic_2/RBL0
rlabel locali 4639 1132 4654 1174 1 10T_4x4_magic_2/10T_toy_magic_2/RBL1
rlabel metal1 4899 1320 4931 1334 1 10T_4x4_magic_2/10T_toy_magic_2/VDD
rlabel metal1 4899 1094 4931 1108 7 10T_4x4_magic_2/10T_toy_magic_2/GND
rlabel polycont 4861 1201 4891 1235 1 10T_4x4_magic_2/10T_toy_magic_2/junc0
rlabel polycont 4939 1201 4969 1235 1 10T_4x4_magic_2/10T_toy_magic_2/junc1
rlabel ndiff 4712 1132 4768 1160 1 10T_4x4_magic_2/10T_toy_magic_2/RWL1_junc
rlabel ndiff 5062 1132 5118 1160 1 10T_4x4_magic_2/10T_toy_magic_2/RWL0_junc
rlabel locali 5698 1466 5728 1500 1 10T_4x4_magic_2/10T_toy_magic_1/RWL
rlabel locali 5262 1466 5292 1500 1 10T_4x4_magic_2/10T_toy_magic_1/RWL
rlabel locali 5683 1548 5698 1577 1 10T_4x4_magic_2/10T_toy_magic_1/WBL
rlabel locali 5293 1548 5308 1576 1 10T_4x4_magic_2/10T_toy_magic_1/WBLb
rlabel locali 5756 1402 5771 1444 1 10T_4x4_magic_2/10T_toy_magic_1/RBL0
rlabel locali 5219 1402 5234 1444 1 10T_4x4_magic_2/10T_toy_magic_1/RBL1
rlabel metal1 5479 1590 5511 1604 1 10T_4x4_magic_2/10T_toy_magic_1/VDD
rlabel metal1 5479 1364 5511 1378 7 10T_4x4_magic_2/10T_toy_magic_1/GND
rlabel polycont 5441 1471 5471 1505 1 10T_4x4_magic_2/10T_toy_magic_1/junc0
rlabel polycont 5519 1471 5549 1505 1 10T_4x4_magic_2/10T_toy_magic_1/junc1
rlabel ndiff 5292 1402 5348 1430 1 10T_4x4_magic_2/10T_toy_magic_1/RWL1_junc
rlabel ndiff 5642 1402 5698 1430 1 10T_4x4_magic_2/10T_toy_magic_1/RWL0_junc
rlabel locali 5118 1466 5148 1500 1 10T_4x4_magic_2/10T_toy_magic_0/RWL
rlabel locali 4682 1466 4712 1500 1 10T_4x4_magic_2/10T_toy_magic_0/RWL
rlabel locali 5103 1548 5118 1577 1 10T_4x4_magic_2/10T_toy_magic_0/WBL
rlabel locali 4713 1548 4728 1576 1 10T_4x4_magic_2/10T_toy_magic_0/WBLb
rlabel locali 5176 1402 5191 1444 1 10T_4x4_magic_2/10T_toy_magic_0/RBL0
rlabel locali 4639 1402 4654 1444 1 10T_4x4_magic_2/10T_toy_magic_0/RBL1
rlabel metal1 4899 1590 4931 1604 1 10T_4x4_magic_2/10T_toy_magic_0/VDD
rlabel metal1 4899 1364 4931 1378 7 10T_4x4_magic_2/10T_toy_magic_0/GND
rlabel polycont 4861 1471 4891 1505 1 10T_4x4_magic_2/10T_toy_magic_0/junc0
rlabel polycont 4939 1471 4969 1505 1 10T_4x4_magic_2/10T_toy_magic_0/junc1
rlabel ndiff 4712 1402 4768 1430 1 10T_4x4_magic_2/10T_toy_magic_0/RWL1_junc
rlabel ndiff 5062 1402 5118 1430 1 10T_4x4_magic_2/10T_toy_magic_0/RWL0_junc
rlabel poly 5751 523 5781 553 1 10T_4x4_magic_8/WWL_0
rlabel poly 5751 253 5781 283 1 10T_4x4_magic_8/WWL_1
rlabel metal1 5751 509 5781 523 1 10T_4x4_magic_8/VDD
rlabel metal1 5751 239 5781 253 1 10T_4x4_magic_8/VDD
rlabel metal1 5751 283 5781 297 1 10T_4x4_magic_8/GND
rlabel metal1 5751 13 5781 27 1 10T_4x4_magic_8/GND
rlabel corelocali 5799 -35 5814 -5 1 10T_4x4_magic_8/RBL1_0
rlabel corelocali 6336 -35 6351 -5 1 10T_4x4_magic_8/RBL0_0
rlabel corelocali 6379 -35 6394 -5 1 10T_4x4_magic_8/RBL1_1
rlabel corelocali 6916 -35 6931 -5 1 10T_4x4_magic_8/RBL0_1
rlabel metal1 5751 115 5781 149 1 10T_4x4_magic_8/RWL_1
rlabel metal1 5751 385 5781 419 1 10T_4x4_magic_8/RWL_0
rlabel poly 6379 253 6931 283 1 10T_4x4_magic_8/10T_toy_magic_3/WWL
rlabel locali 6858 115 6888 149 1 10T_4x4_magic_8/10T_toy_magic_3/RWL
rlabel locali 6422 115 6452 149 1 10T_4x4_magic_8/10T_toy_magic_3/RWL
rlabel locali 6843 197 6858 226 1 10T_4x4_magic_8/10T_toy_magic_3/WBL
rlabel locali 6453 197 6468 225 1 10T_4x4_magic_8/10T_toy_magic_3/WBLb
rlabel locali 6916 51 6931 93 1 10T_4x4_magic_8/10T_toy_magic_3/RBL0
rlabel locali 6379 51 6394 93 1 10T_4x4_magic_8/10T_toy_magic_3/RBL1
rlabel metal1 6639 239 6671 253 1 10T_4x4_magic_8/10T_toy_magic_3/VDD
rlabel metal1 6639 13 6671 27 7 10T_4x4_magic_8/10T_toy_magic_3/GND
rlabel polycont 6601 120 6631 154 1 10T_4x4_magic_8/10T_toy_magic_3/junc0
rlabel polycont 6679 120 6709 154 1 10T_4x4_magic_8/10T_toy_magic_3/junc1
rlabel ndiff 6452 51 6508 79 1 10T_4x4_magic_8/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 51 6858 79 1 10T_4x4_magic_8/10T_toy_magic_3/RWL0_junc
rlabel poly 5799 253 6351 283 1 10T_4x4_magic_8/10T_toy_magic_2/WWL
rlabel locali 6278 115 6308 149 1 10T_4x4_magic_8/10T_toy_magic_2/RWL
rlabel locali 5842 115 5872 149 1 10T_4x4_magic_8/10T_toy_magic_2/RWL
rlabel locali 6263 197 6278 226 1 10T_4x4_magic_8/10T_toy_magic_2/WBL
rlabel locali 5873 197 5888 225 1 10T_4x4_magic_8/10T_toy_magic_2/WBLb
rlabel locali 6336 51 6351 93 1 10T_4x4_magic_8/10T_toy_magic_2/RBL0
rlabel locali 5799 51 5814 93 1 10T_4x4_magic_8/10T_toy_magic_2/RBL1
rlabel metal1 6059 239 6091 253 1 10T_4x4_magic_8/10T_toy_magic_2/VDD
rlabel metal1 6059 13 6091 27 7 10T_4x4_magic_8/10T_toy_magic_2/GND
rlabel polycont 6021 120 6051 154 1 10T_4x4_magic_8/10T_toy_magic_2/junc0
rlabel polycont 6099 120 6129 154 1 10T_4x4_magic_8/10T_toy_magic_2/junc1
rlabel ndiff 5872 51 5928 79 1 10T_4x4_magic_8/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 51 6278 79 1 10T_4x4_magic_8/10T_toy_magic_2/RWL0_junc
rlabel poly 6379 523 6931 553 1 10T_4x4_magic_8/10T_toy_magic_1/WWL
rlabel locali 6858 385 6888 419 1 10T_4x4_magic_8/10T_toy_magic_1/RWL
rlabel locali 6422 385 6452 419 1 10T_4x4_magic_8/10T_toy_magic_1/RWL
rlabel locali 6843 467 6858 496 1 10T_4x4_magic_8/10T_toy_magic_1/WBL
rlabel locali 6453 467 6468 495 1 10T_4x4_magic_8/10T_toy_magic_1/WBLb
rlabel locali 6916 321 6931 363 1 10T_4x4_magic_8/10T_toy_magic_1/RBL0
rlabel locali 6379 321 6394 363 1 10T_4x4_magic_8/10T_toy_magic_1/RBL1
rlabel metal1 6639 509 6671 523 1 10T_4x4_magic_8/10T_toy_magic_1/VDD
rlabel metal1 6639 283 6671 297 7 10T_4x4_magic_8/10T_toy_magic_1/GND
rlabel polycont 6601 390 6631 424 1 10T_4x4_magic_8/10T_toy_magic_1/junc0
rlabel polycont 6679 390 6709 424 1 10T_4x4_magic_8/10T_toy_magic_1/junc1
rlabel ndiff 6452 321 6508 349 1 10T_4x4_magic_8/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 321 6858 349 1 10T_4x4_magic_8/10T_toy_magic_1/RWL0_junc
rlabel poly 5799 523 6351 553 1 10T_4x4_magic_8/10T_toy_magic_0/WWL
rlabel locali 6278 385 6308 419 1 10T_4x4_magic_8/10T_toy_magic_0/RWL
rlabel locali 5842 385 5872 419 1 10T_4x4_magic_8/10T_toy_magic_0/RWL
rlabel locali 6263 467 6278 496 1 10T_4x4_magic_8/10T_toy_magic_0/WBL
rlabel locali 5873 467 5888 495 1 10T_4x4_magic_8/10T_toy_magic_0/WBLb
rlabel locali 6336 321 6351 363 1 10T_4x4_magic_8/10T_toy_magic_0/RBL0
rlabel locali 5799 321 5814 363 1 10T_4x4_magic_8/10T_toy_magic_0/RBL1
rlabel metal1 6059 509 6091 523 1 10T_4x4_magic_8/10T_toy_magic_0/VDD
rlabel metal1 6059 283 6091 297 7 10T_4x4_magic_8/10T_toy_magic_0/GND
rlabel polycont 6021 390 6051 424 1 10T_4x4_magic_8/10T_toy_magic_0/junc0
rlabel polycont 6099 390 6129 424 1 10T_4x4_magic_8/10T_toy_magic_0/junc1
rlabel ndiff 5872 321 5928 349 1 10T_4x4_magic_8/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 321 6278 349 1 10T_4x4_magic_8/10T_toy_magic_0/RWL0_junc
rlabel poly 5751 -17 5781 13 1 10T_4x4_magic_9/WWL_0
rlabel poly 5751 -287 5781 -257 1 10T_4x4_magic_9/WWL_1
rlabel metal1 5751 -31 5781 -17 1 10T_4x4_magic_9/VDD
rlabel metal1 5751 -301 5781 -287 1 10T_4x4_magic_9/VDD
rlabel metal1 5751 -257 5781 -243 1 10T_4x4_magic_9/GND
rlabel metal1 5751 -527 5781 -513 1 10T_4x4_magic_9/GND
rlabel corelocali 5799 -575 5814 -545 1 10T_4x4_magic_9/RBL1_0
rlabel corelocali 6336 -575 6351 -545 1 10T_4x4_magic_9/RBL0_0
rlabel corelocali 6379 -575 6394 -545 1 10T_4x4_magic_9/RBL1_1
rlabel corelocali 6916 -575 6931 -545 1 10T_4x4_magic_9/RBL0_1
rlabel metal1 5751 -425 5781 -391 1 10T_4x4_magic_9/RWL_1
rlabel metal1 5751 -155 5781 -121 1 10T_4x4_magic_9/RWL_0
rlabel poly 6379 -287 6931 -257 1 10T_4x4_magic_9/10T_toy_magic_3/WWL
rlabel locali 6858 -425 6888 -391 1 10T_4x4_magic_9/10T_toy_magic_3/RWL
rlabel locali 6422 -425 6452 -391 1 10T_4x4_magic_9/10T_toy_magic_3/RWL
rlabel locali 6843 -343 6858 -314 1 10T_4x4_magic_9/10T_toy_magic_3/WBL
rlabel locali 6453 -343 6468 -315 1 10T_4x4_magic_9/10T_toy_magic_3/WBLb
rlabel locali 6916 -489 6931 -447 1 10T_4x4_magic_9/10T_toy_magic_3/RBL0
rlabel locali 6379 -489 6394 -447 1 10T_4x4_magic_9/10T_toy_magic_3/RBL1
rlabel metal1 6639 -301 6671 -287 1 10T_4x4_magic_9/10T_toy_magic_3/VDD
rlabel metal1 6639 -527 6671 -513 7 10T_4x4_magic_9/10T_toy_magic_3/GND
rlabel polycont 6601 -420 6631 -386 1 10T_4x4_magic_9/10T_toy_magic_3/junc0
rlabel polycont 6679 -420 6709 -386 1 10T_4x4_magic_9/10T_toy_magic_3/junc1
rlabel ndiff 6452 -489 6508 -461 1 10T_4x4_magic_9/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 -489 6858 -461 1 10T_4x4_magic_9/10T_toy_magic_3/RWL0_junc
rlabel poly 5799 -287 6351 -257 1 10T_4x4_magic_9/10T_toy_magic_2/WWL
rlabel locali 6278 -425 6308 -391 1 10T_4x4_magic_9/10T_toy_magic_2/RWL
rlabel locali 5842 -425 5872 -391 1 10T_4x4_magic_9/10T_toy_magic_2/RWL
rlabel locali 6263 -343 6278 -314 1 10T_4x4_magic_9/10T_toy_magic_2/WBL
rlabel locali 5873 -343 5888 -315 1 10T_4x4_magic_9/10T_toy_magic_2/WBLb
rlabel locali 6336 -489 6351 -447 1 10T_4x4_magic_9/10T_toy_magic_2/RBL0
rlabel locali 5799 -489 5814 -447 1 10T_4x4_magic_9/10T_toy_magic_2/RBL1
rlabel metal1 6059 -301 6091 -287 1 10T_4x4_magic_9/10T_toy_magic_2/VDD
rlabel metal1 6059 -527 6091 -513 7 10T_4x4_magic_9/10T_toy_magic_2/GND
rlabel polycont 6021 -420 6051 -386 1 10T_4x4_magic_9/10T_toy_magic_2/junc0
rlabel polycont 6099 -420 6129 -386 1 10T_4x4_magic_9/10T_toy_magic_2/junc1
rlabel ndiff 5872 -489 5928 -461 1 10T_4x4_magic_9/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 -489 6278 -461 1 10T_4x4_magic_9/10T_toy_magic_2/RWL0_junc
rlabel poly 6379 -17 6931 13 1 10T_4x4_magic_9/10T_toy_magic_1/WWL
rlabel locali 6858 -155 6888 -121 1 10T_4x4_magic_9/10T_toy_magic_1/RWL
rlabel locali 6422 -155 6452 -121 1 10T_4x4_magic_9/10T_toy_magic_1/RWL
rlabel locali 6843 -73 6858 -44 1 10T_4x4_magic_9/10T_toy_magic_1/WBL
rlabel locali 6453 -73 6468 -45 1 10T_4x4_magic_9/10T_toy_magic_1/WBLb
rlabel locali 6916 -219 6931 -177 1 10T_4x4_magic_9/10T_toy_magic_1/RBL0
rlabel locali 6379 -219 6394 -177 1 10T_4x4_magic_9/10T_toy_magic_1/RBL1
rlabel metal1 6639 -31 6671 -17 1 10T_4x4_magic_9/10T_toy_magic_1/VDD
rlabel metal1 6639 -257 6671 -243 7 10T_4x4_magic_9/10T_toy_magic_1/GND
rlabel polycont 6601 -150 6631 -116 1 10T_4x4_magic_9/10T_toy_magic_1/junc0
rlabel polycont 6679 -150 6709 -116 1 10T_4x4_magic_9/10T_toy_magic_1/junc1
rlabel ndiff 6452 -219 6508 -191 1 10T_4x4_magic_9/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 -219 6858 -191 1 10T_4x4_magic_9/10T_toy_magic_1/RWL0_junc
rlabel poly 5799 -17 6351 13 1 10T_4x4_magic_9/10T_toy_magic_0/WWL
rlabel locali 6278 -155 6308 -121 1 10T_4x4_magic_9/10T_toy_magic_0/RWL
rlabel locali 5842 -155 5872 -121 1 10T_4x4_magic_9/10T_toy_magic_0/RWL
rlabel locali 6263 -73 6278 -44 1 10T_4x4_magic_9/10T_toy_magic_0/WBL
rlabel locali 5873 -73 5888 -45 1 10T_4x4_magic_9/10T_toy_magic_0/WBLb
rlabel locali 6336 -219 6351 -177 1 10T_4x4_magic_9/10T_toy_magic_0/RBL0
rlabel locali 5799 -219 5814 -177 1 10T_4x4_magic_9/10T_toy_magic_0/RBL1
rlabel metal1 6059 -31 6091 -17 1 10T_4x4_magic_9/10T_toy_magic_0/VDD
rlabel metal1 6059 -257 6091 -243 7 10T_4x4_magic_9/10T_toy_magic_0/GND
rlabel polycont 6021 -150 6051 -116 1 10T_4x4_magic_9/10T_toy_magic_0/junc0
rlabel polycont 6099 -150 6129 -116 1 10T_4x4_magic_9/10T_toy_magic_0/junc1
rlabel ndiff 5872 -219 5928 -191 1 10T_4x4_magic_9/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 -219 6278 -191 1 10T_4x4_magic_9/10T_toy_magic_0/RWL0_junc
rlabel poly 5751 -557 5781 -527 1 10T_4x4_magic_10/WWL_0
rlabel poly 5751 -827 5781 -797 1 10T_4x4_magic_10/WWL_1
rlabel metal1 5751 -571 5781 -557 1 10T_4x4_magic_10/VDD
rlabel metal1 5751 -841 5781 -827 1 10T_4x4_magic_10/VDD
rlabel metal1 5751 -797 5781 -783 1 10T_4x4_magic_10/GND
rlabel metal1 5751 -1067 5781 -1053 1 10T_4x4_magic_10/GND
rlabel corelocali 5799 -1115 5814 -1085 1 10T_4x4_magic_10/RBL1_0
rlabel corelocali 6336 -1115 6351 -1085 1 10T_4x4_magic_10/RBL0_0
rlabel corelocali 6379 -1115 6394 -1085 1 10T_4x4_magic_10/RBL1_1
rlabel corelocali 6916 -1115 6931 -1085 1 10T_4x4_magic_10/RBL0_1
rlabel metal1 5751 -965 5781 -931 1 10T_4x4_magic_10/RWL_1
rlabel metal1 5751 -695 5781 -661 1 10T_4x4_magic_10/RWL_0
rlabel poly 6379 -827 6931 -797 1 10T_4x4_magic_10/10T_toy_magic_3/WWL
rlabel locali 6858 -965 6888 -931 1 10T_4x4_magic_10/10T_toy_magic_3/RWL
rlabel locali 6422 -965 6452 -931 1 10T_4x4_magic_10/10T_toy_magic_3/RWL
rlabel locali 6843 -883 6858 -854 1 10T_4x4_magic_10/10T_toy_magic_3/WBL
rlabel locali 6453 -883 6468 -855 1 10T_4x4_magic_10/10T_toy_magic_3/WBLb
rlabel locali 6916 -1029 6931 -987 1 10T_4x4_magic_10/10T_toy_magic_3/RBL0
rlabel locali 6379 -1029 6394 -987 1 10T_4x4_magic_10/10T_toy_magic_3/RBL1
rlabel metal1 6639 -841 6671 -827 1 10T_4x4_magic_10/10T_toy_magic_3/VDD
rlabel metal1 6639 -1067 6671 -1053 7 10T_4x4_magic_10/10T_toy_magic_3/GND
rlabel polycont 6601 -960 6631 -926 1 10T_4x4_magic_10/10T_toy_magic_3/junc0
rlabel polycont 6679 -960 6709 -926 1 10T_4x4_magic_10/10T_toy_magic_3/junc1
rlabel ndiff 6452 -1029 6508 -1001 1 10T_4x4_magic_10/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 -1029 6858 -1001 1 10T_4x4_magic_10/10T_toy_magic_3/RWL0_junc
rlabel poly 5799 -827 6351 -797 1 10T_4x4_magic_10/10T_toy_magic_2/WWL
rlabel locali 6278 -965 6308 -931 1 10T_4x4_magic_10/10T_toy_magic_2/RWL
rlabel locali 5842 -965 5872 -931 1 10T_4x4_magic_10/10T_toy_magic_2/RWL
rlabel locali 6263 -883 6278 -854 1 10T_4x4_magic_10/10T_toy_magic_2/WBL
rlabel locali 5873 -883 5888 -855 1 10T_4x4_magic_10/10T_toy_magic_2/WBLb
rlabel locali 6336 -1029 6351 -987 1 10T_4x4_magic_10/10T_toy_magic_2/RBL0
rlabel locali 5799 -1029 5814 -987 1 10T_4x4_magic_10/10T_toy_magic_2/RBL1
rlabel metal1 6059 -841 6091 -827 1 10T_4x4_magic_10/10T_toy_magic_2/VDD
rlabel metal1 6059 -1067 6091 -1053 7 10T_4x4_magic_10/10T_toy_magic_2/GND
rlabel polycont 6021 -960 6051 -926 1 10T_4x4_magic_10/10T_toy_magic_2/junc0
rlabel polycont 6099 -960 6129 -926 1 10T_4x4_magic_10/10T_toy_magic_2/junc1
rlabel ndiff 5872 -1029 5928 -1001 1 10T_4x4_magic_10/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 -1029 6278 -1001 1 10T_4x4_magic_10/10T_toy_magic_2/RWL0_junc
rlabel poly 6379 -557 6931 -527 1 10T_4x4_magic_10/10T_toy_magic_1/WWL
rlabel locali 6858 -695 6888 -661 1 10T_4x4_magic_10/10T_toy_magic_1/RWL
rlabel locali 6422 -695 6452 -661 1 10T_4x4_magic_10/10T_toy_magic_1/RWL
rlabel locali 6843 -613 6858 -584 1 10T_4x4_magic_10/10T_toy_magic_1/WBL
rlabel locali 6453 -613 6468 -585 1 10T_4x4_magic_10/10T_toy_magic_1/WBLb
rlabel locali 6916 -759 6931 -717 1 10T_4x4_magic_10/10T_toy_magic_1/RBL0
rlabel locali 6379 -759 6394 -717 1 10T_4x4_magic_10/10T_toy_magic_1/RBL1
rlabel metal1 6639 -571 6671 -557 1 10T_4x4_magic_10/10T_toy_magic_1/VDD
rlabel metal1 6639 -797 6671 -783 7 10T_4x4_magic_10/10T_toy_magic_1/GND
rlabel polycont 6601 -690 6631 -656 1 10T_4x4_magic_10/10T_toy_magic_1/junc0
rlabel polycont 6679 -690 6709 -656 1 10T_4x4_magic_10/10T_toy_magic_1/junc1
rlabel ndiff 6452 -759 6508 -731 1 10T_4x4_magic_10/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 -759 6858 -731 1 10T_4x4_magic_10/10T_toy_magic_1/RWL0_junc
rlabel poly 5799 -557 6351 -527 1 10T_4x4_magic_10/10T_toy_magic_0/WWL
rlabel locali 6278 -695 6308 -661 1 10T_4x4_magic_10/10T_toy_magic_0/RWL
rlabel locali 5842 -695 5872 -661 1 10T_4x4_magic_10/10T_toy_magic_0/RWL
rlabel locali 6263 -613 6278 -584 1 10T_4x4_magic_10/10T_toy_magic_0/WBL
rlabel locali 5873 -613 5888 -585 1 10T_4x4_magic_10/10T_toy_magic_0/WBLb
rlabel locali 6336 -759 6351 -717 1 10T_4x4_magic_10/10T_toy_magic_0/RBL0
rlabel locali 5799 -759 5814 -717 1 10T_4x4_magic_10/10T_toy_magic_0/RBL1
rlabel metal1 6059 -571 6091 -557 1 10T_4x4_magic_10/10T_toy_magic_0/VDD
rlabel metal1 6059 -797 6091 -783 7 10T_4x4_magic_10/10T_toy_magic_0/GND
rlabel polycont 6021 -690 6051 -656 1 10T_4x4_magic_10/10T_toy_magic_0/junc0
rlabel polycont 6099 -690 6129 -656 1 10T_4x4_magic_10/10T_toy_magic_0/junc1
rlabel ndiff 5872 -759 5928 -731 1 10T_4x4_magic_10/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 -759 6278 -731 1 10T_4x4_magic_10/10T_toy_magic_0/RWL0_junc
rlabel poly 5751 -1097 5781 -1067 1 10T_4x4_magic_11/WWL_0
rlabel poly 5751 -1367 5781 -1337 1 10T_4x4_magic_11/WWL_1
rlabel metal1 5751 -1111 5781 -1097 1 10T_4x4_magic_11/VDD
rlabel metal1 5751 -1381 5781 -1367 1 10T_4x4_magic_11/VDD
rlabel metal1 5751 -1337 5781 -1323 1 10T_4x4_magic_11/GND
rlabel metal1 5751 -1607 5781 -1593 1 10T_4x4_magic_11/GND
rlabel corelocali 5799 -1655 5814 -1625 1 10T_4x4_magic_11/RBL1_0
rlabel corelocali 6336 -1655 6351 -1625 1 10T_4x4_magic_11/RBL0_0
rlabel corelocali 6379 -1655 6394 -1625 1 10T_4x4_magic_11/RBL1_1
rlabel corelocali 6916 -1655 6931 -1625 1 10T_4x4_magic_11/RBL0_1
rlabel metal1 5751 -1505 5781 -1471 1 10T_4x4_magic_11/RWL_1
rlabel metal1 5751 -1235 5781 -1201 1 10T_4x4_magic_11/RWL_0
rlabel poly 6379 -1367 6931 -1337 1 10T_4x4_magic_11/10T_toy_magic_3/WWL
rlabel locali 6858 -1505 6888 -1471 1 10T_4x4_magic_11/10T_toy_magic_3/RWL
rlabel locali 6422 -1505 6452 -1471 1 10T_4x4_magic_11/10T_toy_magic_3/RWL
rlabel locali 6843 -1423 6858 -1394 1 10T_4x4_magic_11/10T_toy_magic_3/WBL
rlabel locali 6453 -1423 6468 -1395 1 10T_4x4_magic_11/10T_toy_magic_3/WBLb
rlabel locali 6916 -1569 6931 -1527 1 10T_4x4_magic_11/10T_toy_magic_3/RBL0
rlabel locali 6379 -1569 6394 -1527 1 10T_4x4_magic_11/10T_toy_magic_3/RBL1
rlabel metal1 6639 -1381 6671 -1367 1 10T_4x4_magic_11/10T_toy_magic_3/VDD
rlabel metal1 6639 -1607 6671 -1593 7 10T_4x4_magic_11/10T_toy_magic_3/GND
rlabel polycont 6601 -1500 6631 -1466 1 10T_4x4_magic_11/10T_toy_magic_3/junc0
rlabel polycont 6679 -1500 6709 -1466 1 10T_4x4_magic_11/10T_toy_magic_3/junc1
rlabel ndiff 6452 -1569 6508 -1541 1 10T_4x4_magic_11/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 -1569 6858 -1541 1 10T_4x4_magic_11/10T_toy_magic_3/RWL0_junc
rlabel poly 5799 -1367 6351 -1337 1 10T_4x4_magic_11/10T_toy_magic_2/WWL
rlabel locali 6278 -1505 6308 -1471 1 10T_4x4_magic_11/10T_toy_magic_2/RWL
rlabel locali 5842 -1505 5872 -1471 1 10T_4x4_magic_11/10T_toy_magic_2/RWL
rlabel locali 6263 -1423 6278 -1394 1 10T_4x4_magic_11/10T_toy_magic_2/WBL
rlabel locali 5873 -1423 5888 -1395 1 10T_4x4_magic_11/10T_toy_magic_2/WBLb
rlabel locali 6336 -1569 6351 -1527 1 10T_4x4_magic_11/10T_toy_magic_2/RBL0
rlabel locali 5799 -1569 5814 -1527 1 10T_4x4_magic_11/10T_toy_magic_2/RBL1
rlabel metal1 6059 -1381 6091 -1367 1 10T_4x4_magic_11/10T_toy_magic_2/VDD
rlabel metal1 6059 -1607 6091 -1593 7 10T_4x4_magic_11/10T_toy_magic_2/GND
rlabel polycont 6021 -1500 6051 -1466 1 10T_4x4_magic_11/10T_toy_magic_2/junc0
rlabel polycont 6099 -1500 6129 -1466 1 10T_4x4_magic_11/10T_toy_magic_2/junc1
rlabel ndiff 5872 -1569 5928 -1541 1 10T_4x4_magic_11/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 -1569 6278 -1541 1 10T_4x4_magic_11/10T_toy_magic_2/RWL0_junc
rlabel poly 6379 -1097 6931 -1067 1 10T_4x4_magic_11/10T_toy_magic_1/WWL
rlabel locali 6858 -1235 6888 -1201 1 10T_4x4_magic_11/10T_toy_magic_1/RWL
rlabel locali 6422 -1235 6452 -1201 1 10T_4x4_magic_11/10T_toy_magic_1/RWL
rlabel locali 6843 -1153 6858 -1124 1 10T_4x4_magic_11/10T_toy_magic_1/WBL
rlabel locali 6453 -1153 6468 -1125 1 10T_4x4_magic_11/10T_toy_magic_1/WBLb
rlabel locali 6916 -1299 6931 -1257 1 10T_4x4_magic_11/10T_toy_magic_1/RBL0
rlabel locali 6379 -1299 6394 -1257 1 10T_4x4_magic_11/10T_toy_magic_1/RBL1
rlabel metal1 6639 -1111 6671 -1097 1 10T_4x4_magic_11/10T_toy_magic_1/VDD
rlabel metal1 6639 -1337 6671 -1323 7 10T_4x4_magic_11/10T_toy_magic_1/GND
rlabel polycont 6601 -1230 6631 -1196 1 10T_4x4_magic_11/10T_toy_magic_1/junc0
rlabel polycont 6679 -1230 6709 -1196 1 10T_4x4_magic_11/10T_toy_magic_1/junc1
rlabel ndiff 6452 -1299 6508 -1271 1 10T_4x4_magic_11/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 -1299 6858 -1271 1 10T_4x4_magic_11/10T_toy_magic_1/RWL0_junc
rlabel poly 5799 -1097 6351 -1067 1 10T_4x4_magic_11/10T_toy_magic_0/WWL
rlabel locali 6278 -1235 6308 -1201 1 10T_4x4_magic_11/10T_toy_magic_0/RWL
rlabel locali 5842 -1235 5872 -1201 1 10T_4x4_magic_11/10T_toy_magic_0/RWL
rlabel locali 6263 -1153 6278 -1124 1 10T_4x4_magic_11/10T_toy_magic_0/WBL
rlabel locali 5873 -1153 5888 -1125 1 10T_4x4_magic_11/10T_toy_magic_0/WBLb
rlabel locali 6336 -1299 6351 -1257 1 10T_4x4_magic_11/10T_toy_magic_0/RBL0
rlabel locali 5799 -1299 5814 -1257 1 10T_4x4_magic_11/10T_toy_magic_0/RBL1
rlabel metal1 6059 -1111 6091 -1097 1 10T_4x4_magic_11/10T_toy_magic_0/VDD
rlabel metal1 6059 -1337 6091 -1323 7 10T_4x4_magic_11/10T_toy_magic_0/GND
rlabel polycont 6021 -1230 6051 -1196 1 10T_4x4_magic_11/10T_toy_magic_0/junc0
rlabel polycont 6099 -1230 6129 -1196 1 10T_4x4_magic_11/10T_toy_magic_0/junc1
rlabel ndiff 5872 -1299 5928 -1271 1 10T_4x4_magic_11/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 -1299 6278 -1271 1 10T_4x4_magic_11/10T_toy_magic_0/RWL0_junc
rlabel poly 5751 -1637 5781 -1607 1 10T_4x4_magic_12/WWL_0
rlabel poly 5751 -1907 5781 -1877 1 10T_4x4_magic_12/WWL_1
rlabel metal1 5751 -1651 5781 -1637 1 10T_4x4_magic_12/VDD
rlabel metal1 5751 -1921 5781 -1907 1 10T_4x4_magic_12/VDD
rlabel metal1 5751 -1877 5781 -1863 1 10T_4x4_magic_12/GND
rlabel metal1 5751 -2147 5781 -2133 1 10T_4x4_magic_12/GND
rlabel metal1 5751 -2045 5781 -2011 1 10T_4x4_magic_12/RWL_1
rlabel metal1 5751 -1775 5781 -1741 1 10T_4x4_magic_12/RWL_0
rlabel poly 6379 -1907 6931 -1877 1 10T_4x4_magic_12/10T_toy_magic_3/WWL
rlabel locali 6858 -2045 6888 -2011 1 10T_4x4_magic_12/10T_toy_magic_3/RWL
rlabel locali 6422 -2045 6452 -2011 1 10T_4x4_magic_12/10T_toy_magic_3/RWL
rlabel locali 6843 -1963 6858 -1934 1 10T_4x4_magic_12/10T_toy_magic_3/WBL
rlabel locali 6453 -1963 6468 -1935 1 10T_4x4_magic_12/10T_toy_magic_3/WBLb
rlabel locali 6916 -2109 6931 -2067 1 10T_4x4_magic_12/10T_toy_magic_3/RBL0
rlabel locali 6379 -2109 6394 -2067 1 10T_4x4_magic_12/10T_toy_magic_3/RBL1
rlabel metal1 6639 -1921 6671 -1907 1 10T_4x4_magic_12/10T_toy_magic_3/VDD
rlabel metal1 6639 -2147 6671 -2133 7 10T_4x4_magic_12/10T_toy_magic_3/GND
rlabel polycont 6601 -2040 6631 -2006 1 10T_4x4_magic_12/10T_toy_magic_3/junc0
rlabel polycont 6679 -2040 6709 -2006 1 10T_4x4_magic_12/10T_toy_magic_3/junc1
rlabel ndiff 6452 -2109 6508 -2081 1 10T_4x4_magic_12/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 -2109 6858 -2081 1 10T_4x4_magic_12/10T_toy_magic_3/RWL0_junc
rlabel poly 5799 -1907 6351 -1877 1 10T_4x4_magic_12/10T_toy_magic_2/WWL
rlabel locali 6278 -2045 6308 -2011 1 10T_4x4_magic_12/10T_toy_magic_2/RWL
rlabel locali 5842 -2045 5872 -2011 1 10T_4x4_magic_12/10T_toy_magic_2/RWL
rlabel locali 6263 -1963 6278 -1934 1 10T_4x4_magic_12/10T_toy_magic_2/WBL
rlabel locali 5873 -1963 5888 -1935 1 10T_4x4_magic_12/10T_toy_magic_2/WBLb
rlabel locali 6336 -2109 6351 -2067 1 10T_4x4_magic_12/10T_toy_magic_2/RBL0
rlabel locali 5799 -2109 5814 -2067 1 10T_4x4_magic_12/10T_toy_magic_2/RBL1
rlabel metal1 6059 -1921 6091 -1907 1 10T_4x4_magic_12/10T_toy_magic_2/VDD
rlabel metal1 6059 -2147 6091 -2133 7 10T_4x4_magic_12/10T_toy_magic_2/GND
rlabel polycont 6021 -2040 6051 -2006 1 10T_4x4_magic_12/10T_toy_magic_2/junc0
rlabel polycont 6099 -2040 6129 -2006 1 10T_4x4_magic_12/10T_toy_magic_2/junc1
rlabel ndiff 5872 -2109 5928 -2081 1 10T_4x4_magic_12/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 -2109 6278 -2081 1 10T_4x4_magic_12/10T_toy_magic_2/RWL0_junc
rlabel poly 6379 -1637 6931 -1607 1 10T_4x4_magic_12/10T_toy_magic_1/WWL
rlabel locali 6858 -1775 6888 -1741 1 10T_4x4_magic_12/10T_toy_magic_1/RWL
rlabel locali 6422 -1775 6452 -1741 1 10T_4x4_magic_12/10T_toy_magic_1/RWL
rlabel locali 6843 -1693 6858 -1664 1 10T_4x4_magic_12/10T_toy_magic_1/WBL
rlabel locali 6453 -1693 6468 -1665 1 10T_4x4_magic_12/10T_toy_magic_1/WBLb
rlabel locali 6916 -1839 6931 -1797 1 10T_4x4_magic_12/10T_toy_magic_1/RBL0
rlabel locali 6379 -1839 6394 -1797 1 10T_4x4_magic_12/10T_toy_magic_1/RBL1
rlabel metal1 6639 -1651 6671 -1637 1 10T_4x4_magic_12/10T_toy_magic_1/VDD
rlabel metal1 6639 -1877 6671 -1863 7 10T_4x4_magic_12/10T_toy_magic_1/GND
rlabel polycont 6601 -1770 6631 -1736 1 10T_4x4_magic_12/10T_toy_magic_1/junc0
rlabel polycont 6679 -1770 6709 -1736 1 10T_4x4_magic_12/10T_toy_magic_1/junc1
rlabel ndiff 6452 -1839 6508 -1811 1 10T_4x4_magic_12/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 -1839 6858 -1811 1 10T_4x4_magic_12/10T_toy_magic_1/RWL0_junc
rlabel poly 5799 -1637 6351 -1607 1 10T_4x4_magic_12/10T_toy_magic_0/WWL
rlabel locali 6278 -1775 6308 -1741 1 10T_4x4_magic_12/10T_toy_magic_0/RWL
rlabel locali 5842 -1775 5872 -1741 1 10T_4x4_magic_12/10T_toy_magic_0/RWL
rlabel locali 6263 -1693 6278 -1664 1 10T_4x4_magic_12/10T_toy_magic_0/WBL
rlabel locali 5873 -1693 5888 -1665 1 10T_4x4_magic_12/10T_toy_magic_0/WBLb
rlabel locali 6336 -1839 6351 -1797 1 10T_4x4_magic_12/10T_toy_magic_0/RBL0
rlabel locali 5799 -1839 5814 -1797 1 10T_4x4_magic_12/10T_toy_magic_0/RBL1
rlabel metal1 6059 -1651 6091 -1637 1 10T_4x4_magic_12/10T_toy_magic_0/VDD
rlabel metal1 6059 -1877 6091 -1863 7 10T_4x4_magic_12/10T_toy_magic_0/GND
rlabel polycont 6021 -1770 6051 -1736 1 10T_4x4_magic_12/10T_toy_magic_0/junc0
rlabel polycont 6099 -1770 6129 -1736 1 10T_4x4_magic_12/10T_toy_magic_0/junc1
rlabel ndiff 5872 -1839 5928 -1811 1 10T_4x4_magic_12/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 -1839 6278 -1811 1 10T_4x4_magic_12/10T_toy_magic_0/RWL0_junc
rlabel poly 5751 1063 5781 1093 1 10T_4x4_magic_13/WWL_0
rlabel poly 5751 793 5781 823 1 10T_4x4_magic_13/WWL_1
rlabel metal1 5751 1049 5781 1063 1 10T_4x4_magic_13/VDD
rlabel metal1 5751 779 5781 793 1 10T_4x4_magic_13/VDD
rlabel metal1 5751 823 5781 837 1 10T_4x4_magic_13/GND
rlabel metal1 5751 553 5781 567 1 10T_4x4_magic_13/GND
rlabel corelocali 5799 505 5814 535 1 10T_4x4_magic_13/RBL1_0
rlabel corelocali 6336 505 6351 535 1 10T_4x4_magic_13/RBL0_0
rlabel corelocali 6379 505 6394 535 1 10T_4x4_magic_13/RBL1_1
rlabel corelocali 6916 505 6931 535 1 10T_4x4_magic_13/RBL0_1
rlabel metal1 5751 655 5781 689 1 10T_4x4_magic_13/RWL_1
rlabel metal1 5751 925 5781 959 1 10T_4x4_magic_13/RWL_0
rlabel poly 6379 793 6931 823 1 10T_4x4_magic_13/10T_toy_magic_3/WWL
rlabel locali 6858 655 6888 689 1 10T_4x4_magic_13/10T_toy_magic_3/RWL
rlabel locali 6422 655 6452 689 1 10T_4x4_magic_13/10T_toy_magic_3/RWL
rlabel locali 6843 737 6858 766 1 10T_4x4_magic_13/10T_toy_magic_3/WBL
rlabel locali 6453 737 6468 765 1 10T_4x4_magic_13/10T_toy_magic_3/WBLb
rlabel locali 6916 591 6931 633 1 10T_4x4_magic_13/10T_toy_magic_3/RBL0
rlabel locali 6379 591 6394 633 1 10T_4x4_magic_13/10T_toy_magic_3/RBL1
rlabel metal1 6639 779 6671 793 1 10T_4x4_magic_13/10T_toy_magic_3/VDD
rlabel metal1 6639 553 6671 567 7 10T_4x4_magic_13/10T_toy_magic_3/GND
rlabel polycont 6601 660 6631 694 1 10T_4x4_magic_13/10T_toy_magic_3/junc0
rlabel polycont 6679 660 6709 694 1 10T_4x4_magic_13/10T_toy_magic_3/junc1
rlabel ndiff 6452 591 6508 619 1 10T_4x4_magic_13/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 591 6858 619 1 10T_4x4_magic_13/10T_toy_magic_3/RWL0_junc
rlabel poly 5799 793 6351 823 1 10T_4x4_magic_13/10T_toy_magic_2/WWL
rlabel locali 6278 655 6308 689 1 10T_4x4_magic_13/10T_toy_magic_2/RWL
rlabel locali 5842 655 5872 689 1 10T_4x4_magic_13/10T_toy_magic_2/RWL
rlabel locali 6263 737 6278 766 1 10T_4x4_magic_13/10T_toy_magic_2/WBL
rlabel locali 5873 737 5888 765 1 10T_4x4_magic_13/10T_toy_magic_2/WBLb
rlabel locali 6336 591 6351 633 1 10T_4x4_magic_13/10T_toy_magic_2/RBL0
rlabel locali 5799 591 5814 633 1 10T_4x4_magic_13/10T_toy_magic_2/RBL1
rlabel metal1 6059 779 6091 793 1 10T_4x4_magic_13/10T_toy_magic_2/VDD
rlabel metal1 6059 553 6091 567 7 10T_4x4_magic_13/10T_toy_magic_2/GND
rlabel polycont 6021 660 6051 694 1 10T_4x4_magic_13/10T_toy_magic_2/junc0
rlabel polycont 6099 660 6129 694 1 10T_4x4_magic_13/10T_toy_magic_2/junc1
rlabel ndiff 5872 591 5928 619 1 10T_4x4_magic_13/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 591 6278 619 1 10T_4x4_magic_13/10T_toy_magic_2/RWL0_junc
rlabel poly 6379 1063 6931 1093 1 10T_4x4_magic_13/10T_toy_magic_1/WWL
rlabel locali 6858 925 6888 959 1 10T_4x4_magic_13/10T_toy_magic_1/RWL
rlabel locali 6422 925 6452 959 1 10T_4x4_magic_13/10T_toy_magic_1/RWL
rlabel locali 6843 1007 6858 1036 1 10T_4x4_magic_13/10T_toy_magic_1/WBL
rlabel locali 6453 1007 6468 1035 1 10T_4x4_magic_13/10T_toy_magic_1/WBLb
rlabel locali 6916 861 6931 903 1 10T_4x4_magic_13/10T_toy_magic_1/RBL0
rlabel locali 6379 861 6394 903 1 10T_4x4_magic_13/10T_toy_magic_1/RBL1
rlabel metal1 6639 1049 6671 1063 1 10T_4x4_magic_13/10T_toy_magic_1/VDD
rlabel metal1 6639 823 6671 837 7 10T_4x4_magic_13/10T_toy_magic_1/GND
rlabel polycont 6601 930 6631 964 1 10T_4x4_magic_13/10T_toy_magic_1/junc0
rlabel polycont 6679 930 6709 964 1 10T_4x4_magic_13/10T_toy_magic_1/junc1
rlabel ndiff 6452 861 6508 889 1 10T_4x4_magic_13/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 861 6858 889 1 10T_4x4_magic_13/10T_toy_magic_1/RWL0_junc
rlabel poly 5799 1063 6351 1093 1 10T_4x4_magic_13/10T_toy_magic_0/WWL
rlabel locali 6278 925 6308 959 1 10T_4x4_magic_13/10T_toy_magic_0/RWL
rlabel locali 5842 925 5872 959 1 10T_4x4_magic_13/10T_toy_magic_0/RWL
rlabel locali 6263 1007 6278 1036 1 10T_4x4_magic_13/10T_toy_magic_0/WBL
rlabel locali 5873 1007 5888 1035 1 10T_4x4_magic_13/10T_toy_magic_0/WBLb
rlabel locali 6336 861 6351 903 1 10T_4x4_magic_13/10T_toy_magic_0/RBL0
rlabel locali 5799 861 5814 903 1 10T_4x4_magic_13/10T_toy_magic_0/RBL1
rlabel metal1 6059 1049 6091 1063 1 10T_4x4_magic_13/10T_toy_magic_0/VDD
rlabel metal1 6059 823 6091 837 7 10T_4x4_magic_13/10T_toy_magic_0/GND
rlabel polycont 6021 930 6051 964 1 10T_4x4_magic_13/10T_toy_magic_0/junc0
rlabel polycont 6099 930 6129 964 1 10T_4x4_magic_13/10T_toy_magic_0/junc1
rlabel ndiff 5872 861 5928 889 1 10T_4x4_magic_13/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 861 6278 889 1 10T_4x4_magic_13/10T_toy_magic_0/RWL0_junc
rlabel metal1 5751 2130 5781 2144 1 10T_4x4_magic_14/VDD
rlabel metal1 5751 1860 5781 1874 1 10T_4x4_magic_14/VDD
rlabel metal1 5751 1904 5781 1918 1 10T_4x4_magic_14/GND
rlabel metal1 5751 1634 5781 1648 1 10T_4x4_magic_14/GND
rlabel corelocali 5799 1586 5814 1616 1 10T_4x4_magic_14/RBL1_0
rlabel corelocali 6336 1586 6351 1616 1 10T_4x4_magic_14/RBL0_0
rlabel corelocali 6379 1586 6394 1616 1 10T_4x4_magic_14/RBL1_1
rlabel corelocali 6916 1586 6931 1616 1 10T_4x4_magic_14/RBL0_1
rlabel metal1 5751 1736 5781 1770 1 10T_4x4_magic_14/RWL_1
rlabel metal1 5751 2006 5781 2040 1 10T_4x4_magic_14/RWL_0
rlabel locali 6858 1736 6888 1770 1 10T_4x4_magic_14/10T_toy_magic_3/RWL
rlabel locali 6422 1736 6452 1770 1 10T_4x4_magic_14/10T_toy_magic_3/RWL
rlabel locali 6843 1818 6858 1847 1 10T_4x4_magic_14/10T_toy_magic_3/WBL
rlabel locali 6453 1818 6468 1846 1 10T_4x4_magic_14/10T_toy_magic_3/WBLb
rlabel locali 6916 1672 6931 1714 1 10T_4x4_magic_14/10T_toy_magic_3/RBL0
rlabel locali 6379 1672 6394 1714 1 10T_4x4_magic_14/10T_toy_magic_3/RBL1
rlabel metal1 6639 1860 6671 1874 1 10T_4x4_magic_14/10T_toy_magic_3/VDD
rlabel metal1 6639 1634 6671 1648 7 10T_4x4_magic_14/10T_toy_magic_3/GND
rlabel polycont 6601 1741 6631 1775 1 10T_4x4_magic_14/10T_toy_magic_3/junc0
rlabel polycont 6679 1741 6709 1775 1 10T_4x4_magic_14/10T_toy_magic_3/junc1
rlabel ndiff 6452 1672 6508 1700 1 10T_4x4_magic_14/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 1672 6858 1700 1 10T_4x4_magic_14/10T_toy_magic_3/RWL0_junc
rlabel locali 6278 1736 6308 1770 1 10T_4x4_magic_14/10T_toy_magic_2/RWL
rlabel locali 5842 1736 5872 1770 1 10T_4x4_magic_14/10T_toy_magic_2/RWL
rlabel locali 6263 1818 6278 1847 1 10T_4x4_magic_14/10T_toy_magic_2/WBL
rlabel locali 5873 1818 5888 1846 1 10T_4x4_magic_14/10T_toy_magic_2/WBLb
rlabel locali 6336 1672 6351 1714 1 10T_4x4_magic_14/10T_toy_magic_2/RBL0
rlabel locali 5799 1672 5814 1714 1 10T_4x4_magic_14/10T_toy_magic_2/RBL1
rlabel metal1 6059 1860 6091 1874 1 10T_4x4_magic_14/10T_toy_magic_2/VDD
rlabel metal1 6059 1634 6091 1648 7 10T_4x4_magic_14/10T_toy_magic_2/GND
rlabel polycont 6021 1741 6051 1775 1 10T_4x4_magic_14/10T_toy_magic_2/junc0
rlabel polycont 6099 1741 6129 1775 1 10T_4x4_magic_14/10T_toy_magic_2/junc1
rlabel ndiff 5872 1672 5928 1700 1 10T_4x4_magic_14/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 1672 6278 1700 1 10T_4x4_magic_14/10T_toy_magic_2/RWL0_junc
rlabel locali 6858 2006 6888 2040 1 10T_4x4_magic_14/10T_toy_magic_1/RWL
rlabel locali 6422 2006 6452 2040 1 10T_4x4_magic_14/10T_toy_magic_1/RWL
rlabel locali 6843 2088 6858 2117 1 10T_4x4_magic_14/10T_toy_magic_1/WBL
rlabel locali 6453 2088 6468 2116 1 10T_4x4_magic_14/10T_toy_magic_1/WBLb
rlabel locali 6916 1942 6931 1984 1 10T_4x4_magic_14/10T_toy_magic_1/RBL0
rlabel locali 6379 1942 6394 1984 1 10T_4x4_magic_14/10T_toy_magic_1/RBL1
rlabel metal1 6639 2130 6671 2144 1 10T_4x4_magic_14/10T_toy_magic_1/VDD
rlabel metal1 6639 1904 6671 1918 7 10T_4x4_magic_14/10T_toy_magic_1/GND
rlabel polycont 6601 2011 6631 2045 1 10T_4x4_magic_14/10T_toy_magic_1/junc0
rlabel polycont 6679 2011 6709 2045 1 10T_4x4_magic_14/10T_toy_magic_1/junc1
rlabel ndiff 6452 1942 6508 1970 1 10T_4x4_magic_14/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 1942 6858 1970 1 10T_4x4_magic_14/10T_toy_magic_1/RWL0_junc
rlabel locali 6278 2006 6308 2040 1 10T_4x4_magic_14/10T_toy_magic_0/RWL
rlabel locali 5842 2006 5872 2040 1 10T_4x4_magic_14/10T_toy_magic_0/RWL
rlabel locali 6263 2088 6278 2117 1 10T_4x4_magic_14/10T_toy_magic_0/WBL
rlabel locali 5873 2088 5888 2116 1 10T_4x4_magic_14/10T_toy_magic_0/WBLb
rlabel locali 6336 1942 6351 1984 1 10T_4x4_magic_14/10T_toy_magic_0/RBL0
rlabel locali 5799 1942 5814 1984 1 10T_4x4_magic_14/10T_toy_magic_0/RBL1
rlabel metal1 6059 2130 6091 2144 1 10T_4x4_magic_14/10T_toy_magic_0/VDD
rlabel metal1 6059 1904 6091 1918 7 10T_4x4_magic_14/10T_toy_magic_0/GND
rlabel polycont 6021 2011 6051 2045 1 10T_4x4_magic_14/10T_toy_magic_0/junc0
rlabel polycont 6099 2011 6129 2045 1 10T_4x4_magic_14/10T_toy_magic_0/junc1
rlabel ndiff 5872 1942 5928 1970 1 10T_4x4_magic_14/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 1942 6278 1970 1 10T_4x4_magic_14/10T_toy_magic_0/RWL0_junc
rlabel metal1 5751 1590 5781 1604 1 10T_4x4_magic_15/VDD
rlabel metal1 5751 1320 5781 1334 1 10T_4x4_magic_15/VDD
rlabel metal1 5751 1364 5781 1378 1 10T_4x4_magic_15/GND
rlabel metal1 5751 1094 5781 1108 1 10T_4x4_magic_15/GND
rlabel corelocali 5799 1046 5814 1076 1 10T_4x4_magic_15/RBL1_0
rlabel corelocali 6336 1046 6351 1076 1 10T_4x4_magic_15/RBL0_0
rlabel corelocali 6379 1046 6394 1076 1 10T_4x4_magic_15/RBL1_1
rlabel corelocali 6916 1046 6931 1076 1 10T_4x4_magic_15/RBL0_1
rlabel metal1 5751 1196 5781 1230 1 10T_4x4_magic_15/RWL_1
rlabel metal1 5751 1466 5781 1500 1 10T_4x4_magic_15/RWL_0
rlabel locali 6858 1196 6888 1230 1 10T_4x4_magic_15/10T_toy_magic_3/RWL
rlabel locali 6422 1196 6452 1230 1 10T_4x4_magic_15/10T_toy_magic_3/RWL
rlabel locali 6843 1278 6858 1307 1 10T_4x4_magic_15/10T_toy_magic_3/WBL
rlabel locali 6453 1278 6468 1306 1 10T_4x4_magic_15/10T_toy_magic_3/WBLb
rlabel locali 6916 1132 6931 1174 1 10T_4x4_magic_15/10T_toy_magic_3/RBL0
rlabel locali 6379 1132 6394 1174 1 10T_4x4_magic_15/10T_toy_magic_3/RBL1
rlabel metal1 6639 1320 6671 1334 1 10T_4x4_magic_15/10T_toy_magic_3/VDD
rlabel metal1 6639 1094 6671 1108 7 10T_4x4_magic_15/10T_toy_magic_3/GND
rlabel polycont 6601 1201 6631 1235 1 10T_4x4_magic_15/10T_toy_magic_3/junc0
rlabel polycont 6679 1201 6709 1235 1 10T_4x4_magic_15/10T_toy_magic_3/junc1
rlabel ndiff 6452 1132 6508 1160 1 10T_4x4_magic_15/10T_toy_magic_3/RWL1_junc
rlabel ndiff 6802 1132 6858 1160 1 10T_4x4_magic_15/10T_toy_magic_3/RWL0_junc
rlabel locali 6278 1196 6308 1230 1 10T_4x4_magic_15/10T_toy_magic_2/RWL
rlabel locali 5842 1196 5872 1230 1 10T_4x4_magic_15/10T_toy_magic_2/RWL
rlabel locali 6263 1278 6278 1307 1 10T_4x4_magic_15/10T_toy_magic_2/WBL
rlabel locali 5873 1278 5888 1306 1 10T_4x4_magic_15/10T_toy_magic_2/WBLb
rlabel locali 6336 1132 6351 1174 1 10T_4x4_magic_15/10T_toy_magic_2/RBL0
rlabel locali 5799 1132 5814 1174 1 10T_4x4_magic_15/10T_toy_magic_2/RBL1
rlabel metal1 6059 1320 6091 1334 1 10T_4x4_magic_15/10T_toy_magic_2/VDD
rlabel metal1 6059 1094 6091 1108 7 10T_4x4_magic_15/10T_toy_magic_2/GND
rlabel polycont 6021 1201 6051 1235 1 10T_4x4_magic_15/10T_toy_magic_2/junc0
rlabel polycont 6099 1201 6129 1235 1 10T_4x4_magic_15/10T_toy_magic_2/junc1
rlabel ndiff 5872 1132 5928 1160 1 10T_4x4_magic_15/10T_toy_magic_2/RWL1_junc
rlabel ndiff 6222 1132 6278 1160 1 10T_4x4_magic_15/10T_toy_magic_2/RWL0_junc
rlabel locali 6858 1466 6888 1500 1 10T_4x4_magic_15/10T_toy_magic_1/RWL
rlabel locali 6422 1466 6452 1500 1 10T_4x4_magic_15/10T_toy_magic_1/RWL
rlabel locali 6843 1548 6858 1577 1 10T_4x4_magic_15/10T_toy_magic_1/WBL
rlabel locali 6453 1548 6468 1576 1 10T_4x4_magic_15/10T_toy_magic_1/WBLb
rlabel locali 6916 1402 6931 1444 1 10T_4x4_magic_15/10T_toy_magic_1/RBL0
rlabel locali 6379 1402 6394 1444 1 10T_4x4_magic_15/10T_toy_magic_1/RBL1
rlabel metal1 6639 1590 6671 1604 1 10T_4x4_magic_15/10T_toy_magic_1/VDD
rlabel metal1 6639 1364 6671 1378 7 10T_4x4_magic_15/10T_toy_magic_1/GND
rlabel polycont 6601 1471 6631 1505 1 10T_4x4_magic_15/10T_toy_magic_1/junc0
rlabel polycont 6679 1471 6709 1505 1 10T_4x4_magic_15/10T_toy_magic_1/junc1
rlabel ndiff 6452 1402 6508 1430 1 10T_4x4_magic_15/10T_toy_magic_1/RWL1_junc
rlabel ndiff 6802 1402 6858 1430 1 10T_4x4_magic_15/10T_toy_magic_1/RWL0_junc
rlabel locali 6278 1466 6308 1500 1 10T_4x4_magic_15/10T_toy_magic_0/RWL
rlabel locali 5842 1466 5872 1500 1 10T_4x4_magic_15/10T_toy_magic_0/RWL
rlabel locali 6263 1548 6278 1577 1 10T_4x4_magic_15/10T_toy_magic_0/WBL
rlabel locali 5873 1548 5888 1576 1 10T_4x4_magic_15/10T_toy_magic_0/WBLb
rlabel locali 6336 1402 6351 1444 1 10T_4x4_magic_15/10T_toy_magic_0/RBL0
rlabel locali 5799 1402 5814 1444 1 10T_4x4_magic_15/10T_toy_magic_0/RBL1
rlabel metal1 6059 1590 6091 1604 1 10T_4x4_magic_15/10T_toy_magic_0/VDD
rlabel metal1 6059 1364 6091 1378 7 10T_4x4_magic_15/10T_toy_magic_0/GND
rlabel polycont 6021 1471 6051 1505 1 10T_4x4_magic_15/10T_toy_magic_0/junc0
rlabel polycont 6099 1471 6129 1505 1 10T_4x4_magic_15/10T_toy_magic_0/junc1
rlabel ndiff 5872 1402 5928 1430 1 10T_4x4_magic_15/10T_toy_magic_0/RWL1_junc
rlabel ndiff 6222 1402 6278 1430 1 10T_4x4_magic_15/10T_toy_magic_0/RWL0_junc
rlabel corelocali 579 1942 594 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_1
rlabel ndiff 422 1942 478 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/RWL0_junc
rlabel ndiff 72 1942 128 1970 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/RWL1_junc
rlabel polycont 299 2011 329 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/junc1
rlabel polycont 221 2011 251 2045 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/junc0
rlabel metal1 259 1904 291 1918 7 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/GND
rlabel metal1 259 2130 291 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/VDD
rlabel locali -1 1942 14 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/RBL1
rlabel locali 536 1942 551 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/RBL0
rlabel viali 478 2006 508 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/10T_toy_magic_7/RWL
rlabel metal1 -1 1904 14 1918 1 10T_8x8_magic_0/10T_1x8_magic_2/GND
rlabel metal1 -1 2130 14 2144 1 10T_8x8_magic_0/10T_1x8_magic_2/VDD
rlabel locali 536 1942 551 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL0_0
rlabel locali -1 1942 14 1984 1 10T_8x8_magic_0/10T_1x8_magic_2/RBL1_0
rlabel metal1 -1 2006 14 2040 1 10T_8x8_magic_0/10T_1x8_magic_2/RWL
rlabel metal1 -1 1904 14 1918 1 10T_8x8_magic_0/GND
rlabel metal1 -1 2130 14 2144 1 10T_8x8_magic_0/VDD
rlabel metal1 -1 2006 14 2040 1 10T_8x8_magic_0/RWL_0
rlabel ndiffc 73 2088 88 2116 1 WBLb_0
port 1 n
rlabel poly -1 2144 6931 2174 1 WWL_0
port 2 n
rlabel pwell 42 2006 72 2040 1 RWL_0
port 3 n
rlabel ndiffc 463 2088 478 2117 1 WBL_0
port 4 n
rlabel poly -1 1874 6931 1904 1 WWL_1
port 5 n
rlabel poly -1 1334 6931 1364 1 WWL_3
port 6 n
rlabel poly -1 1604 6931 1634 1 WWL_2
port 7 n
rlabel poly -1 1064 4611 1094 1 WWL_4
port 8 n
rlabel poly -1 794 4611 824 1 WWL_5
port 9 n
<< end >>
