* FILE: 10T-toy.sp



* SPICE Header file for TSMC 3.3 0.35 process (scn4me_subm)

.OPTIONS post NOMOD probe measout captab 

**################################################
* Only Typical/Typical spice models included
.include '/programs/micromagic/mmi_local/ami05.mod'
**################################################

.PARAM vddp=3.30	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 25
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "10T-toy" generated by MMI_SUE5.6.37 on Fri Nov 19 
*+ 07:57:02 CST 2021.

.SUBCKT invM A1 O 
M_1 O A1 Vdd vdd p W='0.14*1u' L='0.15*1u' 
M_2 O A1 Gnd gnd n W='0.21*1u' L='0.15*1u' 
.ENDS	$ invM

* start main CELL 10T-toy
* .SUBCKT 10T-toy RBL0 RBL1 RWL0 RWL1 WBL WBLb WWL 
XinvM net_1 net_4 invM 
M_1 net_1 WWL WBL gnd n W='0.14*1u' L='0.15*1u' 
M_2 WBLb WWL net_4 gnd n W='0.14*1u' L='0.15*1u' 
M_3 net_2 RWL0 RBL0 gnd n W='0.14*1u' L='0.025*1u' 
M_4 gnd net_1 net_2 gnd n W='0.42*1u' L='0.15*1u' 
M_5 RBL1 RWL1 net_3 gnd n W='0.14*1u' L='0.025*1u' 
M_6 net_3 net_4 gnd gnd n W='0.42*1u' L='0.15*1u' 
XInv net_4 net_1 invM 
* .ENDS	$ 10T-toy

.GLOBAL gnd vdd

.END

