* SPICE3 file created from sky130_fd_bd_sram__sram_sp_cell.spice.ext - technology: sky130A

