magic
tech sky130A
magscale 1 2
timestamp 1655151891
<< error_p >>
rect -91 235 -78 251
rect 10 249 23 251
rect -24 235 -9 249
rect 7 235 37 249
rect 98 247 251 293
rect 80 235 272 247
rect 315 235 345 249
rect 357 235 370 251
rect 458 235 471 251
rect -106 221 471 235
rect -91 117 -78 221
rect -34 199 -33 209
rect -18 199 -5 209
rect -34 195 -5 199
rect 7 195 37 221
rect 55 207 71 209
rect 143 207 209 221
rect 144 205 208 207
rect 55 195 70 199
rect -34 193 70 195
rect -43 185 1 193
rect -43 173 -25 185
rect -18 173 1 185
rect 39 185 89 193
rect 39 177 55 185
rect 62 183 89 185
rect 98 185 113 189
rect 160 185 192 205
rect 251 193 266 221
rect 315 218 345 221
rect 315 215 357 218
rect 281 207 297 209
rect 282 195 297 199
rect 315 196 360 215
rect 379 209 386 210
rect 385 202 386 209
rect 369 199 370 202
rect 385 199 398 202
rect 315 195 345 196
rect 360 195 366 196
rect 369 195 398 199
rect 282 194 398 195
rect 282 193 404 194
rect 251 185 319 193
rect 98 183 319 185
rect 62 173 134 183
rect 152 182 160 183
rect 192 182 200 183
rect -43 165 1 173
rect 55 169 134 173
rect 215 169 319 183
rect 354 185 404 193
rect 354 178 370 185
rect 55 165 319 169
rect 369 173 370 178
rect 377 173 404 185
rect 369 165 404 173
rect -34 149 -33 165
rect -18 145 -5 165
rect -33 133 -5 145
rect -63 117 -5 133
rect -91 109 -5 117
rect 7 109 37 165
rect 72 155 280 165
rect 239 151 287 155
rect 122 129 152 138
rect 215 131 230 138
rect 251 129 287 151
rect 98 125 287 129
rect 113 122 287 125
rect 106 119 287 122
rect 315 141 345 165
rect 351 144 366 156
rect 369 149 370 165
rect 385 145 398 165
rect 370 144 398 145
rect 351 141 385 144
rect 315 128 351 141
rect 357 133 385 141
rect -91 103 -15 109
rect -91 101 -17 103
rect -91 99 -78 101
rect -63 99 -29 101
rect -91 83 -17 99
rect -15 97 -9 103
rect 10 95 23 109
rect 38 95 55 111
rect 106 106 117 119
rect -107 61 -106 77
rect -91 61 -78 83
rect -63 61 -33 83
rect 10 79 72 95
rect 106 88 117 104
rect 122 99 132 119
rect 142 99 156 119
rect 159 106 168 119
rect 184 106 193 119
rect 122 88 156 99
rect 159 88 168 104
rect 184 88 193 104
rect 200 99 210 119
rect 220 99 234 119
rect 235 106 246 119
rect 200 88 234 99
rect 235 88 246 104
rect 297 103 314 119
rect 315 109 345 128
rect 357 122 415 133
rect 357 117 370 122
rect 385 117 415 122
rect 284 93 330 103
rect 284 85 294 93
rect 313 87 330 93
rect 357 101 431 117
rect 357 99 370 101
rect 385 99 419 101
rect 313 85 318 87
rect 10 77 23 79
rect 38 77 72 79
rect 10 61 75 77
rect 122 72 138 79
rect 200 72 230 83
rect 284 69 330 85
rect 357 83 431 99
rect 297 61 314 69
rect 357 61 370 83
rect 385 61 415 83
rect 442 61 443 77
rect 458 61 471 221
rect -113 53 -72 61
rect -113 27 -98 53
rect -91 27 -72 53
rect -10 49 23 61
rect 29 49 59 61
rect 72 49 147 61
rect 205 49 280 61
rect 293 49 323 61
rect 335 49 370 61
rect -10 47 160 49
rect -113 19 -72 27
rect -107 9 -106 19
rect -91 9 -78 19
rect -63 9 -33 19
rect 10 9 23 47
rect 38 45 55 47
rect 29 9 59 19
rect 66 9 74 19
rect 80 18 90 28
rect 93 20 160 47
rect 192 47 370 49
rect 192 20 272 47
rect 93 19 272 20
rect 93 11 96 19
rect 160 11 192 19
rect 93 9 259 11
rect 278 9 289 19
rect 293 9 323 19
rect 357 9 370 47
rect 442 53 477 61
rect 442 27 443 53
rect 450 27 477 53
rect 442 19 477 27
rect 385 9 415 19
rect 442 9 443 19
rect 458 9 471 19
rect -107 3 471 9
rect -106 -5 471 3
rect -91 -19 -78 -5
rect -63 -23 -33 -5
rect 10 -19 23 -5
rect 66 -18 74 -5
rect 107 -14 245 -5
rect 107 -18 200 -14
rect 129 -19 200 -18
rect 209 -18 245 -14
rect 278 -18 286 -5
rect 209 -19 223 -18
rect 357 -19 370 -5
rect 144 -21 208 -19
rect 152 -27 160 -21
rect 192 -27 200 -21
rect 385 -23 415 -5
rect 458 -19 471 -5
<< nwell >>
rect 98 125 251 221
<< pwell >>
rect -106 87 70 251
rect 78 164 91 171
rect 282 87 458 251
rect -106 -19 458 87
<< nmos >>
rect 7 165 37 193
rect 315 165 345 193
rect -63 19 -33 61
rect 385 19 415 61
<< npd >>
rect 122 19 152 61
rect 200 19 230 61
<< npass >>
rect 29 19 59 47
rect 293 19 323 47
<< ppu >>
rect 122 155 152 183
rect 200 155 230 183
<< ndiff >>
rect -18 165 7 193
rect 37 165 55 193
rect 297 165 315 193
rect 345 165 370 193
rect -91 19 -63 61
rect -33 47 -10 61
rect 97 52 122 61
rect -33 19 29 47
rect 59 19 93 47
tri 104 42 114 52 ne
rect 114 19 122 52
rect 152 19 200 61
rect 230 51 255 61
rect 230 19 238 51
rect 362 47 385 61
rect 259 19 293 47
rect 323 19 385 47
rect 415 19 443 61
rect 66 -5 93 19
rect 160 -5 192 19
rect 259 -5 286 19
rect 66 -19 143 -5
rect 209 -19 286 -5
<< pdiff >>
rect 160 183 192 207
rect 113 155 122 183
rect 152 155 200 183
rect 230 155 239 183
tri 239 155 251 167 sw
<< ndiffc >>
rect -33 165 -18 193
rect 55 165 70 193
rect 282 165 297 193
rect 370 165 385 194
rect -106 19 -91 61
rect 97 42 104 52
tri 104 42 114 52 sw
rect 97 19 114 42
rect 238 19 255 51
rect 443 19 458 61
rect 160 -19 192 -5
<< pdiffc >>
rect 98 155 113 183
rect 239 167 251 183
tri 239 155 251 167 ne
<< psubdiff >>
rect 143 -19 160 -5
rect 192 -19 209 -5
<< nsubdiff >>
rect 143 207 160 221
rect 192 207 209 221
<< nsubdiffcont >>
rect 160 207 192 221
<< poly >>
rect -106 221 458 251
rect 7 193 37 221
rect 122 183 152 205
rect 200 183 230 205
rect 315 193 345 221
rect 7 143 37 165
rect 122 122 152 155
rect -63 61 -33 83
rect 29 61 38 95
rect 122 61 152 88
rect 200 122 230 155
rect 315 127 345 165
rect 200 61 230 88
rect 314 69 323 103
rect 29 47 59 61
rect 293 47 323 69
rect 385 61 415 83
rect -63 -3 -33 19
rect 29 -3 59 19
rect 122 -3 152 19
rect 200 -3 230 19
rect 293 -3 323 19
rect 385 -3 415 19
<< polycont >>
rect -63 83 -33 117
rect 38 61 68 95
rect 122 88 152 122
rect 200 88 230 122
rect 284 69 314 103
rect 385 83 415 117
<< corelocali >>
rect -106 61 -91 251
tri -27 215 -5 237 se
rect -5 230 10 251
tri -5 215 10 230 nw
rect 342 230 357 251
tri -33 209 -27 215 se
rect -27 209 -18 215
rect -33 193 -18 209
tri -18 202 -5 215 nw
rect 143 207 160 221
rect 192 207 209 221
tri 342 215 357 230 ne
tri 357 215 379 237 sw
rect -33 137 -18 165
rect 55 193 115 207
rect 70 183 115 193
rect 70 165 98 183
rect 55 155 98 165
rect 113 179 115 183
rect 237 193 297 207
tri 357 202 370 215 ne
rect 370 209 379 215
tri 379 209 385 215 sw
rect 237 183 282 193
rect 113 155 187 179
rect 55 151 187 155
tri 187 151 215 179 sw
rect 237 169 239 183
tri 237 167 239 169 ne
rect 251 165 282 183
rect 251 155 297 165
tri -33 122 -18 137 ne
tri -18 122 4 144 sw
tri -18 109 -5 122 ne
rect -5 116 4 122
tri 4 116 10 122 sw
rect -106 -19 -91 19
rect -5 -19 10 116
rect 55 95 83 151
tri 175 133 193 151 ne
rect 193 131 215 151
tri 215 131 235 151 sw
tri 251 137 269 155 ne
rect 68 61 83 95
rect 117 122 159 123
rect 117 88 122 122
rect 152 88 159 122
rect 117 79 159 88
rect 193 122 235 131
rect 193 88 200 122
rect 230 88 235 122
rect 193 83 235 88
rect 269 103 297 155
rect 370 194 385 209
tri 348 122 370 144 se
rect 370 137 385 165
tri 370 122 385 137 nw
tri 342 116 348 122 se
rect 348 116 357 122
rect 55 52 83 61
tri 83 52 104 73 sw
rect 55 19 97 52
tri 117 42 154 79 ne
rect 154 51 159 79
tri 159 51 185 77 sw
rect 269 69 284 103
rect 269 51 297 69
rect 154 42 238 51
tri 114 41 115 42 sw
rect 114 19 115 41
tri 154 23 173 42 ne
rect 173 23 238 42
rect 55 -5 115 19
rect 237 19 238 23
rect 255 19 297 51
rect 237 -3 297 19
rect 143 -19 160 -5
rect 192 -19 209 -5
rect 342 -19 357 116
tri 357 109 370 122 nw
rect 443 61 458 251
rect 443 -19 458 19
<< viali >>
rect 160 207 192 221
rect 160 -19 192 -5
<< metal1 >>
rect -106 207 160 221
rect 192 207 458 221
rect -106 -19 160 -5
rect 192 -19 458 -5
<< labels >>
rlabel metal1 160 -19 192 -5 7 GND
rlabel polycont -63 83 -33 117 1 RWL1
rlabel corelocali -106 19 -91 61 1 RBL1
rlabel locali -33 165 -18 193 1 WBLb
rlabel polycont 385 83 415 117 1 RWL0
rlabel metal1 160 207 192 221 1 VDD
rlabel ndiff -33 19 29 47 1 RWL1_junc
rlabel pwell 323 19 385 47 1 RWL0_junc
rlabel corelocali 200 88 230 122 1 junc1
rlabel corelocali 122 88 152 122 1 junc0
rlabel pwell 443 19 458 61 1 RBL0
rlabel poly -106 221 458 251 1 WWL
rlabel locali 370 165 385 194 1 WBL
<< end >>
